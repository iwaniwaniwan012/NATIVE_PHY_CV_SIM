`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LZhgbdYFB9OlSTgsUxcj6hGTTJHKZu8nGproYnWQGgV9covCwcCnI304jWnMBQtR
esr8a1bmc2rToIr69+Bd0QkaiaB6uk0B6PXjLbBktNmniKut+qXmL6jREvx+QWPK
cLDXS657l6blVjmDFODF+JNRyAb3CFNwJNloiwTLNwY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7360)
c3ASSqdn9zCcWbWzLkWE8KcpIX79Frk8vKPwz4qUc/vgSBZ0VFLRquxB+XwuuGld
zI0cWHyc2kuGPqIKdrhrTBG7D/RERe716lTzZIU9bJobvelnE1y5PcrSiHEhX/jG
L5Fr9vtr/eLlRIFCnxca8OC5fdPFhgXstVWSVky60dyHt3YMpjOjAQWg+AJmo/Wd
uB3JitpvPoAPViTvmvLrawgUoTZmzkY6PEDTt2+tQufwspAD8jLPwauMRzZ2FWFF
UR50709dlAKH/l0s4DfP+jvzYYtkS82pm5+LaEUYgHZF9x2ErYXP6tiK+VjLYWk+
4OW/AnIVJ1h8B9G1Gjc3fuJY4iBypPQkEKv2GJFWj7ytRXJvGDaXtw96sXhom6/4
7rVNIP9umaL2Jrfk7aSGW/6O4ZRwnI1iUe7tU5Fc+M7OhxDFx3FfQldxDUZGoEOJ
ncOzmoaDVIhZlTklGSYbUToyfVNeUDzQY1pFFdOmxAHhxNs1+JQvssHDs9JTzh7r
qoITCSnsU9EHdeF9m8tXR73gfEf7iQxWa+o+ktZZQM+iDKfg66AS2ATchq3r6RpO
FGw1SaU5rCGXUHbcAMq1Mr8da2txZGss1qJtmhHMrOshz+YM094G2w+5Rh7QdHY4
AzcyxbbV1sxgfo9sMmQUuhxFV7xrkSqZ+9tvT0QjuVcpPYzrCaOn1ImDNGiiZt8e
NQMV9sShSnH/2ZfvWe9UciMtw4KeMIuldtl9xCFzTHz7kmBlLJhCq5TfexhrNcMZ
smHuV7D6ShkE4SlxY8p3FqVcGNdzPA8vDsL9sj895ra+KgNnrr3Hu15yp/Q0JS3I
xzebXAe8ye5yd6q0RFXO3vJcUkA8Il4dLBb0/RRvNbNNuJ7bZpBdlPeBcJxhwSBB
NEJy52UPZ9wRXMQhm8jRpGDWEScNqz0cwIPCOOFE/jAkx/k9sczEgcY7o2t7oIvZ
4aBboMz5dgrZAsU7zfs0bNnxcwOcBQWKEGbvx21/lGZpKCZOWA0bOqlvSkb5jNOV
Xrw3KXEpy3Qiv3EJbCkDg+Q4RKdigf3t5oUgX8rZkX6FeXUs9DgVSAIAYN6yEUnc
9SSycqx++MsuP1VTj8nP9cut06xmA/KL6w6IfESE/fygtarYK/ipPG0DT0baubOO
8Hla2j2Cv1feYQ63Nmhgulk4wmW8s4RmcxgoLhmpKnVv4NeTwgaiGUBMQGGsu2Tk
WgJCKS8S8yWp4V3BShPmaLfYYm9W1gID78DP6XPqI+uxVigqLMZwDnGwZyPoIhsm
Cbf/8/Sg6m3n6fwvx06WFDppYj5yfYTb4k/OcE1LhX12xnk29t5UjXRn+KnRzE+k
8MURoCATOaOuEW4p+8ehxRwwQrkCq/7tC/hktmVLknycSoYVDoT3L0yd0O6P+kus
sFMYjmLa45DiVb8q2/zwutz+j/Hh/nHM3ZSZzXV7OhvHNGOMXOr/iKXHkMpMUhGx
dhStKnCZiZE5z8R9QeNQaEqrOcnmhIviRr1CJHZety5BGU73G3i/x9lZgn3ylfrQ
RB4FJBpz0F6xmXSEQtUYqkVxL1+G5vyG3uzJRYAIXhP6WrGwoPn8UcvdOOF8bQe4
sqBKDjWgb5i7elLMI86HVufRam0agFxgbIpeJBsMmv/Ezfz8rvY840IxbfkgjJ0I
i4YUQolJAkL6ZnMhMU16Uxy9kBO0+SlHBZHFYWbiVFDgpdZkV/qWTca1TIIyLqd0
JtyX5Q9DmBoA/kSynigXxtcw05HEm8GOFqTz+kjO9zEs/7LYSZ/nASDaJNuDK1ZN
AKUtZ0LWyJp5MNwIi7A7R7m6pdQItQlpB4C5DICYsTt7Lk1seJ6kudRv4eqWwmOy
OPcFbjW6Xkp2OVHRqjDJQ2iayUtonvwGIahR696ZVEmQntBaLhUTI0TjvnP8UCbm
5E1IGRosov2YFAQ6QBFx0WBxAeQ5EV/vy9ldjM2Wge+goHUJiuDhPJNL+az6tPLI
PgjIKJlHHsUljizDxGXc/4BBDzPpbENDnmreIg3y+DP4Rk1cfZRL002bEei09XEn
clZsMe0Mqx2fO2gSWondiSGDJD7u/BAM2baN9iazaKEI+ShwITtDzmJjvACmG719
vz5m3+/W2g6o8u2i1Q2NjC4aUIz6K/XpllrXP/Lieujnd3A7KbJ1VW15I+plgTuc
Vuf5nB8y7fbA4CMTQvOtFKtkigxLlRrjWiHeOSrXBtuCnf+dYLtPMprlXLkvBHSM
MDytCP2mvt/aIfwJgGH/i8HXkTzd1c6fwG7QmqTB1GnI50pBP99SZ2bw9+dNuBmX
r6dexo53uPds+xNR5sEO+ChSDKgDdyS879/eQqBuIDsNl4erDB11P0S08XKIvn9i
XfQ7rybMj+1qnpwdMenpVd1Zu8EmMoimos+mmDuYNhoDfjO+To0sWbPmK6WyEpIR
Z91rRrhtQnyMnUiZCUQWi4inMYlSH6NHGgfk7sYGIfZkCixfM/N3TRcVAb6rdN4V
FW39p3hzsZj6ftKk23k41Hn/VLRDZPRtDew46xtZx0/YYnDPnJWzvpmatncpbmZt
Zd0W9BAqxwXfzCrgNiaKBcZiowArj5OcHYMmbmZJBsG0WOMrQfACWMctCBalnAI5
SviBeLj4R/lSmRWFiS2WW8czG3LVxbGwkGHBDLiXM1BwOyxa91M/TZ0i9WerXVCr
V0VzyHsYvrL8XwaXYYmUvaHyOg53NqikpR+LZorpDj9tK4w8AuEa86PFYdy6s4nd
CHOlFvSTDuYI3U4WQrz5Iql3Z6oAkFyL/ZFDG3IHaU8/PPIXWAaWNs27Q0V3WR34
6pTfrcpZCdDljmx4UNQ5VeQ0/7tZOvfzsjOAPALrnIoteXp31l1ub4GMAS4Se06U
aXzeNcj2Fa/V02VDy5/XVfN45l+LZKmxf/zqoRQNJJdGdKhklXxN76lkHIWZy4at
f6IIkFDMUHsk2GwDR0Kuz2Z+40/93/Y2n/3GU80rpb1oqXS69kQU4lfLzKuZNHcX
zWNFWjdJ7b4GD/X38ScDH7nB3wqSyPPRWm+GQo5mGmq+WZN6oAhrPVoBGHXSfBsh
tcBdC5eFQwsH5GTqDoJNGTODATu5J6D0E+dNUnkrk4hlxfaF6vP0x0Q4dtTjbXUO
MZzjk5A2kGCO06IGG/vbsDlU8pV0XelVpObrk8sIcq1fR1SSAE+6xnpESJmpLWBL
MenNg/3YMgiNqFwy3qNBwKeKsNgJ3+NeZ5Y1G87JQZ/qT7X++t+lfucUpnEe6N6u
5xV6Wrff9pjmFOG8H/J5uj6xg5ocN1IR6r1e4hDJJ4mgYHBe1SyFIBDsSjYfGT8O
VUSPb4mMumKLyuGnjqWRsneW41qiMd+na6R1ZhHXKOTKmdWubYWuBNLmGbqWrVC5
8K9G/vCl/fE1102OUTCrxDeJ0ukJr1H1Ny4n6laAg6bA9WfMWqbrj0F+p7VX7Nv0
48wjxR7USPiVzuHBzKn5djzdPb3M0iyYOTr15+DaIXEw9dK2PhpGwGcsrk6m5uYS
tDnMDeo0sA4596q1M5Ox9XO1BCISrEKru1aPX+m7dYUaXm31MoRGHvbKKXvw15Nu
xrfIRJPyc6maAgn6gEyO/FLGdKT+V5AS5Jo6NPHE+E44IylcAW9FLx3uuY/0x9QI
By+QA9/sy8lpIm/AhmCaHrSmeGfkk9aGvQ+c/AJ15CowaUnMV0BIxA7taul9tGpp
y5azqGrL3t9kBk2nqDGebxf1r0uBhfPS0Qpd9uz2F/FkB7HZNIOt6AnYkgf7FwNG
g7iZqMs0oYSJbUyibcSfCa9bPgsTUwhCdPBL5ZB8aY+HnirvnVa/QT1oPjpZ9txW
uVY+dT+CJuK5XId8s0khj4NEuMc7UsAUupT7C4M4uDGAWtjFm+8vSvtRb1ulndjX
lf2ORCJr/5p1oCf+WKIiDeXIaU0t/75nkhIB4daMUCxdkyakox0G0NhQAuTuVzML
watoNCoAlp7g/OM9I10IxFvl+bae+vTWLM3/OQB5kwr3Con7d7YGugjI+bXvXH1P
yrJZ8pjSLbxjI80qEKe68UHxNi1+RjxaSWvuInLyeFKMsbxisTEdVU8KC/NtPHwd
7lEYWtlIHNiAWh50h8J6wVQtL3E6fMlRuLI6O0Uz/fnpV2vCxJP/NoMvv4MbTKaO
zvrd9TsKyNLZ4FSAG5AqHfQDUatgtRHHW/TrdSDo65RDvHrvchahOrzt7wROF91i
CL06fJXerJ5YElkesBfK9JM8q2yl+XV1Psn4gDBzuWeOqLF+PRPxrkbdXLykV/4c
1dFmzjcYWoL36qeZZRAuHiUv1jUcFZfyl2w/P0APjHriy/PdZXU5sdgfhyGNbT3A
Dpno9NDBNC2w5VoV8k9fSr3rJC5gtGTYIENF8sGyxMSH7rod70/wzNvEo3gqnt82
dzaDzOfTD23SErR7hsFq3wirenaQzlZdh728L/7Tufh0pVeOsaqBr5c6pF/cnMsv
sc+F8Nx8X/zB3w4hXJorbAf2vYKIYGprj6X3rj4XqL0Sm+V/0R/riU9No1+avYRO
F19Shuk/ksYUIGekMdVe+jjnlMhsgP+0oyWOxM1tuEMpw4hoPP9I26desbHpbSMZ
037WELyBw1SAKsrW/OJ4XjUidiDMJ24EdBBW/SKm47KRYjcz0fYWi75l/aOl/xOY
hg+xn6xQOwSyAYGiM78T9ornoIUJWklb/8KHuq9eoQBrqGF2gK4mNixksaPtd8rN
0HN6mzfY/nOjwYDVnfseMliKIuiGPUcFDCe/H2k3/s0SHO3RW00vsfsvw5XWg5/H
VEF7lyuK9nEjlZNowA4uV3Rn2smA1weIO5BzOFO/ypYf2hMJTXdPpwmXQvErTJki
//004Lc5TOyAvXkf3ZGE1DBfqmsFvujpX3W07DnyMGIrdZy2q931wDIR6IOkL6Gi
QWDkeZDJbYJe+EyZWjTgpQpSXYTx63Mq2//+udKqzg59HfdJO/1Hp7jZHTNhTaJl
pcBymA4cLDhqTNtuam6OCIVc4w/WgQnK2xLrcZHT6lGuo9GAZLgNm+x2/LvMheek
RPNi4bZGJ3S3pr85yxawwdTtk6R4nzvcqRfoU/MRnZeZNFO+bJnE2btXMfSCVdtJ
qy8itU84ovO1gs01BU7fRTcZFiKsp/0cB9Jdgwbz2Wx6ZAHWhPYgOakPW7UryaHv
ZHhUHhLatprmjClm9DTqndDbDStsxmCN89kImT8/zjGThjZu1u78Bz+TVTbQaLHO
0TAd1jnRMvUtINMfYvhUpcg38s6ymNapxLbVbrQVoXYmauWLaggxLgkOmzDfpzSZ
+pGRJDdvrTVTPhPF9VacqhWkgo+bI7Twg+Blyp5/OdGxKFj5rj9HX1KFZinwoI2u
rddcqr1QFvysW56/mbWs/rR00vEUmhm7E0Zrm8XOKtjGE5n5ErYVFvlr4KW1QJDn
Rqmuaf2czPt1qPZCdqV1At5oMpVKWHm+sAMdfUXXb5GEH5BYAdB0PhMb6GpB7P1W
LelxuHGPubnip+yCYHLbkalUGefx06Kpc2r8j3X8gQss8p59aVWcGDQE3Iv+sODH
MuPBKBu9ug2Fp5GWQCxDXfyEj65QkwrrY3ZgXyPG0eaLBtLrQ2/pMzycPvzdxIQy
gBM/DG8nYEI4440lfn5cq3g04BRxf6RI60m0jHfRRZNQxlO2pgjA9FUdowSGittT
6XuYygI9s6m75Qz+D+nGy/rv/pDNAErRuQ7BoNG7SwqtaELqso+agj1ZwV+ddGrt
CAhIMSGh4MknDZyJQwW0u0rRwGne+Os8lYWd0/ldtWupOKBuvRubr1zNJ8wypBPn
IOlwtHgt3THBr2g00ARgtcPx8sRv8Do6l4UTvnfQRs+w/ICEt8qNQuggu53sLE2k
gT6VYI1kexLDV+IFaFD4NBNKRY6sJE1I2V7qCIcZHLnzmWSTybDaGTs0C2q9eAUV
Y765qwvIjLxhrjsihdAJSjvnqxNU3LJGABRJXiGV+IeTaIOKLKE01O9iQX7r3TPo
PdqztLGi6cC+c0xSyhrgAnCVIVIXneT4I72dcwaVSHFmR88xIGetLnQPd5O/hO2q
5SHJq6081BDrBDKVs7Cabyobmc/vdvMLL/P5oV7XG+CRCZX8obvfeskwmTyhDA0U
LbnN+TiM9wcVo0y2F7sSi1z7qeA3AhKwnrVdR7rvLQWB+ffF+LjQ3p/NuYOvwBJQ
NhtKsBNV7JI3aFYV1NrApJKWLxkqEWWR4jFM+0kX+sKa8hJYtGxQv8vVrlTsE9yH
Eol867Wb6XFg92aKRseAWjp7lFiGRKBldhRzfzSELCOiQvyBzfjFJO/5DqSPWVAv
OO1FLNykzqZ57NDsT86SwXNNNwIjTeiKjXo7RFkkIlt88cZvtEZNLKiPJL/dHHnm
nGO/eT1ub8QfeVQ9c8HTtws5Mw5TAUWYE01TBRtXONCJCHgNp0dczTBJPYdf7D+Y
wgMVNGxo34VBPIR0Xrcu2BqRXgUwJjoflMVU3KMEuSkaWuolNC+Km/2aChO73xcq
kL9DAZ3Zf52Kr+wECB4SbIvAfy+nlxQ3VuYA+I36kBPDkp+b6kWhiWaKgzwmwtAh
Uwf+zC3iGmr6W16z0sYBS9mQSf+yYgcJ8WFB3OQgs9YMJ9V9vcNVn3qhtBRbUDQW
2Zr7677UDHC6OWdCinb7KINQbWjLf7KZlCAeXXiP2nIY5RYoccPXrYWO8hPzccSS
55g+md+LRSZxPjeXP7XdShuNkK3Se2hWO/HMGYg3lhLwtr2Bw0b+nGWdDGrCzAo+
Jfv/ZKAsxErK9kyjM15xZieEy5CzmLBhK1CSOWJ68LwO5yuygZxs6194CyTGOpeT
Eyl46HAcSTBGE7tPSqH8nKDpLZwoCWptWrQUUY5X8Pqz/qfunLUUuEK4x+w8Atk8
a2e9lYLOFYvAom1q/9mxp5V+mGQwoIZFo3n2cbpECvCqu6wzKhXdehfjW/I89K3j
1W5idpGoOLBULA10TXLXrGvZY/Tm9qUKhVjqUZ9HSmCAYX0zo/GjGk8dcagt/xE8
OhswB9C5UNr7t9yVyWIaFbyEAWqKeyxLLJKRC4kGdHUBgO4o+7++uo5Q0Pv60+lR
8Zx1+lOapIdT7rrOKoGD+Aorhe1ZvZzaAY7Da4aPaWWQzBiHv/x5xG2ua9VxbE0S
qA5TQqNGwRRoBO13dBwMFg94odqPtsj98ElXgImF6Yva4hLtA+yBc7rOODPaQYOE
3IinBBWtYhqk1ocbTZ4NYeQmFHTPADMhJ18inbnTSkKwk5DLArpBnzX4Woo2Vc8F
/3ZHT4BPrDQGRZeM3kfkTpA2M3AFkEvWXC1q8Ji3yc78FEueyTzZ3GAGPXKTNi0J
HVEmrz0xjf7Cs+NuPJdZ0igq3vamNaDKNlQ51Qkn1VoGtE9UJOMEFDSuk/B3AUf2
aAuVaU1iOn2NoSs1Tq5IxQkzLBTtGgntCRwtMSXaSFlfyEVanBitwT/4xWAmT8zf
6i5ySnK0WrBLYUdvg4XjRUcHcnO0J365GFyKklkbznm89xoW+/zAKZ0ysOhCPEcE
6NvAhX2hH3yaUeV5fzLJKN/bliXTgkW93Cb0lb2BFdpTBzJRFbwumz+BPcp9JvFa
uvzMYW6vHZ3cJHYpRBEPRSHbDBPeX8weVOs5pAd0dSVokz3hSX83FefHUHVfKmBl
bGfx7jUIEnAZD/ZXsZNByoA9Kr+rFmAJUZ07noHd7XyMPgBR0WxSlPhoTvPyw3cA
TmVBYAVH3pkBI/CSLuIwefV/f79DjvIjyncuJYDSXI+JhjjGiy3nUuQNwVpe5DIs
ntibM+eoNlpJGZ7FHCfjA5XijlFdooK9qCkkeqG+SNOyAy+Asoj4Ipa1q+OF2OVi
mMWVMCwBvmc4fHDAEosykFDifPnyBhF0Pbq1esSpTmjIun6tg7hQX7UIozCoyxhG
h9F+IAV4+eoUfTipw1x67YCVn+iVPhdAXqEirWj/NPonWPaaQWAN8tEK244yjknJ
0pL882KR9yC3ELUtuRI1uUaj2CCrBf2TVUDF72f1WJioYuxFFiR+e1U7EFn3dwAC
SJTY8l4clRuua+Mzf3Qlq4enG/+t6f3QzV6JX90MJFCYsuoGA4Gpff0Og14Wm84U
FUqVZbOxcoXciCPzBqm3cANLCEfizs1R9q9gwGEXW6nwse13J2g7RXCxI+68zGOc
1bW7qaZzwdtDfeLWc4zLs9DU8pzl1mtPGvs62SI2pId0Aq0c+ONWeoeOdyeq3Dh2
lPFgZH38bFEcYgGUoM812gnNa/2GvOcjBguqE3Q8LQ6sg3InhwaeOgPDWMruYysG
2+ljM2UX8ylEFJirI99dlWjmXAxT1OjtcXBHCEcg6eR3F6KS2imJnmOwMNQfG+e1
fO6+EB4c5rHKL284s0PV/8nco12M6lZtE+6m3K+LrDO+r8l3RpeE5v0ea1DuwLj0
QiC4zB/g5hnHjzu8BgoZdB1YdkM0+9IdQ2Lu1OHuorQsQLP3A/1lPj+jPmU/JCg8
yE4iV1CvDqnQM2xtN7UfhbFItj7sAQMjFZH6d1LThxynl+9VtFvf2yBCS8K1rNtT
SS+0Rgvwd2Om7migwvXkRVFeDVFu9qmRMwV4MVS9s8Z7wHwzX7gba4QwYo8+N8qH
oNpnZk8/VIR4VK0VpXSD8Wj/ESxRWN/YutfHQc5fmURa4Moj5qjV2shmqiY4qkac
FnvracOcEC0TEhAwRvxBJm8pwFpuzHJqSvMAM07Nk+g9GVWfhDEXZd+is+wdDAFj
U3EDRp31OzURAhHipPkfwqxsjgZX9nzHcsJwnbWsBd4MsbDUBmdwYxHasI7fvv/E
NkW8PE0m3KKRhmzFZt48BGmYmvfhVLdk5lIDYCerVfRnHWadA5YKdzW/1YvClrED
UyrkVRkuq0mAqbfr68xCzf9E5eEfO6MpD5rdiLHcPInhaJK7zP153kH95bkBJURH
Jp3q6F1RTCftJ17sVM0dSuCaDTLVML0NEGwClKgsuSstj8G+CvwUDRRleNWL42zS
Lx4Q8gvZD7w45GyDnmfxLq4V0UunLjVnpP3ggkbJnJ1tshy5vUW1Ifc3o4m94iJH
Wp3Sp0hfi7OymhMEdS+0OGWHlRkJxc86EpZeaxvk8yvFCtoCVdI/cw/Nr0eWjREQ
d6lDz4gyNtXjG6yc+NJEnzEDhrHfxxXvZJyE3+977Akx314W2ZcOexlCxloj5TIg
umB7qMGJf6OCpA4swCydF+PHoaN01sT1D6Vbsdi+DqfzGlYx4VxFh3I1Rl1f/NXX
a/BggmmbnljIYEVvVyhGZgCGab6uzLRdnBC6AQdhHT2QblYCDbZ19aXGKL+VLbDg
IgPxjBU/935Lju498W+LbOPtkfEWRz/Ax6ualaTHuZVKguvEAaIJFme2vOvqvOmd
8NTLCv6HhnS6wQ3uoVXE5/ep8c1PoTIuzMZEXNRxn/vw7si8ZGAbsVYPUzWdsgUx
4gQSCoM3NIQbJ9Sf+Idt8179eT0LvYN2OREqPe7ViRd4gXRK3DeEWckfQBeTbICi
92UGcTWV4TXCR+Kg9L6SH/GrxI8o8ZFjK7RB0zt1J/hSSKXJ7G5L+qCuXc9XRhFk
Yu6ycv2qLVFizylv6eyEPCH8sncK0spa3BbyDCSkFlNGYDKq3No4jnRKkpBkyKlR
lDzehaLAuYSGw2AjxsOO4h/7gVndbKbJBiatePIUQ2/8d/qOsqn7IhFGgeSaIt7x
aSvT68jxCRGim+1NDnmkUUp2f82oVn5LoMs3EfiZYzA8G5+79NSPPk9vC89gJvBO
tBGT/nWVXyp+n96yymi7vA==
`pragma protect end_protected
