`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DSfW+W74d8kY6OqghxTFmKXCfrT710+1j3ZXHkyeNkR8j8fYNLBdlwIoHDdUxqYn
ury2noyNIQjpIpkSGwrmWGlQpAhoKjjaBEUtcITfRGdGFaNSeTOCh5v0AeldYZ5X
Yz5BL3fWOpvc7rjv/AF7v5yAy2sA5XLtKgZuaRLMGxY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7088)
ovKRr1DYaO21kSF/Fqqq+Ba3XHS5eVwLsA6pugRIVkA1wZVwTuYq01nugSADMbEr
tZiyN5zc3VR2i0TU0+qBKwecc6F2J5Cqs7OfueFo3KXYy/Lhc+LpoxnV2SZdJ8hT
5D5eGvtKiR6zRaIk6vn/2+9n5/eCc+JVoAVc0W368mijgXUP6eW0BYQagc7u94sw
0NvaUB6jyPSn2YgW2dtG98wTNq2gd1tLgqs26rdVZszYMGEfwM2P1IQyRL/vSENe
xeHK567aAV9zenBzj75VifFTEPIzS4qlhxITHp3duyYGiUBBo5SX6PaVRmmi99VY
/dizY7StOw4RhqHCMyVdQ8PbFguLjIDr1gAk8IQNxmAc4CUgm1b/r4Iz409qmjcp
hY1o25n5iMN7T/BQOoLNqAN3KHldNSreCpUc1RK6+LlDqzxAhJAYc86xQ7c+4iqq
xECM04nPpWqjurlqwIFMz9fIe24Ze4Y4RRbWJCDY1wW4Phi8iycMAf8SA0Ne/eLY
uai0KqrgnEZ9d4owreFcHnLShdA1mSNAuf/tYCnQVaFCcFSajQPwxtPjeBzwOaEX
mTsq2AwGY4pX93EDZCq3/TOZ91xmpwxPLpcjTQ2bkiWjf9vh+NSA5ilJOjqbz3t8
9SiIGr+g2C/UsvfRS+RXpNycozzNThjnKcaaeiWadzRwI6F6siQeyNJr+tD4x+yz
b4p+YL7K6ghPAqa+WDwm93bkI8GuULn1+pRH+YJI1gN6voI+pQ60FgXlkI1GOXKt
FdYLwdP+QnIa6H6ZfEw2G7VLuz+oldLosCP3hccC5oyKBnXVED8HL49j0CXdQK9T
+fJBkUDQEqQRBSubeM8O4ToJTfBS9SDyHl4bnnAdsH53934YQT8pc9PYiuHcatx1
BIcBJ1Zhyg5zrWhEElvCPubz6bF0I3vpH9R7yYCaJ4dP0oAs430gdKai5Z2z353u
J/yFdqsUnZ1xLVRYWM+knVLevsWDapNLO3SpI15wACu4mnhFjXj9AamgXErL0Zgz
4U89sDjZbIYHwfXXXiPzvpysT6x5uvO5Sop0k3MapPH2WkevH6ELCNMEfLA8nhBM
wOCF3UK0XzLZUo2qmQfZZ7DcAyehB8MnheabN3SnpztSPjy713aUm8/KihLsa91t
Yk0IH77AVSLLkOapsXvUt2ASxf8vaY3rOgMH7D8Pn2DlHLUnYE1NGgZqXsq6SKDs
8v2rEmBv/NnMqJwVdT4qo4FKxI1a0xSixz+48+eLHRggaBehdFczECH5OHDpG7qH
xERZhLVvnErNpD2WDYJmBPCGLZseUItJobzKSJI0Abz/qPa5kNY1/fMKkV6iZqjF
a08sRtFenPx/RagqHZoMgg4H1ceh8GR08saHKsyj1YT4AYKXWGRj9Vxw29inKupP
KMRoZuWjH2I/E06ocTC2x8GoQbcRhAvryTgj4rGnnzC9lMzFRmopKE+HD1NEISpY
sMh3VbiA7XiQoNjMdHVTu2Y36eP6zV2xiHDfBcAu/20TMtrHAYIdjtbrwLOmeK8f
/49F4y52M6UarTmF9b+psVy9mISnJ6lgl5TcSFqhZ1ZyCNikuj1zCa6uM+7j+REo
3VW3rAT5J+84V7s0+PYK2wJ9rxZ79VYXiZjMR4r7twb05weJSV35PNVu1f8pxxp7
kOtdukcNjd/K6Ngxd+Bgzh25PkwXLIIWDLb+P3heVWz8rY+e1+FXePdZr3eI7vFa
VC+129nTk3xAz5krydbTcVqqgIDNvAJ0hqO+FBKd1OHVAOuT3d8JUYpapoZvZ1sF
S/rZUWLEQaSkw3YI29PILrtPhG0lc1Gz4fPc+XtSBz0KZZv6RCvmHOkiplm7LLHJ
aHvEe9aGS5CJgDnfR6S+ZPKgZ5hxWrU8rz+ay9mvFVWlzaJLozl8FxCjUCBIKU0W
Gz/FoXQlTnAOoOQXGmiyXpv5WbWMmSQq8resYiOBDhUvOhEs76z2UOaZvBKR33HZ
g674aGG/qj9W9BY0+yAKPuEbJaR2ryRqlHqHJ6KgxjwdhNFn+/+FR2NX4otNFlBl
jrB807EKLkFuF+7yjER4cxpJ5zlf5fLaC6TB4ni/z27U9fUcPwsTp5SlhvTXPKnv
/7cklCH8nQuPql0i+qDbrj2Z8M+0sZQ24Ng978SA7APH5A29dCjgTZGxLPC1DwSb
RgIsJAZKKvEYnlLxYYb5XWEZtqTUBBl/zOJAFRtu4nlQh63zxOsUHnHxs5Oo7jBJ
dk8+x403M8DIcGMqGG8WCaNAkyL4LDUUEvr0VQyQH6yeRHEfALXHe1VfdKM8Z5hm
JFoHmWQZ8i5d1xEFbm7UdMiHXhFfoWKGGNGfimopJ9r/DK6S1bBXtjGEsx9+n/p+
xzSvoTGFpoPjUZie8MmDokKEAHiprF7tQ+UEBJ9zQkqVuEIJVjb3P9U3Eb3/Z4Qq
EfKGJbmv9q+aOqCnfFeXKNn8HmzwjSQ9hzYxui0FSHy1UqqLPtT8ACPucoem8IoR
tLVU/pcIT9Nx6umioHBW2prHB6+Z0H3xlrANV4jJZpKNvv0gRMhNNuBuFBx3dhS7
u2lJOQgWHpEdyDTHn0KIhJQaxKzFsqJCJ1ZIwTChNw6ANM1zLohGTTfyqpJyeLnB
vD9B2DNsm9lxjLJc5iaKsmWgzaG3+tEg5ZbHrQt11KMgt9CnegkF4UVkrwfTxZZv
Y2NhIodwMQYG1UoZx7u+Un/wzIAOcIIT0T3bV9e9LZy+wULz35IQX8Ye2qKbfqmC
yXHHmoT2t79vIFC/cHRv7WABh/vic3q7/XRLe1GiFPDPGmRiQHvsKKDb+VrxJXzQ
eEswoEIVSyrqNEvs1GW0glEhiJF2y1N953eK461JsutVsXfxQG4E2+ZKdE5X8Gul
4C49+QtYuVHnkOK2d6sVOy1vVatiNN7KIwXwBr/iSn7zwvmVRPNTWfgaZe8/01eV
HEIFOXLgdsC5DPtJAEJbQMNo2xsVDydVQQNXc0UhaBar7aErSeimR9rnIkUTnM9C
6ge3sduMCGQGSVuNJtRMAMI80F8QJPBGWSRWxDhdxRSpeYz8AWaVMdrUyQSubeL5
Wd1eN0kqhsNmphs704iXzDf6mGkxEU0QGtg1bLFb8y/Is7KBxXpcGn99iozJIUPb
HCDQJHAOxM9xfzvqGLJu27Id1IIb3WNvCHAM+LojKOl8GRKMVLl3omIIGyy4T4lb
61CajTiN7GfFLLIg1w1oZYrSQbsDIOzGQhRjg/Ng+oZWsnJkZRwoZwZWCvIrUVgx
OCEXUgDmBGYOUYe8b3BSCPLOlSZ9EMTW2JpIll2Popz0urLXnw79n3/R48SgPmnL
RGyR5mZNT/pJruRkiqFf60QkUK/uuVk86U/JVA9Z0sEZX7/XaqpJCeGaOb/jixFW
SIrWFd6xSACcrmFvkKOkcPuGbcql3kj6EtVapWjGHxmMx92NwTZ8pgZMXyEQxq6J
008ceCLPGKlX+3HxF1AafghPBPVkOo9wK1rwfPHiZN9EnyFQ/biNkT95hyi/e3BJ
i3gxoKZYLVCdPYU6fLXN0Uy6TGE3muPTiAh5Lq8sPLx4Bgegui8BDTDSzzn+tsbV
8U7JHP3JTKKOSHeZ1ib1BoBXBtdXptwPBj6MqLayidvCBgK0HXTyjmmValFLFbPx
qx8oOFt50A0fvfVCKQkVDiCcIZp7bzMgPArijf/mnnXHXtolMuBiwQ49OjTXFxgz
w68os774X45vWil+iTzKNIK7JRuxeQuvXRSaS2lwO/KbDVODi/xJ9RIS39K0OpJc
WHG2uQlRC27a/0SSxiODgwHtjKcI8NNBKiGFW22afn6RhEd0gdgqgaQAk6jaW4R2
vTlDK7cYSG30gJZSvmlYcDIspY+PW+spQLP8THe2wF0EDO2tXuWYnPT3HOyCJdVa
c4Wg7VIRwuhVobQkKhGjFz2cBBdh5/fDJv58R0xuyP6IFWNwPo7hZERZLhoXzdWl
Kpv74kQpmIg0SEqdhVfQ756VzjPJu4JYD/bFifdk6wK+nI9Pt0mrbqzgnmxy36O/
5iNmbNktQpLgHAkBi6ZOWmzRfTBxYgpZmDXJEoqPGhBZFGUEpPJ1FoFoYPKHNd5q
ULcWYZoN/qQIxZRm7SXUFaXdoEtWRDbQsK9GS6NoyEE9aHn9K/4pDIjZkBUrhkba
Tf2ul7LHd3vtJpPRgEFdWfHCTlxy9tbTxlMc0CLqkQ8yDgvni4NuT5IUtjwzCoW/
UFHrzxcjWhpQIdFD8badWthGWx06aCEimHm3p1Gv3uiq4YIxYSXkIOF2Eh4pHpj3
HaicDblxHr9PFXUWlFz8YcdbTxSRgy+Ek0kZCCFwRvO65sKZgLAjtLQFWTl9fIo6
u61aFvSlYzLC2/2e6M+kSFxPi9FGknfDeYsOGcLGMlOAHVn3yJ2MeR7JIM8Paxud
r5SCHZMrD4+eoHHCYCyq5ehqYeiTZYZVKYdsJm0JLghpQepKLzwAmhbmPsIb3xY0
Zn2yb2XtJxzxb4axtVlGHUwd1kUnPivS9kjgktvPLLJamF9kxocjxzO1sWrnxkE8
1LJodc8RqgbwXEn17silFZsuwozYCHCJbwbrrHY1uEz5Szb+G5/zz3VQl8KgGX/z
wJ8L3DUwJzAhJl/Wr1blmp69YKLA/Y+BMxN7g2fDNqRzVc7QZnRTWVcH6Uln7dgB
zu4DG+3XzkkfT3uEUmP8EFu0wfA9jErNcZqueEs2QPFMTQkUQJS0i/sC3bWSOh2S
D8zsCYZs2tpUktRKXqZVx3Kr0yqp9KLtQ28IkMJTS8CAMdkLRdUZcwtxVIdjmV6U
PyyR4dCGrMlA8YQtGi/Q60nxnu7ZyguaUmB1DWRMaIBI/j5eQ6bWFDavP0OmdNTp
w8f2WC8Js6zShcz5pfMxy5wmTsTQkCYCIChzbcj4KQfOKjLa+YnI6f87Q6UI7iDW
+iJBklF4SvPD1/+stDDayj37gs0VeA9nFtIQh1BWRbs/a62Nhkam/FQ0tczOOIoj
S9rZ0uU9NANSo4xNoKFgi626JMnJj6B+MNx4DG4SiylLKb4kEdPY0VFKKS2/rjb8
tAd+MtvIc56CgZjjGVuP92p8YNSU/Xe0mkhw6KmUrM5T5qboE4s7a05aSD6qhhIM
kgxArAywR53dPGZAu5OQMu1PodkKx6XtrcqvWxV13iogAX61J0tw3wGerKreLBkQ
vgur1DooIJiAScNKWCmb7EHcKjaekfhtnMDIrwnlVGeN5QweXNZcuOtRSdVYSlE8
sa+tECvi1elTHCiaGcXzpp1iqAyJwh4kdKa8ajPk2RCDk3lzUomphQrwzGwqtoBO
mBOyxm/FhhnSpSY7GBx9IrZGkIjgrOAQGBJRQO91gS18WIKRr2HH9XkEIazOgAm1
GVj0jWuZX0Se3A7n7KLzIt94QmbvKsAHB6+3RA2KbriX8jicBJIxAXUmIUgfgy9h
aYJaH6DAH6wI6PvXc5gMBkFAavbMntitGMpG5EtrYI40tXISKicK9X6ZpkJxTtA8
Mrg+zWmz16c9dH+GH7eAXxL9GtXx6ccsw0ycq+Sr4l85Ffy7gkGkvBPxOFUC0ZmZ
cE1tXhHyfh8x9byKsjhsDD8g1qoPAe3IXJz7AN1/rRXNhtWIhjFVLeBfcxSjA7TU
+ZesyokipwypiaJYctfhavttp95EwMiddSGsObnYERuT62f2Cr7YLwLD8yltwj+l
Nu0W0CaLY1gNg6dzVfQ54F4dnGcuv7S4GOQP4/cTWx31xeOeueCW5jDXiTfyhfW7
DsmRsB8gECza78ebHoD/Oei6MFXKEOwpBDA7qPNz0g/YH6OvzA8fg7UEZs8sc9Mt
vXRhxe147xDzQeMyZnKk7pzczysqAEZ+cGl0WyevhU3204QMUlt0VgwC+MEkGvO1
rsl8I5RilnyDSiK8574P9KSJ2Rvx1Rjx9LaB8qAJ+Rtof3j6U1pMpKrImFYf9hx9
PCwFjr7cUvaf1x9eKk4GBxCfT6ZIUwFwdOz+F7UbQzJ9p9UfAdCh/vi1NnDid4YJ
Mxezzl7aA431PUkc86dMDp1FLy7EahGP0Jn/Sw9cJ2dvtKW8GnnsUmjIB+YIUP4f
h+tuelHgemVYR/oeFR6Nu2e27brOpSXx0K51PGsuGn52k9jsgIGWoZgT6BylsZCz
QdvJn+gtnATleiYA2oZMkqSNgMnagQrQkT1raWRkSOax77JaTBmX4+/P9x4g1kcD
ZwdbWlqgNP+W4AMN93f0aIY/VPE6JzGHwFPoobyRNNkVTJ+LvCjpND2v5dYbB23Z
W4udfarj/tYeam0TELSWF4BZ1AQgfvYZiE3/5OTFUaJg1RrlWXv8gPTzI1tf8pxS
wnI6G0Ufpd1kBrX1R3bWWG/vHiJkRcORrGUK5GIYnK48iBSxb3TImFvZedXaxDo1
yqZ8EZGdktnlJRH+cVHYwcfO13Dj0UAQDqtTr9Mwit8xlQGre2IOhPHXi+aGZMDv
dX8O2nyLLcbNoTHxGI66VaI2NDn+DSZCuv2e75HZdatJTlUWJUblP4oXvEmKAK9a
jXj3+RzHFxW9QMyRub+Up73HKJ6v7dzRX/t6k3QUxuYTrmEk6K8SluDgMWhyW8Tc
zi01AzZkmSltpjC2x+ZzOijURsNODVRTGknH2FveeKD0tFhbtVcJSGoY38GKDjZt
cFq0ZT84MJ0PUHXSNjBkIpoPe25+KYpfD9ns7q2QWGVuLmiN517Y0p/P39eOH06P
Kuf4sq0WUK5JSKvgF6CqUR3BCvGnYhndzaqxxdfXERPCmC9rM4rTqjliFWyqJe0Z
XH90KbGcxAvo3Fu1afZLh5UQ/uGf8P9d9x4wtyl3FPa5C79GC9TfCSI1/l86xS2U
kaCWrURl4P5SSWdeaLIhUVMaW9zVPEZ6sBwKBKn10I87J58IXpKfQkK1YcijbIw3
2OzdG2Q3YN60f7OtUJwjUkUfeFXldwtTFGuCm/vwUaOSYalrVw5R5nefhUAM9/I5
O/O4bQupKsLtyNdGSen+MZWNGGD3B2TspyaQ2w1paWLaCBr1gjdB0PSPPb+wCKJg
bhthpyinn02f9QC6Zf5VQUhJ88qWShN9VDg0/wfvaKvL78W7uuDJBHMneCOgvc3I
kpB8k+IxfshePzd/Snx9IX5UZTtIdy3nE8ZWdmZDjV5X46LBgowriYpBCu782Ql0
SSpF1xRhgxKEvdBSrVxIuXVKWnRTNU8VYMK6PMR0G5ZuAVH4diDvTEl5mTra+J23
MoByNChDGntk0NgP6Idm+WhDmQ3fnEWGwE/7ykc+V4JZZBo7YLGwe08HowfrR9NS
fmqNdyM4NADLU3+rd0Gk56i1XuHh86quwewZj/6p7WZW2V1sYCeHs8qmwwpVVoJN
Y2QipTEMb99zmYvEjnhbLVIkpegPw7vqymmVw9nuQK+Igm3BaQp2amlTcounR7fX
soXjEvMuinV/svAjUbf4rC86+3WgMW11hdh70LXzY7ynmFJjVKXBH2ZDsWfOcp9R
sfxEEQqlqOD/smuvosS2lTc2MN0XflxLZQo16uBxsVd/xYGTevlX/9tOG1M3rI/w
BeqAJEWmuyDvRc8zT6Hss6swHXJYgn+w0SqSvoUO/h6zgMTSq98VOHH/2SWZvRZw
0lDAehHBN0C3o/bllvtbbctutTwGkQQPYVar2XpQwGaQNf9/ZeGTx/q7FjuqFUDk
g4bqWVAo4eNg474x4jpMVlhUve5mBQc2xo7h967S7KKHX8WGdBYmUuSFjOJimxws
KzfAPj0vcnqahY/YXm1Sqf2q8pZ61Twf0wvLJRRoAQCv8pcK4hNuxdTuyV2GfMd/
opNPmWeVlip6+R44F0Qp6g2CSskzUbKg6fcCqbCskwr1ymxwg+3Iq0O0y5+xfIjw
LiBFrD5KxZVDtokI8YVa+ZEZj0PdXzCgBuO+tWxRd9a6DRzr5ZILcu12537YhfF0
0cQCYwEVD+D05afRitKODSqj6SPcKfrnx4QBWq364Y4legCv9DK8vyDxc441Ve46
Ui47rJLmKKOveWWG/00J3g/HL2nu1WiDq7hqKnebC08GWQVmjHCUJlR8xAjAAPpC
Abf/9BkKE0YwelBJjV57jx85kCXyY/pF+/F55UmzpT9JvdoYJIGmBnvFsgsnwcXY
K62Hdcpd1POrQwTh7LwXa0GRyBr4TP17PENn1dAZWUJLkBPup7a0Bbd0Jh8vobFK
uUfi9tlw0/deoU5aawxIQNUnAI8ORLr0MiBnxx59rf1aVOTCZSZNaUics0Frk1mi
w/liYzS4+89WtsXi7aTYy91C6qWspUydHROV290MEfH85p97poJiyqM6W8rFHgQB
w0C1kpAdrydZLoeUVh3lGyIJjHBdZszMGAfdx6Yu4o6uEDA3TYC6hsh4GxN/Gb2x
bzzB9CvWQlfzW7XT+rfO9SpV4lfW/ROQOIc5eqcgz46pQonyEBzzWmNzUkv0Ro+W
SDEI4mieMKG5fux7tc+2ao0C6ZZgYex/cvOsf1A4HiV88kU2rLahXBD1mwlNV/Qk
5ffZaPaDCwIe19PsBKvF0ZzyIq5HHvIwROxsOC71ZBnXo1sN5QVvQplu8MyowYQ5
yJxcot/9eJrAs7TLvLnEmx2e4A5sSNkbKKUHXWEG//Vgs/ALNlu6yMNb+fjLbxX/
kfBgp7wR8UCyOvSA4RDxgXG6xpaFnjpJRu37PHLRYnne2Ryh128g7lptsB9+G5pe
gbPC8vdNgNmArg68C+YmjjjLQBXFhsp1VrQGzR2aOVG5bL3LI+TtkXfH8B4bDrtl
QCXM+tsm+pZy0LFzKFt655McPQq7WQGmj95hDN1Pp0L1+yU1dJk82+uhwdFw8wRt
PiLlktY47rE9eOO7Zx4FgaFrhzaqzngEc6xYlG8iZmBnrEbKEwCELqO8pf530114
3hqsHqhZ6n8GKP8waOeN2aICBikJAKSUn48NYtUygPbnsnHztnMXi2wkpyZr3bDE
MmaSsM+qRrEBYagAtARrTesnv0lD0FaQcYYOZSUtXpBcMzuoXLt4Ar+y7NHOBY4c
XR9FrYSYyooHl5YsD4afGCZWa0PR5V16ycq5aKb1mBtvDIZ4qv54FzQSh/tCtYKk
ynoUoaskBM/kTdTY/9HYTiRGYKG+lRihBxPGUNCLmSJfWwhJmimq6OIuyY3s4w+B
QZKx/YM2Zb8btzNV/XSb2Mngnfq0JD5ecLZ4kOYqnp4q08P6jYN1InKeFF73kIy3
4Z3NiFpOdZDhpWWOIZH1Ctq4QcrPXKWOkQ20Ks1JIQyAPXK6h7hPP6PZRwmroTCP
aYmgNUyZ3NbS5tMuGmis35OoL0FTtiSGC/zSBmSeHUdYovAR1igmD2kBdUyCYLe6
kbVyhG3Ew9HLCvuvw4trbA04IEAt5TFbUHupgZlSyODGWQXdx0zf9WO7S5NH6Zqd
EPiXrja6nUdqkXr4td7/hJiT4oXCcmHebcjt2BET5ao=
`pragma protect end_protected
