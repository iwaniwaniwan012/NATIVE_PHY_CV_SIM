-- Trans_Native_Phy.vhd

-- Generated using ACDS version 21.1 842

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Trans_Native_Phy is
	port (
		pll_powerdown           : in  std_logic_vector(0 downto 0)   := (others => '0'); --           pll_powerdown.pll_powerdown
		tx_analogreset          : in  std_logic_vector(0 downto 0)   := (others => '0'); --          tx_analogreset.tx_analogreset
		tx_digitalreset         : in  std_logic_vector(0 downto 0)   := (others => '0'); --         tx_digitalreset.tx_digitalreset
		tx_pll_refclk           : in  std_logic_vector(0 downto 0)   := (others => '0'); --           tx_pll_refclk.tx_pll_refclk
		tx_serial_data          : out std_logic_vector(0 downto 0);                      --          tx_serial_data.tx_serial_data
		pll_locked              : out std_logic_vector(0 downto 0);                      --              pll_locked.pll_locked
		rx_analogreset          : in  std_logic_vector(0 downto 0)   := (others => '0'); --          rx_analogreset.rx_analogreset
		rx_digitalreset         : in  std_logic_vector(0 downto 0)   := (others => '0'); --         rx_digitalreset.rx_digitalreset
		rx_cdr_refclk           : in  std_logic_vector(0 downto 0)   := (others => '0'); --           rx_cdr_refclk.rx_cdr_refclk
		rx_serial_data          : in  std_logic_vector(0 downto 0)   := (others => '0'); --          rx_serial_data.rx_serial_data
		rx_is_lockedtoref       : out std_logic_vector(0 downto 0);                      --       rx_is_lockedtoref.rx_is_lockedtoref
		rx_is_lockedtodata      : out std_logic_vector(0 downto 0);                      --      rx_is_lockedtodata.rx_is_lockedtodata
		tx_std_coreclkin        : in  std_logic_vector(0 downto 0)   := (others => '0'); --        tx_std_coreclkin.tx_std_coreclkin
		rx_std_coreclkin        : in  std_logic_vector(0 downto 0)   := (others => '0'); --        rx_std_coreclkin.rx_std_coreclkin
		tx_std_clkout           : out std_logic_vector(0 downto 0);                      --           tx_std_clkout.tx_std_clkout
		rx_std_clkout           : out std_logic_vector(0 downto 0);                      --           rx_std_clkout.rx_std_clkout
		tx_cal_busy             : out std_logic_vector(0 downto 0);                      --             tx_cal_busy.tx_cal_busy
		rx_cal_busy             : out std_logic_vector(0 downto 0);                      --             rx_cal_busy.rx_cal_busy
		reconfig_to_xcvr        : in  std_logic_vector(139 downto 0) := (others => '0'); --        reconfig_to_xcvr.reconfig_to_xcvr
		reconfig_from_xcvr      : out std_logic_vector(91 downto 0);                     --      reconfig_from_xcvr.reconfig_from_xcvr
		tx_parallel_data        : in  std_logic_vector(19 downto 0)  := (others => '0'); --        tx_parallel_data.tx_parallel_data
		unused_tx_parallel_data : in  std_logic_vector(23 downto 0)  := (others => '0'); -- unused_tx_parallel_data.unused_tx_parallel_data
		rx_parallel_data        : out std_logic_vector(19 downto 0);                     --        rx_parallel_data.rx_parallel_data
		unused_rx_parallel_data : out std_logic_vector(43 downto 0)                      -- unused_rx_parallel_data.unused_rx_parallel_data
	);
end entity Trans_Native_Phy;

architecture rtl of Trans_Native_Phy is
	component altera_xcvr_native_av is
		generic (
			tx_enable                       : integer := 1;
			rx_enable                       : integer := 1;
			enable_std                      : integer := 1;
			data_path_select                : string  := "standard";
			channels                        : integer := 1;
			bonded_mode                     : string  := "non_bonded";
			data_rate                       : string  := "";
			pma_width                       : integer := 10;
			tx_pma_clk_div                  : integer := 1;
			pll_reconfig_enable             : integer := 0;
			pll_external_enable             : integer := 0;
			pll_data_rate                   : string  := "0 Mbps";
			pll_type                        : string  := "CMU";
			pma_bonding_mode                : string  := "x1";
			plls                            : integer := 1;
			pll_select                      : integer := 0;
			pll_refclk_cnt                  : integer := 1;
			pll_refclk_select               : string  := "0";
			pll_refclk_freq                 : string  := "125.0 MHz";
			pll_feedback_path               : string  := "internal";
			cdr_reconfig_enable             : integer := 0;
			cdr_refclk_cnt                  : integer := 1;
			cdr_refclk_select               : integer := 0;
			cdr_refclk_freq                 : string  := "";
			rx_ppm_detect_threshold         : string  := "1000";
			rx_clkslip_enable               : integer := 0;
			std_protocol_hint               : string  := "basic";
			std_pcs_pma_width               : integer := 10;
			std_low_latency_bypass_enable   : integer := 0;
			std_tx_pcfifo_mode              : string  := "low_latency";
			std_rx_pcfifo_mode              : string  := "low_latency";
			std_rx_byte_order_enable        : integer := 0;
			std_rx_byte_order_mode          : string  := "manual";
			std_rx_byte_order_width         : integer := 10;
			std_rx_byte_order_symbol_count  : integer := 1;
			std_rx_byte_order_pattern       : string  := "0";
			std_rx_byte_order_pad           : string  := "0";
			std_tx_byte_ser_enable          : integer := 0;
			std_rx_byte_deser_enable        : integer := 0;
			std_tx_8b10b_enable             : integer := 0;
			std_tx_8b10b_disp_ctrl_enable   : integer := 0;
			std_rx_8b10b_enable             : integer := 0;
			std_rx_rmfifo_enable            : integer := 0;
			std_rx_rmfifo_pattern_p         : string  := "00000";
			std_rx_rmfifo_pattern_n         : string  := "00000";
			std_tx_bitslip_enable           : integer := 0;
			std_rx_word_aligner_mode        : string  := "bit_slip";
			std_rx_word_aligner_pattern_len : integer := 7;
			std_rx_word_aligner_pattern     : string  := "0000000000";
			std_rx_word_aligner_rknumber    : integer := 3;
			std_rx_word_aligner_renumber    : integer := 3;
			std_rx_word_aligner_rgnumber    : integer := 3;
			std_rx_run_length_val           : integer := 31;
			std_tx_bitrev_enable            : integer := 0;
			std_rx_bitrev_enable            : integer := 0;
			std_tx_byterev_enable           : integer := 0;
			std_rx_byterev_enable           : integer := 0;
			std_tx_polinv_enable            : integer := 0;
			std_rx_polinv_enable            : integer := 0
		);
		port (
			pll_powerdown             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- pll_powerdown
			tx_analogreset            : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- tx_analogreset
			tx_digitalreset           : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- tx_digitalreset
			tx_pll_refclk             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- tx_pll_refclk
			tx_serial_data            : out std_logic_vector(0 downto 0);                      -- tx_serial_data
			pll_locked                : out std_logic_vector(0 downto 0);                      -- pll_locked
			rx_analogreset            : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- rx_analogreset
			rx_digitalreset           : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- rx_digitalreset
			rx_cdr_refclk             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- rx_cdr_refclk
			rx_serial_data            : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- rx_serial_data
			rx_is_lockedtoref         : out std_logic_vector(0 downto 0);                      -- rx_is_lockedtoref
			rx_is_lockedtodata        : out std_logic_vector(0 downto 0);                      -- rx_is_lockedtodata
			tx_std_coreclkin          : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- tx_std_coreclkin
			rx_std_coreclkin          : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- rx_std_coreclkin
			tx_std_clkout             : out std_logic_vector(0 downto 0);                      -- tx_std_clkout
			rx_std_clkout             : out std_logic_vector(0 downto 0);                      -- rx_std_clkout
			tx_cal_busy               : out std_logic_vector(0 downto 0);                      -- tx_cal_busy
			rx_cal_busy               : out std_logic_vector(0 downto 0);                      -- rx_cal_busy
			reconfig_to_xcvr          : in  std_logic_vector(139 downto 0) := (others => 'X'); -- reconfig_to_xcvr
			reconfig_from_xcvr        : out std_logic_vector(91 downto 0);                     -- reconfig_from_xcvr
			tx_parallel_data          : in  std_logic_vector(43 downto 0)  := (others => 'X'); -- unused_tx_parallel_data
			rx_parallel_data          : out std_logic_vector(63 downto 0);                     -- unused_rx_parallel_data
			tx_pma_clkout             : out std_logic_vector(0 downto 0);                      -- tx_pma_clkout
			tx_pma_parallel_data      : in  std_logic_vector(79 downto 0)  := (others => 'X'); -- tx_pma_parallel_data
			ext_pll_clk               : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- ext_pll_clk
			rx_pma_clkout             : out std_logic_vector(0 downto 0);                      -- rx_pma_clkout
			rx_pma_parallel_data      : out std_logic_vector(79 downto 0);                     -- rx_pma_parallel_data
			rx_clkslip                : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- rx_clkslip
			rx_clklow                 : out std_logic_vector(0 downto 0);                      -- rx_clklow
			rx_fref                   : out std_logic_vector(0 downto 0);                      -- rx_fref
			rx_set_locktodata         : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- rx_set_locktodata
			rx_set_locktoref          : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- rx_set_locktoref
			rx_seriallpbken           : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- rx_seriallpbken
			rx_signaldetect           : out std_logic_vector(0 downto 0);                      -- rx_signaldetect
			rx_std_prbs_done          : out std_logic_vector(0 downto 0);                      -- rx_std_prbs_done
			rx_std_prbs_err           : out std_logic_vector(0 downto 0);                      -- rx_std_prbs_err
			tx_std_pcfifo_full        : out std_logic_vector(0 downto 0);                      -- tx_std_pcfifo_full
			tx_std_pcfifo_empty       : out std_logic_vector(0 downto 0);                      -- tx_std_pcfifo_empty
			rx_std_pcfifo_full        : out std_logic_vector(0 downto 0);                      -- rx_std_pcfifo_full
			rx_std_pcfifo_empty       : out std_logic_vector(0 downto 0);                      -- rx_std_pcfifo_empty
			rx_std_byteorder_ena      : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- rx_std_byteorder_ena
			rx_std_byteorder_flag     : out std_logic_vector(0 downto 0);                      -- rx_std_byteorder_flag
			rx_std_rmfifo_full        : out std_logic_vector(0 downto 0);                      -- rx_std_rmfifo_full
			rx_std_rmfifo_empty       : out std_logic_vector(0 downto 0);                      -- rx_std_rmfifo_empty
			rx_std_wa_patternalign    : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- rx_std_wa_patternalign
			rx_std_wa_a1a2size        : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- rx_std_wa_a1a2size
			tx_std_bitslipboundarysel : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- tx_std_bitslipboundarysel
			rx_std_bitslipboundarysel : out std_logic_vector(4 downto 0);                      -- rx_std_bitslipboundarysel
			rx_std_bitslip            : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- rx_std_bitslip
			rx_std_runlength_err      : out std_logic_vector(0 downto 0);                      -- rx_std_runlength_err
			rx_std_bitrev_ena         : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- rx_std_bitrev_ena
			rx_std_byterev_ena        : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- rx_std_byterev_ena
			tx_std_polinv             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- tx_std_polinv
			rx_std_polinv             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- rx_std_polinv
			tx_std_elecidle           : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- tx_std_elecidle
			rx_std_signaldetect       : out std_logic_vector(0 downto 0)                       -- rx_std_signaldetect
		);
	end component altera_xcvr_native_av;

	signal trans_native_phy_inst_rx_parallel_data : std_logic_vector(63 downto 0); -- port fragment

begin

	trans_native_phy_inst : component altera_xcvr_native_av
		generic map (
			tx_enable                       => 1,
			rx_enable                       => 1,
			enable_std                      => 1,
			data_path_select                => "standard",
			channels                        => 1,
			bonded_mode                     => "non_bonded",
			data_rate                       => "1250 Mbps",
			pma_width                       => 20,
			tx_pma_clk_div                  => 1,
			pll_reconfig_enable             => 1,
			pll_external_enable             => 0,
			pll_data_rate                   => "1250 Mbps",
			pll_type                        => "CMU",
			pma_bonding_mode                => "x1",
			plls                            => 1,
			pll_select                      => 0,
			pll_refclk_cnt                  => 1,
			pll_refclk_select               => "0",
			pll_refclk_freq                 => "125.0 MHz",
			pll_feedback_path               => "internal",
			cdr_reconfig_enable             => 1,
			cdr_refclk_cnt                  => 1,
			cdr_refclk_select               => 0,
			cdr_refclk_freq                 => "125.0 MHz",
			rx_ppm_detect_threshold         => "1000",
			rx_clkslip_enable               => 0,
			std_protocol_hint               => "basic",
			std_pcs_pma_width               => 20,
			std_low_latency_bypass_enable   => 1,
			std_tx_pcfifo_mode              => "low_latency",
			std_rx_pcfifo_mode              => "low_latency",
			std_rx_byte_order_enable        => 0,
			std_rx_byte_order_mode          => "manual",
			std_rx_byte_order_width         => 10,
			std_rx_byte_order_symbol_count  => 1,
			std_rx_byte_order_pattern       => "0",
			std_rx_byte_order_pad           => "0",
			std_tx_byte_ser_enable          => 0,
			std_rx_byte_deser_enable        => 0,
			std_tx_8b10b_enable             => 0,
			std_tx_8b10b_disp_ctrl_enable   => 0,
			std_rx_8b10b_enable             => 0,
			std_rx_rmfifo_enable            => 0,
			std_rx_rmfifo_pattern_p         => "00000",
			std_rx_rmfifo_pattern_n         => "00000",
			std_tx_bitslip_enable           => 0,
			std_rx_word_aligner_mode        => "bit_slip",
			std_rx_word_aligner_pattern_len => 7,
			std_rx_word_aligner_pattern     => "0000000000",
			std_rx_word_aligner_rknumber    => 3,
			std_rx_word_aligner_renumber    => 3,
			std_rx_word_aligner_rgnumber    => 3,
			std_rx_run_length_val           => 31,
			std_tx_bitrev_enable            => 0,
			std_rx_bitrev_enable            => 0,
			std_tx_byterev_enable           => 0,
			std_rx_byterev_enable           => 0,
			std_tx_polinv_enable            => 0,
			std_rx_polinv_enable            => 0
		)
		port map (
			pll_powerdown             => pll_powerdown,                                                                      --      pll_powerdown.pll_powerdown
			tx_analogreset            => tx_analogreset,                                                                     --     tx_analogreset.tx_analogreset
			tx_digitalreset           => tx_digitalreset,                                                                    --    tx_digitalreset.tx_digitalreset
			tx_pll_refclk             => tx_pll_refclk,                                                                      --      tx_pll_refclk.tx_pll_refclk
			tx_serial_data            => tx_serial_data,                                                                     --     tx_serial_data.tx_serial_data
			pll_locked                => pll_locked,                                                                         --         pll_locked.pll_locked
			rx_analogreset            => rx_analogreset,                                                                     --     rx_analogreset.rx_analogreset
			rx_digitalreset           => rx_digitalreset,                                                                    --    rx_digitalreset.rx_digitalreset
			rx_cdr_refclk             => rx_cdr_refclk,                                                                      --      rx_cdr_refclk.rx_cdr_refclk
			rx_serial_data            => rx_serial_data,                                                                     --     rx_serial_data.rx_serial_data
			rx_is_lockedtoref         => rx_is_lockedtoref,                                                                  --  rx_is_lockedtoref.rx_is_lockedtoref
			rx_is_lockedtodata        => rx_is_lockedtodata,                                                                 -- rx_is_lockedtodata.rx_is_lockedtodata
			tx_std_coreclkin          => tx_std_coreclkin,                                                                   --   tx_std_coreclkin.tx_std_coreclkin
			rx_std_coreclkin          => rx_std_coreclkin,                                                                   --   rx_std_coreclkin.rx_std_coreclkin
			tx_std_clkout             => tx_std_clkout,                                                                      --      tx_std_clkout.tx_std_clkout
			rx_std_clkout             => rx_std_clkout,                                                                      --      rx_std_clkout.rx_std_clkout
			tx_cal_busy               => tx_cal_busy,                                                                        --        tx_cal_busy.tx_cal_busy
			rx_cal_busy               => rx_cal_busy,                                                                        --        rx_cal_busy.rx_cal_busy
			reconfig_to_xcvr          => reconfig_to_xcvr,                                                                   --   reconfig_to_xcvr.reconfig_to_xcvr
			reconfig_from_xcvr        => reconfig_from_xcvr,                                                                 -- reconfig_from_xcvr.reconfig_from_xcvr
			tx_parallel_data(0)       => tx_parallel_data(0),                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(1)       => tx_parallel_data(1),                                                                --                   .tx_parallel_data
			tx_parallel_data(2)       => tx_parallel_data(2),                                                                --                   .tx_parallel_data
			tx_parallel_data(3)       => tx_parallel_data(3),                                                                --                   .tx_parallel_data
			tx_parallel_data(4)       => tx_parallel_data(4),                                                                --                   .tx_parallel_data
			tx_parallel_data(5)       => tx_parallel_data(5),                                                                --                   .tx_parallel_data
			tx_parallel_data(6)       => tx_parallel_data(6),                                                                --                   .tx_parallel_data
			tx_parallel_data(7)       => tx_parallel_data(7),                                                                --                   .tx_parallel_data
			tx_parallel_data(8)       => tx_parallel_data(8),                                                                --                   .tx_parallel_data
			tx_parallel_data(9)       => tx_parallel_data(9),                                                                --                   .tx_parallel_data
			tx_parallel_data(10)      => unused_tx_parallel_data(0),                                                         --                   .tx_parallel_data
			tx_parallel_data(11)      => tx_parallel_data(10),                                                               --                   .tx_parallel_data
			tx_parallel_data(12)      => tx_parallel_data(11),                                                               --                   .tx_parallel_data
			tx_parallel_data(13)      => tx_parallel_data(12),                                                               --                   .tx_parallel_data
			tx_parallel_data(14)      => tx_parallel_data(13),                                                               --                   .tx_parallel_data
			tx_parallel_data(15)      => tx_parallel_data(14),                                                               --                   .tx_parallel_data
			tx_parallel_data(16)      => tx_parallel_data(15),                                                               --                   .tx_parallel_data
			tx_parallel_data(17)      => tx_parallel_data(16),                                                               --                   .tx_parallel_data
			tx_parallel_data(18)      => tx_parallel_data(17),                                                               --                   .tx_parallel_data
			tx_parallel_data(19)      => tx_parallel_data(18),                                                               --                   .tx_parallel_data
			tx_parallel_data(20)      => tx_parallel_data(19),                                                               --                   .tx_parallel_data
			tx_parallel_data(21)      => unused_tx_parallel_data(1),                                                         --                   .tx_parallel_data
			tx_parallel_data(22)      => unused_tx_parallel_data(2),                                                         --                   .tx_parallel_data
			tx_parallel_data(23)      => unused_tx_parallel_data(3),                                                         --                   .tx_parallel_data
			tx_parallel_data(24)      => unused_tx_parallel_data(4),                                                         --                   .tx_parallel_data
			tx_parallel_data(25)      => unused_tx_parallel_data(5),                                                         --                   .tx_parallel_data
			tx_parallel_data(26)      => unused_tx_parallel_data(6),                                                         --                   .tx_parallel_data
			tx_parallel_data(27)      => unused_tx_parallel_data(7),                                                         --                   .tx_parallel_data
			tx_parallel_data(28)      => unused_tx_parallel_data(8),                                                         --                   .tx_parallel_data
			tx_parallel_data(29)      => unused_tx_parallel_data(9),                                                         --                   .tx_parallel_data
			tx_parallel_data(30)      => unused_tx_parallel_data(10),                                                        --                   .tx_parallel_data
			tx_parallel_data(31)      => unused_tx_parallel_data(11),                                                        --                   .tx_parallel_data
			tx_parallel_data(32)      => unused_tx_parallel_data(12),                                                        --                   .tx_parallel_data
			tx_parallel_data(33)      => unused_tx_parallel_data(13),                                                        --                   .tx_parallel_data
			tx_parallel_data(34)      => unused_tx_parallel_data(14),                                                        --                   .tx_parallel_data
			tx_parallel_data(35)      => unused_tx_parallel_data(15),                                                        --                   .tx_parallel_data
			tx_parallel_data(36)      => unused_tx_parallel_data(16),                                                        --                   .tx_parallel_data
			tx_parallel_data(37)      => unused_tx_parallel_data(17),                                                        --                   .tx_parallel_data
			tx_parallel_data(38)      => unused_tx_parallel_data(18),                                                        --                   .tx_parallel_data
			tx_parallel_data(39)      => unused_tx_parallel_data(19),                                                        --                   .tx_parallel_data
			tx_parallel_data(40)      => unused_tx_parallel_data(20),                                                        --                   .tx_parallel_data
			tx_parallel_data(41)      => unused_tx_parallel_data(21),                                                        --                   .tx_parallel_data
			tx_parallel_data(42)      => unused_tx_parallel_data(22),                                                        --                   .tx_parallel_data
			tx_parallel_data(43)      => unused_tx_parallel_data(23),                                                        --                   .tx_parallel_data
			rx_parallel_data(0)       => trans_native_phy_inst_rx_parallel_data(0),                                          --   rx_parallel_data.rx_parallel_data
			rx_parallel_data(1)       => trans_native_phy_inst_rx_parallel_data(1),                                          --                   .rx_parallel_data
			rx_parallel_data(2)       => trans_native_phy_inst_rx_parallel_data(2),                                          --                   .rx_parallel_data
			rx_parallel_data(3)       => trans_native_phy_inst_rx_parallel_data(3),                                          --                   .rx_parallel_data
			rx_parallel_data(4)       => trans_native_phy_inst_rx_parallel_data(4),                                          --                   .rx_parallel_data
			rx_parallel_data(5)       => trans_native_phy_inst_rx_parallel_data(5),                                          --                   .rx_parallel_data
			rx_parallel_data(6)       => trans_native_phy_inst_rx_parallel_data(6),                                          --                   .rx_parallel_data
			rx_parallel_data(7)       => trans_native_phy_inst_rx_parallel_data(7),                                          --                   .rx_parallel_data
			rx_parallel_data(8)       => trans_native_phy_inst_rx_parallel_data(8),                                          --                   .rx_parallel_data
			rx_parallel_data(9)       => trans_native_phy_inst_rx_parallel_data(9),                                          --                   .rx_parallel_data
			rx_parallel_data(10)      => trans_native_phy_inst_rx_parallel_data(10),                                         --                   .rx_parallel_data
			rx_parallel_data(11)      => trans_native_phy_inst_rx_parallel_data(11),                                         --                   .rx_parallel_data
			rx_parallel_data(12)      => trans_native_phy_inst_rx_parallel_data(12),                                         --                   .rx_parallel_data
			rx_parallel_data(13)      => trans_native_phy_inst_rx_parallel_data(13),                                         --                   .rx_parallel_data
			rx_parallel_data(14)      => trans_native_phy_inst_rx_parallel_data(14),                                         --                   .rx_parallel_data
			rx_parallel_data(15)      => trans_native_phy_inst_rx_parallel_data(15),                                         --                   .rx_parallel_data
			rx_parallel_data(16)      => trans_native_phy_inst_rx_parallel_data(16),                                         --                   .rx_parallel_data
			rx_parallel_data(17)      => trans_native_phy_inst_rx_parallel_data(17),                                         --                   .rx_parallel_data
			rx_parallel_data(18)      => trans_native_phy_inst_rx_parallel_data(18),                                         --                   .rx_parallel_data
			rx_parallel_data(19)      => trans_native_phy_inst_rx_parallel_data(19),                                         --                   .rx_parallel_data
			rx_parallel_data(20)      => trans_native_phy_inst_rx_parallel_data(20),                                         --                   .rx_parallel_data
			rx_parallel_data(21)      => trans_native_phy_inst_rx_parallel_data(21),                                         --                   .rx_parallel_data
			rx_parallel_data(22)      => trans_native_phy_inst_rx_parallel_data(22),                                         --                   .rx_parallel_data
			rx_parallel_data(23)      => trans_native_phy_inst_rx_parallel_data(23),                                         --                   .rx_parallel_data
			rx_parallel_data(24)      => trans_native_phy_inst_rx_parallel_data(24),                                         --                   .rx_parallel_data
			rx_parallel_data(25)      => trans_native_phy_inst_rx_parallel_data(25),                                         --                   .rx_parallel_data
			rx_parallel_data(26)      => trans_native_phy_inst_rx_parallel_data(26),                                         --                   .rx_parallel_data
			rx_parallel_data(27)      => trans_native_phy_inst_rx_parallel_data(27),                                         --                   .rx_parallel_data
			rx_parallel_data(28)      => trans_native_phy_inst_rx_parallel_data(28),                                         --                   .rx_parallel_data
			rx_parallel_data(29)      => trans_native_phy_inst_rx_parallel_data(29),                                         --                   .rx_parallel_data
			rx_parallel_data(30)      => trans_native_phy_inst_rx_parallel_data(30),                                         --                   .rx_parallel_data
			rx_parallel_data(31)      => trans_native_phy_inst_rx_parallel_data(31),                                         --                   .rx_parallel_data
			rx_parallel_data(32)      => trans_native_phy_inst_rx_parallel_data(32),                                         --                   .rx_parallel_data
			rx_parallel_data(33)      => trans_native_phy_inst_rx_parallel_data(33),                                         --                   .rx_parallel_data
			rx_parallel_data(34)      => trans_native_phy_inst_rx_parallel_data(34),                                         --                   .rx_parallel_data
			rx_parallel_data(35)      => trans_native_phy_inst_rx_parallel_data(35),                                         --                   .rx_parallel_data
			rx_parallel_data(36)      => trans_native_phy_inst_rx_parallel_data(36),                                         --                   .rx_parallel_data
			rx_parallel_data(37)      => trans_native_phy_inst_rx_parallel_data(37),                                         --                   .rx_parallel_data
			rx_parallel_data(38)      => trans_native_phy_inst_rx_parallel_data(38),                                         --                   .rx_parallel_data
			rx_parallel_data(39)      => trans_native_phy_inst_rx_parallel_data(39),                                         --                   .rx_parallel_data
			rx_parallel_data(40)      => trans_native_phy_inst_rx_parallel_data(40),                                         --                   .rx_parallel_data
			rx_parallel_data(41)      => trans_native_phy_inst_rx_parallel_data(41),                                         --                   .rx_parallel_data
			rx_parallel_data(42)      => trans_native_phy_inst_rx_parallel_data(42),                                         --                   .rx_parallel_data
			rx_parallel_data(43)      => trans_native_phy_inst_rx_parallel_data(43),                                         --                   .rx_parallel_data
			rx_parallel_data(44)      => trans_native_phy_inst_rx_parallel_data(44),                                         --                   .rx_parallel_data
			rx_parallel_data(45)      => trans_native_phy_inst_rx_parallel_data(45),                                         --                   .rx_parallel_data
			rx_parallel_data(46)      => trans_native_phy_inst_rx_parallel_data(46),                                         --                   .rx_parallel_data
			rx_parallel_data(47)      => trans_native_phy_inst_rx_parallel_data(47),                                         --                   .rx_parallel_data
			rx_parallel_data(48)      => trans_native_phy_inst_rx_parallel_data(48),                                         --                   .rx_parallel_data
			rx_parallel_data(49)      => trans_native_phy_inst_rx_parallel_data(49),                                         --                   .rx_parallel_data
			rx_parallel_data(50)      => trans_native_phy_inst_rx_parallel_data(50),                                         --                   .rx_parallel_data
			rx_parallel_data(51)      => trans_native_phy_inst_rx_parallel_data(51),                                         --                   .rx_parallel_data
			rx_parallel_data(52)      => trans_native_phy_inst_rx_parallel_data(52),                                         --                   .rx_parallel_data
			rx_parallel_data(53)      => trans_native_phy_inst_rx_parallel_data(53),                                         --                   .rx_parallel_data
			rx_parallel_data(54)      => trans_native_phy_inst_rx_parallel_data(54),                                         --                   .rx_parallel_data
			rx_parallel_data(55)      => trans_native_phy_inst_rx_parallel_data(55),                                         --                   .rx_parallel_data
			rx_parallel_data(56)      => trans_native_phy_inst_rx_parallel_data(56),                                         --                   .rx_parallel_data
			rx_parallel_data(57)      => trans_native_phy_inst_rx_parallel_data(57),                                         --                   .rx_parallel_data
			rx_parallel_data(58)      => trans_native_phy_inst_rx_parallel_data(58),                                         --                   .rx_parallel_data
			rx_parallel_data(59)      => trans_native_phy_inst_rx_parallel_data(59),                                         --                   .rx_parallel_data
			rx_parallel_data(60)      => trans_native_phy_inst_rx_parallel_data(60),                                         --                   .rx_parallel_data
			rx_parallel_data(61)      => trans_native_phy_inst_rx_parallel_data(61),                                         --                   .rx_parallel_data
			rx_parallel_data(62)      => trans_native_phy_inst_rx_parallel_data(62),                                         --                   .rx_parallel_data
			rx_parallel_data(63)      => trans_native_phy_inst_rx_parallel_data(63),                                         --                   .rx_parallel_data
			tx_pma_clkout             => open,                                                                               --        (terminated)
			tx_pma_parallel_data      => "00000000000000000000000000000000000000000000000000000000000000000000000000000000", --        (terminated)
			ext_pll_clk               => "0",                                                                                --        (terminated)
			rx_pma_clkout             => open,                                                                               --        (terminated)
			rx_pma_parallel_data      => open,                                                                               --        (terminated)
			rx_clkslip                => "0",                                                                                --        (terminated)
			rx_clklow                 => open,                                                                               --        (terminated)
			rx_fref                   => open,                                                                               --        (terminated)
			rx_set_locktodata         => "0",                                                                                --        (terminated)
			rx_set_locktoref          => "0",                                                                                --        (terminated)
			rx_seriallpbken           => "0",                                                                                --        (terminated)
			rx_signaldetect           => open,                                                                               --        (terminated)
			rx_std_prbs_done          => open,                                                                               --        (terminated)
			rx_std_prbs_err           => open,                                                                               --        (terminated)
			tx_std_pcfifo_full        => open,                                                                               --        (terminated)
			tx_std_pcfifo_empty       => open,                                                                               --        (terminated)
			rx_std_pcfifo_full        => open,                                                                               --        (terminated)
			rx_std_pcfifo_empty       => open,                                                                               --        (terminated)
			rx_std_byteorder_ena      => "0",                                                                                --        (terminated)
			rx_std_byteorder_flag     => open,                                                                               --        (terminated)
			rx_std_rmfifo_full        => open,                                                                               --        (terminated)
			rx_std_rmfifo_empty       => open,                                                                               --        (terminated)
			rx_std_wa_patternalign    => "0",                                                                                --        (terminated)
			rx_std_wa_a1a2size        => "0",                                                                                --        (terminated)
			tx_std_bitslipboundarysel => "00000",                                                                            --        (terminated)
			rx_std_bitslipboundarysel => open,                                                                               --        (terminated)
			rx_std_bitslip            => "0",                                                                                --        (terminated)
			rx_std_runlength_err      => open,                                                                               --        (terminated)
			rx_std_bitrev_ena         => "0",                                                                                --        (terminated)
			rx_std_byterev_ena        => "0",                                                                                --        (terminated)
			tx_std_polinv             => "0",                                                                                --        (terminated)
			rx_std_polinv             => "0",                                                                                --        (terminated)
			tx_std_elecidle           => "0",                                                                                --        (terminated)
			rx_std_signaldetect       => open                                                                                --        (terminated)
		);

	rx_parallel_data <= Trans_Native_Phy_inst_rx_parallel_data(25) & Trans_Native_Phy_inst_rx_parallel_data(24) & Trans_Native_Phy_inst_rx_parallel_data(23) & Trans_Native_Phy_inst_rx_parallel_data(22) & Trans_Native_Phy_inst_rx_parallel_data(21) & Trans_Native_Phy_inst_rx_parallel_data(20) & Trans_Native_Phy_inst_rx_parallel_data(19) & Trans_Native_Phy_inst_rx_parallel_data(18) & Trans_Native_Phy_inst_rx_parallel_data(17) & Trans_Native_Phy_inst_rx_parallel_data(16) & Trans_Native_Phy_inst_rx_parallel_data(9) & Trans_Native_Phy_inst_rx_parallel_data(8) & Trans_Native_Phy_inst_rx_parallel_data(7) & Trans_Native_Phy_inst_rx_parallel_data(6) & Trans_Native_Phy_inst_rx_parallel_data(5) & Trans_Native_Phy_inst_rx_parallel_data(4) & Trans_Native_Phy_inst_rx_parallel_data(3) & Trans_Native_Phy_inst_rx_parallel_data(2) & Trans_Native_Phy_inst_rx_parallel_data(1) & Trans_Native_Phy_inst_rx_parallel_data(0);

	unused_rx_parallel_data <= Trans_Native_Phy_inst_rx_parallel_data(63) & Trans_Native_Phy_inst_rx_parallel_data(62) & Trans_Native_Phy_inst_rx_parallel_data(61) & Trans_Native_Phy_inst_rx_parallel_data(60) & Trans_Native_Phy_inst_rx_parallel_data(59) & Trans_Native_Phy_inst_rx_parallel_data(58) & Trans_Native_Phy_inst_rx_parallel_data(57) & Trans_Native_Phy_inst_rx_parallel_data(56) & Trans_Native_Phy_inst_rx_parallel_data(55) & Trans_Native_Phy_inst_rx_parallel_data(54) & Trans_Native_Phy_inst_rx_parallel_data(53) & Trans_Native_Phy_inst_rx_parallel_data(52) & Trans_Native_Phy_inst_rx_parallel_data(51) & Trans_Native_Phy_inst_rx_parallel_data(50) & Trans_Native_Phy_inst_rx_parallel_data(49) & Trans_Native_Phy_inst_rx_parallel_data(48) & Trans_Native_Phy_inst_rx_parallel_data(47) & Trans_Native_Phy_inst_rx_parallel_data(46) & Trans_Native_Phy_inst_rx_parallel_data(45) & Trans_Native_Phy_inst_rx_parallel_data(44) & Trans_Native_Phy_inst_rx_parallel_data(43) & Trans_Native_Phy_inst_rx_parallel_data(42) & Trans_Native_Phy_inst_rx_parallel_data(41) & Trans_Native_Phy_inst_rx_parallel_data(40) & Trans_Native_Phy_inst_rx_parallel_data(39) & Trans_Native_Phy_inst_rx_parallel_data(38) & Trans_Native_Phy_inst_rx_parallel_data(37) & Trans_Native_Phy_inst_rx_parallel_data(36) & Trans_Native_Phy_inst_rx_parallel_data(35) & Trans_Native_Phy_inst_rx_parallel_data(34) & Trans_Native_Phy_inst_rx_parallel_data(33) & Trans_Native_Phy_inst_rx_parallel_data(32) & Trans_Native_Phy_inst_rx_parallel_data(31) & Trans_Native_Phy_inst_rx_parallel_data(30) & Trans_Native_Phy_inst_rx_parallel_data(29) & Trans_Native_Phy_inst_rx_parallel_data(28) & Trans_Native_Phy_inst_rx_parallel_data(27) & Trans_Native_Phy_inst_rx_parallel_data(26) & Trans_Native_Phy_inst_rx_parallel_data(15) & Trans_Native_Phy_inst_rx_parallel_data(14) & Trans_Native_Phy_inst_rx_parallel_data(13) & Trans_Native_Phy_inst_rx_parallel_data(12) & Trans_Native_Phy_inst_rx_parallel_data(11) & Trans_Native_Phy_inst_rx_parallel_data(10);

end architecture rtl; -- of Trans_Native_Phy
