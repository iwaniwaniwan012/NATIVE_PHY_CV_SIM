`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
f9ticm+1cl7zuActyfaDuJnzPg+lw5aoE/MuBS3p116KpPGw2ILgy5OB+1070ODv
MF0Dt1nAgBPDW0S9R8Pq1O/dAlctrok5pFqoEiXwrn0ZDYXbsxecexicKK86LmBI
93du+LyqLg6axbK8fYBuJx9D2fUoUqf39ZJ3J9as+I4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21472)
s40NmCUu8kK6/ahy6hlXtIWLInv0qlcZ38jcEFfogGhUoWh+NlLjbBlCgTjX9EUS
1/ok4IfwPR9cpJMYZbKQZ8KPdI1vknXIMRa39C0JxIDGpAApzW/0qrN0NQYsHcYU
VTZgZmvLqzPFNfQ9oEBgbDu3WmOLjaI8Iz2w2+CYaju+VEXzJdtOz7NkeNua9X6K
uVkExkU3C5vXMuZMLkhpfSt3MaJm4uU29XQUVzlGgQXZn8p5cEDOH3ZGoozCE21Q
sRIcSP85qPnvZHW4rcpMfRaTj4GbAl90H9M23YgGcwGPaodTFAN5/G7Rh3hyFurT
hp53bREqR3c7efwbEzUF9/eWuLoh0GmWdR6LcFMjN8l1IhqNi+PjosL7ISc1Grgc
Ou9w/GmJ71MMOrPRpU2lWaLeOJFKGhgafPFDV4SAYwUX1lgx/9A18CPA3IC0aEBl
btBEWWL/SiGwA5pGOY2OuWRGrMgBJPOaFzmUnaSVJeBDShBKLgzhNNb5u9BHoacZ
OJOczF0wmvEyTPbFSkoDT9psYpailtgrliwCKKOWU5lrMG1YATJ6CbNKEChrRI8f
BwEdYtMlT2GTAssCZ2wsGSmeAsyYzh7T7FKa/9nrK6KE4ThPgfhCFIq5BOc1kuOQ
PLPwLipVzLCZfzERoHmawFqaisxilRGan9u9k2TflNGcx7U+m/yoCNMMIFklUrvh
407ACLM+mPqrS6/+6QcatanWW3nZWMRFVCJFjGe3D2Xuz6fWveQDmQdNBeOKcxS3
OqhB5eakL0lCiKWTzPAjeO8hPXfaWfBrvTsfH777vDJ8HexBmkZbQfnHHm9Oj3WQ
xns/WszvWk2FmfI7CmTLnEt9uN9YQegm53o0A2fHJ0K6WD5mz73jc5HDX9ltXbhg
08pDy7P64lc49rNd9NnWYu++P32PpiNoz5ELRh5RzDQy+jYBTJfDgIVytbUh3rb/
pLdwgkda9EhCDXPLf2PSh5iDdz+dRvvFx1ulWLdwVM6BzAAqXIL+8ZBEb8mEmKwb
6bguZ+rvO2xRYvZ76hG1oRV7aedl9q45aq4baAzYLglfo8IQAXmbhE9PaZoW0+yL
F3JNJynLdSBIgqSJSbp4DBcZC45EvBjc0X9WO+zmVO6ATnWLR24CXuo8yI5ikxmZ
9s5JGD5BAab6ECwvOpQgoX7of9z4KOxX/pN2k+VIkbpcPpAJ1ZJYJgWK8wBdWukb
WaT0Omi/qf1eIuTeWNkLCQBv1pvCAQk4e/+FBUjDRf7TSAFknUVhEHs0mIaUMXUK
0JJQKoImQPq0ERDLNGy+k157x+Z1vyRpJ5kZRM/ALSEwzBoGf/wO+9KoIcddt1k7
12tYhkWAU3JVw2Xi6WgXy2XLCEn4/woydJFdFj0I0Yc2bDR4xav1NzWyxTTnlRT0
AiyON0TcVEMYq24EiyppEosKuSkKemA8bh4siMiMsDd2eVu+EeYqU48rPXwSQ9yu
3AitO5tntilSytsD6ItAW+/AW7TH5yvJ+lqsFesRkmBA+FBgUx7z5zq5Ceb78hpt
NYXoeaRtldTWZ214cNHtKmbbNLLG45IzHPDJY/hOBdz4L3hhEK8BbIuXFV1Z2iHa
m1CsPETfO4CItaGpPzfzvbVLqwXiGiA3yxJ/0jOSK8DJa8aoF/g9yFttbyw+KA1z
ZDGyAEhi5qEdnj4Sv6Gs3Tn6FTVSzeDMWn+UcctJ3ZiUTeIXGGyg/MmwjRctDncN
nzfTgElBcbTB4v/4KvMesSEK5tzg6AjQKQTXgOixKAqrbl4Nq8knwQ45YHMvHGUE
XqpuoqKwbe1c3ZhyYyTsJbM7htcOB97iIAqVlgGtN71jr/0CyVJ9J2/ydcDu9Iav
OAOv3YCse1h2gIpR/Twa6HizL0vYyXY5601GJPoVuKC8hY5wP6vdnQL5Haq05YKg
P5pWJGcTTzAXFF9I8ru9MhoBuRhYg+CHR8i0TfhOx+3kmGbssS5xvREVbETsLvKU
oFDCjmqRm+PsCJdlnV0ZpxBZRhexPZnHG3d/T6DjrCK1AW/nc3VUisMQvA7jEOkq
gJyyUjeY8gf+J+uz0lW/mlvPWeKhKprCz/SWGsDxxlUGNy7bvH5LDdHOjboP6ELo
l5g8Xl3PlHOJ2YYeWzMjayAWhJWnluFV1OjptLTBDXz4roB7vPAqRDRTdExNAkPX
LYKDEzQgXPWFmbqSiTAvu2ECGEByFRU7aITR6B88PqXBK5RgoWI4sae5H2OViOMx
ZPUKunpUqi0Z4JcGxrkBP7biL1taHFZx/Ws4k6uIJ2RbHlTSyGMJxk2bbPjGUbsK
cTiLvTj8Q39FYowoG20UEV4ShBmbzs8vehe1GG42qVWvwMikT/Ruw7Q31huo4IaG
FYLhsyWUaRmPCMIzRXVwiypJi2MifljZABUZQlt6RVrSR9vb3fEKGmlHIVnLbI4/
CMQSodknVYcmRgVSMyi48rIYrqICpO+t7BpkZzX1gx4g/rObmaGqcXc64AFA+wp/
lwf16GJWzeDun9YBmi8GzmsSaDqPxrDOgZ6Ff5hEuz/1Qn1mDwfUmVmZfn1Yw1TL
z4VG1VyEgG+zLSeHAgxy6tRX9uwg52gidSo7HWCO6uHRJwR4dEUguxXDUwZW3A9a
bzERYuGYK9b9GV/jQ4Y31MrUjflmgetkurrqhwnSeeV0YU9QLN7CngOfwiO4Vib6
pAY7l3DfAjXnrBYENj1/7QsHZjcrD/bsn05KjErA6NOpIAMp5AXqhObtdQ36mDrO
cQgQVQex1OkYnVfgXdSi1rh/C+XH4FTm+NBM12WhA376yNnZet4Lcs+HvoTP1KLn
UTpiVHXBpM4i/yg71pAC7zNYH3zJTCXodQ+hKSaLPudt34jqQ6U6aicm2s+VjxVT
nao4OkgvHkWVltJlUgQX2GIuY0MbFqehY/XW4o+puwT6hUzp/vFkhECeds4fl2/M
qTyIwoSUHqOo84su47ecLXYUcpj4ADmlLOrxF1bZcF0Vij5GI7IbGKifOLLvP862
6aRkp0Cm2hoBhaceqCRdCfUCHt1T1lorkrjhP8d9b6VJlOR51k6j5JlFH9xIbU5d
CnoyOvIcW4q9GoMEntEyhWe0q/nFtvm5YbUoXvN2wk5q1eJXKYr9X+zexEYzNcTt
fw+eTtiwnZiYwcXSAc/ffXaXxPYxqVH0lAqbAIyhEoDNt7q8QNjnDEGBna465Zle
4J3KEUta6EhIlGScetY3/9L/sBEVoMdVm5DBPQKasqD1h90aWZLQhigX2njz3+XR
7+yPTpJvrYiDxZBAE3yKE8jgl9Jvc2i9lHxVKRhPqhrA9z0kFOprYsM5micVJO+b
OxQg2COSjQeWePrqyxWyIWFisZ2YiPSW9SDpr+gVYETcGtZcdx7TvXrU3+kl9UaJ
1mOeCGIE18FBJ5YUT+YXI9li5bDnrGWZCSWLdVNnnTzSq+31yKuDMLjC9S0jsyy/
F3Cpw/6dyYqGloSMq1EGvLSHJRWX0i9okoCLy0yClRq2qZT2hrQkAlyUOShf91Jw
GAMrvJxu3sdCRj/t0EeYD41DA54ic63T0VnS90LXkMjQux/KNuB2lJv2YYE4xvoh
IFEYcM17l2CLyMqusAWJYytKxezu+3KVolO1P3N3bgZaU22CQuQ8E25QhljJnURf
BvYubQ1k8iwqbiTCbY2nLvqsp3qPbuCSni6PHx4qKDeyD2U/TdXNIiJfHAh7mVWA
DwquM7cA4BefO8Kq4NRPmM4KEuURQkE03RuYWZo/A/VMB8g2Gh8eIW9DtLew6MEk
uPVoean1rmkjaYhK1BltO71wc2MBkKOpYPDjkXX9tqc+ayWveQYgdBAr+YdMaDI4
EZflGu/8p6IH3QWxCVKC2ZU8STN44NCF1GFI+M0bHHU2BYFxKhk08oUpNit4cGxM
qQx6y8YrpaRlOHF5pzhRIS2oXXZnqvbIAIbn5SKnUMwJrqUWnn5o9FGz8DWb5C4u
tbs47T/EvD+n8wS8IavEponEmn+4UunMKGc9EQFZWvGtOHyfsZKRjhDZPZvh8wxr
4l6UHBqXJpS1eluAUQCIIcVKBll/R9J6BDSHlpLiwBXFmpoc85kUSNsxA46NVSy0
/YpcdBmKSEIba4yq0eFeliUP/VhHUQvRNlTT1sFXUMbo9yPK6SSHr+vhh+f2AhGK
nMYLr///fCmzTB2YXx6dAl6xNimuLxYWjqWI0SWBUrwsYi1e35ON0j8/Gsc7rnGl
Llu6KkMFEeqvwZWFuCvjKG31JJ5TTw2b4Rd22J8J9hdfRQDFKE35xcgoj8IJuQQl
7KehvVq7i7r8b7gH6jd9cXgxlf7yLi5LU2fA9jRW2ftz8GcyVQpaFM1Zsnv5pVpP
nwvkDeDSrr6JmRkxlJylWXT3hNoDbSz1nFQaCfMHoVzi8qcnGoBZlT7FIYFadMPw
n/4v8bsBWVRd1cYfyjvJ1CWeHY6S/VHvQfUL2iGxn6kCUFqi3k7aWxhpvMhkEi6T
kfQvSOOOqZMxVpwYnawV/d1y1jHG9HbteFyl79hSJwX2WrZartzdePsZxBiTYXQd
T44bP30AqDqCyGCmkABmKle/C6xDPkbx9kWz/AOFWnXvGZNwRhJSMAjTAIkmbLc3
u7dC2qkb0rKa3k6MtsF7wRKXcpwGO2ft3nyMmlFNJem9QaoKYSe0bsT1Hcy9FM1N
/WLM/5RCCqdG6zblGiZuAtlvucppHz/e6HsU2kmESOQCiYEICAYHs6h9fhGuk0Uf
PMtT7/cPfziP28BnO1fi6YzJAI4cdUNLpaSUjY7NQC2UKMKCrWuy1HllwBtrmNom
kXVUibhMTGF093girKa2smzaSbtDgQU0kKt4B/efI4mZCayEzd+s96aDntS5J96I
+lAGZy2tHsAK0wedRL/E5LcyugiceAJ9DoY7hQ5JruRug7oEi1eow4J0os+08tXA
ykhPMAme5wPD+zY5i6UbDBlgZrbCOxzfHyjZpeLyorgFHIwLBzPC19EHe3TtQuSf
Sri9+fkXFstkzS4zwENlbtTW2VZ7vVB4kniVwBbr7UHT5TP5dAi5oO0enSCRmvSj
Kemy/2uYMGM3CBte5vEL5J2OWH61rpxLzDqFeyrzHumO0LRT0ZAvsXrxMQEEds+n
yMfX5u2+CjOtDMdIGjjx9OkpYNRWEWNG3jwoBbZKCIuHBjp1GufCHcYa0svnST+F
8vs9E9sk5zNjyEfwFY3vNszgPYSHy1DGP3kAGJnoVbP0D/am52I1oXw1leW1Zc5Q
nrrYxsJLDnC83iKewsZ+v+J6Hq6drRqhNS2ksAOqkqCnYivgL0JwIGZf1Q/5zxFW
QRWg7qcNZy96xU3XnId4mL/t4vfs9o9urmGSqxujhs1ezXifIsWHWiNh7iQf2Qd7
73/i5f7rtvWs5f+KpvWRYd09M/viVVpD207HLEi3cOFjh+gD9uwcHnP669iSIu5S
rzB3FJFTEgcO4YDTX+eiPQnSyOmeaVgeXIb0ZchaXVFBDYYlOGQ3kyH16Dx2d79+
2OwJiHEjUmZqZvWiuSVxL1IBUUNsYm3G0Bdlite/SX7b5hQe+FRcao3DO61UxwRt
YUJDJw7pOumC5Vp3Xgs6UQLLWgyNlHFlAgpOhMcWcj8/3mu0xb8jl6QSXUiiqNfV
M2JcbyeiRPRmZ8gXQYi63aI1FOzsdJj3wpc7pRBMZLDsT5xYC9thpLHPO+n8TZOL
EOd6HJahkLFvBBwMaORfhlINwH/D5OomHqc0PGgvYSRY4G3Mx54bEAtGsEsBlVQj
P8/0a1Uya3NFB4HJJrFSqZVUSbT39EZxfiqP8FvqSec/Iys0E7kiOsSfpa4wdRV7
2au4Jj2LqNE/cRZcA9CHYLbGFgHUX4bMUpB1IoeP/D7K/nGbCJ1+Lov0K3pztJLq
seUZdpcUclWsSFe6l7aLeFS1AlCefSxYeWoguVT0Ms2PyVa1741wiG2RIfRGjywv
4zuu7yhCZYUReIYzIcywjCBJSdRZ2gzKXnV/OnuwIC0vOYYmAJ/S4zDxXju0z5jr
/ui8b3Gn+JIx0+E2Sli0OZdLOM/O6RJ8wN+Jm3KBIU9H1nhu4wTqCeJbrRFBmx2q
8UC8NrriyQAXq9NkJeHuB2GwtmTKibcxHH9AXfL9mE1vfm6PSG+NqMTOOBq5QEjM
ce4vLUPeEvTyUom9a60m0PebfnfF+pAclhNVa37bj+2jAXb9NdJouCqVAF249Sdl
LbqxIh9LfZeixXXqqG+1urbR+N33DI7GHH+1gi5Mv3IiK1sr074Sl0svyTwB8gcg
zvYbuvk47VL2HSRdJDncamly0CfTrh0F+YB/iXH1wGaGO4CrtUdFxzh/fCf18zYo
0Yu+dFYODiWdBaCgSwzVGGxAcaKeNywkX+r8dThGkI4EUvLZFSuhK7zaIpcV6ikg
1ah90C8jrTgjuHR/c2DomuGbLHh2l7GazkmeVLjV3MJ1DT/NI5zUDhQEkBhncMXP
a7Yt0QdD9eDZACBcfMtZ/6GmNMUu/32EvVAM9c4gtO2NELYO2PAk6s6sIDfluUzw
8ZwsI9XCdZvDgWqHuCyrAsnWVIyB67hU+Q79vSuV6vaFoZ5Nzh3e5+xHIt5bqrpT
9gRa5i5Gjaky8jP9ivR2a8rjSibmJPkxqh2wvOQTQpLqPe7B/NCw90dVk+txT6Xb
n0c6460F/MchqoW2PyosyIFMdpjPaZoDGvk47kk9+/rm7UN5nX9fBr9NJ36slHzL
4a7sF62MUvs2m9QIq4pqeuKPWTXpvmG2DREadoGtj5TVq5OnI7Hvb7fhQQcjS+Go
AWD2F2qKnyr6LSkvpHAhQZhGKlNJaXrNd11ZRzxJng7ph9ri5Jl4I/VAggsvZCYy
2YqawbAU9QGQmKV9L7pznBBy6E2Pk9UHBRQ1cfPS909GIv/x5kg4vCloxGGRlRfU
hEf+hp4gGqMefVXt2ybbhcxK8yr1VH0IleK0bIrxVaUCakYQ4Ds3k7PqTXyJRylQ
amdQJWycSTqw6M/oFbILccenyXTK+b1NPcVWFO2Kpb7HU9SVTUv9VwmSoAASoaSh
kn+78PE7x2FJjZeI9W8XdoKt+1RKzRotOFj1cChEvWgqE6VvzZ26PXk1Udk9PkUx
VCQYyDI9XEzt3GYeyg8isN5qY9YgS1Aa8z1NgH4v0TqmnX0Mncy122wE0+14AIrh
zI/d/FZCDM4s4GOhQEphNxSJDD466E3aG0PrdxtMowGFnpsHwpxx7IrINUjR7OLh
U5scs0ObJTUk7U4jFz0G8jkomYUDgEQDPAAJlOJkPfEJBD7FHPvCeRimC+3GvLxV
/+B1kqiVz7OnkGSs1l+rSLGxeuTR9ALFmXeiQ3r9SompfPDcqYAO7f0xp3HeLUT6
W5DCScOi3EauIQ9900T7KKTnmaGD5SNTrSMqZiYsCVKgmgcmFaiusIU43EO3Xe2D
aJH2QIfN3qWtmsx+GCOM96HWtB9bY+oTMYhJ2gcH5PHH+Am18m7OgSQfHt/AXYae
PwgCMPFwT1659x+ZMmgcJIqHr/tmP4WY4JUzQJnidkcWvZJ412+ACWvKjEqX3gjg
vSaF9srMMaJBIWJ6Zm+527wWzKHwqAECCpDQBZOXZUDMMD0mgZhYznx0qptKy+xE
v3Eohb5x439wR5CIv4GqNaMpp/au0MFeyAtLcJNypjfWC1XVQWi9IBgx/T9vkBDz
hiW/YA7XyM1StCDTSDMCiNpKc1W3PX11aK5Lyh9mbS7iAtPLv80/+pqD+ST1eAuX
IVaXYN2KA4/MTFDTlDk8kQBzKpkp7aFf7y+naFok2RCBEYsxxSE/0cENFEz6Y8aj
bQpUZNElC5p8lyJuStSYilxfrVB2zAvdPeezYvXAda8+8XmhWZjyf8p+54zjTu04
KbOjbmq5AxsQm5SSLcx+IiZumy8aiBBjM7RwUx1qQdct2YbWMkIFVwu0EgQ3bwfT
7FM0c7HfIUwmbnhC8uqO9JemeFdBcWBfbaCqiQa0MFPT8+7S2Cfj6+nx3l8q7Zt2
jrKTJzd+B34JPwbGLD7KJb40vCu4QAB5lZxVrBRBgWMcmWowhBosg/iz6+DFvpuD
4bJtQX8rG15bJPvdNNnw4QNt9zNFPp7ZZ6qS+Eb/2DD2fb5tuRY3DcSaZFJapEre
/6ByuPu0YaMHOIr8O2odtLQCu8kwWpTE66RBT2J240fv8ui0qzdmQ6k4O+OUqCiu
FwGfyuar6NdBrDB9H8r1cmf98rn6w40sbgig/uSBdO3eyCyj0iv0UrV64y1gXCGV
MHe/5biynOyVNysGN6hywy8V6CTLwH//PlZXM9fMp/YCMDcDzL4XZded63e12sl1
nWFpYx2uaBTUmZeLe6mvVS8pS7bzlQZlfgEnD35LnsIj87ozIbpjnAgUfdRhjWKB
J0xg5ha1c/j4x5DX2pOJ79SD+X2wqnittKdH9nf0SnQL0Au8VNTJQ+/i/BPRJNOJ
18YrtZ2O8A4IO0WSgKOprrjSxa8URVFjkUGLkUcrUyFSbqSbr/BlLdH4ERIRGv0q
gWBJhtWIqij/11wSl036GzeSldAPvC0/Yp00c/w1UyzRhTJRx4na+8tXrNHWpZWD
18/E08yh8F1ETwcktadPGRVS7g8in5swu0JC9yqydcdDt4Mj1sV90SfzoXHwWJYQ
8Tat8NFS3fr4SWq7xuFGK8pX/0x55S54rLvdsImkb1jV+dtKWNl00I7q7l7Cvyxx
sSwXrnhPNRANDVbUNqGPOyoyPKO4blI9jKJS77x7w2KGF0PFLkcknvlyDNFBpd2j
pQ/iyYu2Xnc79JcNJ13mr8psAbVBzWQaXyAGASmySS3waTfn9xiHGh7Gy7BnaNp2
pujVFv4jWboI222nEO/VuzaceHK0auDTVqQjBSemAFGIBT/4t7sqE12UNIsRdgQx
nW60ZeQcPi8IvEAaRSZmEMd/k/bBOUWpi72KlCtVf/AWTVqbUTH0cJ//xzV2Xd6R
qQpKFLXdypDgLFq2GEcTY+3Io7l8woE1tNWJF41IE5Ixo/91WuUtIoIgeyoZ7Uzi
Kyy5MZJ5LqoT8704ppH4bZP+2/x1RLPgPRUJwJeIJWeCKQoWChIGNpDk52WUTPSe
m/OvSCeuE+k/SbzKhNP4YsYA+zDhACPFzo6a9BAU7aQTVUObeAxtpGfq3jDbKj15
N2ZKsjGb58Zupmba+JDDCMp49/IyVrxrvxEIBJg+lmHtsrznR2AxiOAtzF4iIdw8
jf2eGnKsFRwub9U6f+X00cgOLvFUxcDj8TaCAayXrF7Xlq/zn6A/CRuqll/qAGo7
ylxbgh6SzlpQ1WCxo4LSSUG184W542+cmyO1u0V2iOCp9WPq6FeV92VryDTnSXAp
OKXSJxs4loClzmY0xK63WBi4sCYJnMzB8CLeZyNh1ddQ0ithgSBQUn2g2nHw2/KV
bfgqmbPso4MwkcU6A3uEOPMdChEjSFw5YzSFGFv9hcoJIU3MR5aV2oc3nm/fcR9K
DntVVe9tnC+5p9E2hq+q5wW2LFcWiOD9LjYUXTWkE4sDiONiB3B/Sv0GmFlQsDAQ
9ZIFFeeQ6EZmefl5pPr5liksvbfGQbGINP1Kmv/LeCvv4SR9wPRQXa2uS5AKTPb4
sFrs4rdvawx6u6pZnaesKZzylesXyk0v+v3ndh9BXTnT2vJDpls1nFM1JKkIV5F4
AT/+p+sOgqBqL0v3A5oi5ZDsWI/CmyExYojg0n1MHnTPeOWALm2/WNU0FXrmpr7e
3lPdDS/+8sAM8q9qcL8hZQQeGMDkOkFbJaZQu9frqB6dZ5nkPeXnyeoHE7JmIbrU
QnwjoISDmZfNSfHUfyW/nRYQOdm+z6hCv3+5BuewFTUoK4zfjGL24IWtpi2EGM3E
Dx48PSpPmEylcWT465EZXbBoFLO4oQSQFMNDQDvWx2j+E/dF0+dtJFfov6uFLM5f
DudtBQPxUU+YJsTxv4c8TbYzv+UuGcahMr3BLJ7L6i//a9f62XNY5UqWPRo7AWVh
9Jrqc34+/oseGISg8kvZJpgyT9MOLuXqX0XNWOe8f+FxKM0obRGSgSZNBdnWyiLT
MVo+54IC5mKpeWVMPaDN/dCWM78NgHkiOzUqySrljxkDD8BEIMfZ0QKThPFbkuFQ
dDAvJ1j+btzbGuPBECeDhA7Zk55tnV9Cj54hvkkLwCvrscyCTQErMlKlqxiPeIpK
TafYouuRZFRXYIqxR2X2BNbThKHihYWj+z9ahY6YvuWYkFQqKGFkZggp+ByrWA7F
+XYAQr6tgMuZmW0BaX/mPH/SIGU9X6Utlg1sQzDIbfHj4iYIN2K/xdmhTN+zV/4b
wkR4zpsRDqKrrlBfCpuwLQvRR213yc8Z74FO+3ErcG5t/LM3zNid6w9vopGb2Ogz
8desmYfKGXC+p24i8OCVdRhGdyigP4rMvZETtevJwnz4xuWYFhAnrXeubS9XoLzs
Qy9Lr4V2gKFPXRtzH3T8eUfKb5bFuJxhNnCcWyhFPLuW2GgqFie2uwboty9Nf6Cz
jUur/ej5F6WAnO4owAiuZB96NprK+fH/F9IsY/0KgDMg7+fWPz+eI6PutDQ28vwR
3/NJYFIWbw+KIDArtlImnv5O6M/oDslD++7qRAhoRgHOs+3+k6kYxzmI63tLplTB
hb5HjJ6EKZAFPh1lF1VxiuNgep1Sn8Q9JUa/ugabOeL5oOglwq/wKTfBcRiuCNt+
zsHLvjDziPX6mK89FdNeaxU2uaxwCpJqzP7ioe9wSd7Sdma8QkF8FODKofFNdxgg
sfG8hnzPW9Js0LeohEl4cyr9el5pfLP40kjQR+d6DPIXoXu75QdI8rghyqOiUrTE
bslfCuHUUoBrSZ/s7dbfN0BSoGfYCAMgIZSEScANKDF1yJBeL7LoyGlBJSgicYfn
rnOHRpJEUp524wJgNWj5YcjCs+5/Ms+TIxY7JgCs2GqlubSF9tuzowQbOa8hK62w
cWtrD1ec9AbDcDodSlssJO0MoqHwEjJ5vimDqb34qrsyMQqkZs1KxaeYLZUIIWJp
hyfteNlhCAWhXche729khY4Hx5gq5z14M+dANFupcwXLI4GHCL40jUOjVsqv6+SJ
1TFN92rja9ci7MTxEKJQokJUdI7J4f0DHgzPaY94CiX2Ug2iV5Cvlfg5PP2FQsfm
mmUYFiu9N9j7rM1KrDeHPgMpYES1L2mSnFBt7m2DssGVypCl8feb1/oSpIwrSnX/
pZcAULXvasoPS2KR/r3DS9Ivz5fS6KHUmgfXYKe91LO0bU455r3npcWRzNurXpBm
+PPm2GfEkw+Wghh0UIZIHLX+QlzPD8jpeTwMlVOHtPSC0F+yth6GjY94Sb2V8lhC
225k6SP6ZIzfYAzVg+3vmNbN6lGUqUuiZvDLNMWni7oqeIjZ1VfTkx+H4YnEXs/0
vcd9HJkSrk6BDZNSLicWT1DJh8fvARQtXueIznSiDoZI1VVptHPyTIk5LTnGcGV/
9027Q4BUgStLXMSWRPvRiihR2y8iC+vO6A/hJNyIye93hBbEWdnnDA2uAKCKbyl8
371FLohnywcp1g/Q1l3wfm2TKxyx4AFU6pK13Qvv4NibEjB3jpzVG0LZ5hiJUZYJ
GX4Vw9I6sJP9qvuIPeRHZDc78DpeUZc0lgMuEZwglbUNLiKIO6AGu00o4O0SsSy3
4ptiwIuxM2W8ns5kwYKmbp2KiahNHYNEx2q/JL8o0YDemYh3gfbfppPKCkIYAiD3
IiYmRTnCakD7g8TrEolEC87PvCFBCO7pL4RAhFCl1gbpe2bJNcOFUunDqN5u0hPP
Znl1Xjumj+aiJEEYLJofXlJSfEs8XYuS9nIUsXbknbBSeuYyO4i63rGjq+7GA7Tr
1rk6H5h/tdcMigkW7j/2sQ550HSkPmpxXkuIL7/cjERQ7OoUebX8dqnFmyszOtpm
mPhObBvNOAhwCTVPBcaajvQsiq8F3pRpc8sQLOZuxn5atSW8BPPxcwmZ7/MyH6w0
bZ3pBMCVY1s3ZTJD4mVkDt/lM6q2M+qfhltOMIPAdeyy1rhoco16Q0KckKXqgWEe
QPLO8EjlOlX/+fykQFz9ImYZg7zPxhjHzZ5fvDKRUATqO/Y7XGhH3OoNzHyvz45C
v30hOdjfRg3+YydXR8lI1D6j1ElkKNqKUm+YulYoFd/luwNwBJEXYZ4Wq/o6kJ5d
iI2C7QoRLoOI3rvTs7eEQ74yMNeOiMEKTQ5H754mhvNGKIwBiBchWEEunTrY3Osd
I8aJn43irZ5cq4W42MF8C+DkPQ2gl+irwdPLZm/KfoSVz6ZkLf2WgC87s2wHF+8q
2DlLT/GAjP3pC0IxlNU+4cSKjE29tFEL6HKgmA9Al6gTm3s7zkTHOqIcP5PHR8SJ
CAMZSjW5mqCxdCFugoWZyNijCgvSlxepm+JzFwuEXQBmiQAUHJPH4eY4eSdXtOyI
HbFSY1PfniLIyeSW7298ErGY7OVdTLKSoNDy3NnuaUeRtjhKjyTM1fkVKJa+Mi2a
4kwBlMJZXkYMYXG8Dk4C4Kdc/f2FkFCwNcf4QRoiXWSBkomTCRVtAzm+ZAGMMpGx
JpP+5Z/t3btXSTxOcOqTCPLOad94NblszzLoa+2SD0OLAMAqJnI9IP7qR6eyF2B+
5wPYrRaDliJskQdo9UF+qegW937RwdMCJguK8MKWI9AY4bdjBpaAWg52CTqV+l7d
QQBQCy97UeY/mi6Fs4AEtp90TEi4Q2qwCfM/YlEBHx/lSNiMxZF2bwcYip69XPeS
7WFUW6nDOhsODLWBeGPO8eVWbU/ZP4gE8bmZ2I47Z/FFBRwJf3wNpDyzILWokDVW
V2kiCKLMvIh9wVDHju6UwdV0gYe1fQ1kSSC0Y+dgGYhBxkBc3dyuE7faQbgnG1EQ
cY7bJ95ykYklMBtVGzmu5/rTykVes1Ax9Uoc+QvZGwcFAt2ymkYL1A1XBXtkA66k
9/cBcVIYTdY9fpHM+iDWNJ6GN3L22j5Ak2LrHDT1K4tsce6671VRWvP6C7QKCYGO
L6iOTfMCTjPebru7bARQMcP8wut9RsD1otRzt4X9yxX4e+PCRlnv7RATjz+ZNWl5
DaWqfu6WbziLPmgz3dkhkeBEc5lAAIAuNCi8lWi+8JiS6os65I5rzPKBif1IssoL
xTD20LkVst6546VDFwHV/wS8Bvmz+OdaG5BOk6O5TH8y/gjK5I5LWJ4kz7qz6xHr
e6+KmqvVsNkwYqmAf1uzPaNzo/mSV9PqnL0iCokvkL9HuSVfsnCCYIDUfOCMTv57
FmpAt8EBb2gfHGUzMUFtPWBpnGsPW1ExLYx6NUuzPG37WcAktwjwCZMYYK2lZzWV
OcxPrsX4Oz23R1E1j4+SQvtwFb6ngap14fOJqhZ9pv3kDtWrB1IUKGY4wiaV/N/E
vWKSz3Nr0Vjkfs4pkY8wmvGN53KrIEX51b2CmBpg5r+Fjwd8hbUG372/B1tSl/KQ
/lA3V2f8ailiciqBmdTFlZW2cTSohoXxFPBJRKFZDjXj/foOZ3jxJ4sXZ5qwfnSF
rjXspVL+CRi4PWK89To2aa4fqQy0JToO5xOOmwoEp3PKf5OAaw8oAispXVc+DKwA
cAUdI05UEQ3m+AefR6rTU0wl+sxH3YIEuqAHX6K5gDcw+rbvKgjh3UhcfnGf8io5
5Ajdgi+gJ6lGQYIC/lOOfEW4y4hE1T2jNeXcDWyTt8PgMsEPpdRMFzWzQRsyxINY
FFASRdJPSb/qeoiC1vucRu903ZtehOzsQQPW2kY1OSEOG2CJq3ZkNf0ZlOiZRgfg
+NGffZpXKvxQUA5oC21pveHc4juKTGYJF6ZtnG9sCNALF8VadBTm1afCLaYnW8q7
ijlpRJLSXddFroFcnFt4yneI3oxO1ZhMOIxv/3zfsGDGfZNJiolJMotdLDt9X0pb
1A6VSyDZ483kBO1o9iS633p9UHvDlCJHgAbSzgBTKR/MGW/hcLIPASFxjBb/irH4
gPGxf1nSM4MMF6hXHMTNP4PgC/z2ejFsrvkOb+GRZNtsu+6AErLZWMNjXH8gcTny
/86sCC+cZ7xMGS8pW4oBSP36NXwmKpcZ2NyMBlfp2Fz4+sJxBt2iVkSWZnhdhnai
MAuReaulwed9wClwrWi4DeQWCvXtdzDBSSHtTXZ3puEvSf/9UrU9eAIJi5FBz5Xd
LnTjLHcGE2TbYz+ZHCxFCnleu7++KMaZSWo5l2lE/rlVaPuE6AJzuREX8nrhkwBt
9ykRF4ewGg753NtMGLIiahr5q8XIClguOuv+gNL8WNCT6ShywotobLb7lXZ8Nvnz
AZobnwOdl42L0pqtrGLnbemq+2dOSJj6deQ4PYmQQUXNYtxOF7Dmi0ffLvyBod0R
h1Jf5ekEbognVEp2hNett/4JOP0gayNhn3DFu8UWw0e4IJfTIHfTVru+9oKVbaT5
4+T2l64asJC7aomzB+M+beviwUBH/M0aYjz9MdefvM33PSDVt0aRioD0kPgUeyKK
vELdeN70kfcsckDO6zLSSjL/JJ6LFDt6FBvX2A9CM8WrJ2Fv2eZln3BW1BtYGNF2
gATefyYaFpaEzts87kvUKcbairHEaLESX6XSF0/gAKUr11xAwW0hEAhnrOsyKoxt
zNlW/CmPnNN6Sby1z3v1LqzylvgnooR0uuY+5E5AOHiOxjP6bkJHUK/QcV2YpxIf
Nm5+IxwrwEi7vFU6dEGyzd/KqCQI69LpHH1bZtMUqxA+OU4b7jGqsGZztJiw0pjm
/NtWbTSp4TB2ErKufqXYbmqQ9sNR4pT2nPYOT0LRaJ0XnUdd6h7MWmLU8B435Vu0
NOMKKCcZ5h3R1R+hYuCHDCUhjpYOAnoCDSIraEmbgVYl360eBOnsl+7QX26kJUkd
sYKi2X4r13HzVsRnYE2sbMFIIq3isAS6GM3Yjd9ibAByskUyGGT0KyMZ4Tk+QAAu
VnqBj9numHp7dJtSVDrN45ktb/bb8fYK3J5IGgve3hNT0hzAswpId6UtjWzgyoQ/
x+orgMdFVssUySCX9Hb+lf+j3InA46pvVydmRyMYtkFIwwyCIjzfIyTCuDFdvEsr
PhvNkJeSu1yMMHulnHiA/OWrIkkaUsxrROfiYARisYNFsrDtB/kAA80B8FWbQh37
Or1Jpm61L2gCeAAUq0pi7VTAR7U+znkldJjyBRV0UQ5xGfDMQ4jybFlDHXW4qDOD
Vtffe9B85z3NY7/8ZFtsTIESChtJWVA2EV6o0ulSfeYO0C5pM5KBCI+Uz40qvSNS
e6BRAB/eMy7TA8wBpspwjDnJ2C7I42Wcn1cS4TynL+DM1d2Fxy6/229pH5ihJI6X
uo4ZWt0Q8JjOAtyMuO7xF7mORxcopgg3GUDwMB2Ca+24o7X2N/fO9tKFx6DPs9Mi
9VrKBe1SgWceVjqm18biKyXZifhwqbaqB/NFK5M/2iS2TqII/vPDfm0rzzQzdJ3x
GcUCbptfLyzhlowA/dpJkE4YAekZ7o9wLlEs3HQdCEFntp/Zj0gXSQH+0M1+zODV
enmr8Zbp0LCwakc0LPF6cP9tMdBgdssNzxloXGuKJoT7WLEBDrcQwyIAiqmtzdsK
xdZz8FgTHkv7JFuDfj12cpd0Pj+/uUQJxqvVHxfIWQ58SpNNNJhiIx6qft4vmeaC
FCOihcbksN1bdRyTFHlhCCfHcCqbovUnTsO5C9TPi6fJFU7fhhho24j+jKywbVIW
FKSp6TOGEyfywisdzFk67KI3k2aCiZ5OU7JH4rUgjHUaT7nE7Dtnx9E15ohzf1Gy
4F6GVbVdf7bc4V6Wey0X7bin6kPEo7qsMkQwIZvgvsohFC+PPOBgjFJo/EIfHHCk
qYKJe/cBolsN79kkdNOKRhVGjspb5C4NDugdJPEyxRVoFF+zNFOHHIzBeg6O1ytw
Xvnaw0q6JlnhahO9WtXEPjvAyQb8il9wJXPEMje70Pk8S0LGJLhYB5bhbl+jlzzy
eMGgpWrsmNekXSEhiREF9PSXC2EGgenjSkyGEECTWJClSXt1+Q1vzz7b2SO3UKh1
ipugdCBnmqzlg4yoZe1NTSk1OUE7kf1zRxreV7l1XU1OeLDKvX6hqaxR0n/ft0hy
Hi8bgs6M1kFMMG6GI/A6vkWLVc++3g1ET4YeqYXhs7nInIABZs28L3ZrRNTPMg6t
O5joUq6OMsOagljfDFsgJjFw/pSTSOEcKTBY/vVxwRToBSZ3l2odEqFngjXGz1f4
ZxbmBNpCFvqzX1ZW+CSztuqgDT4uO1DGtWk0sazwFj6d8CZ4n/g4ZRLMll1scj+I
1QSv+scnGieVVLZArywmuk9NEtmJDXFbWjaQjWCbit9PvVqF1WfaMIcGNKmdof3k
bXNwVB8MiH4awfnbCPh9soOvENGyxZTuRyyZMGmAtYsRIOSJ50Fq05M+X35FNveC
wU9kCpxPkaMYUQO67iSc4/pkuAoI+0w50OSxcU5EQ39XTtdUHaakwRsHHu4WH8PY
DTAb8snbmXsY1C1JGi4m/uCj/crmVTNBFpE48xPvDuRxoV4ZV2FK96UdbEjyob3I
Hp3nX+fMZfF5iBEIyZ9WB7YXnPbQaBgvwYNdphWDtQe8ezhwnbOAhuFOHdqV/ilu
6Q4UQpJklVQvwoGuMYKLbZ/FV0aFHpPI99IHFdIcp7Pg1sYhEIskoX2PSS3u56+z
2kLkXSE2hitvMI+bmRAk0kn3S8pRg46QrUc7s+zVHzWKJaO2Xz0dH2V1GRZ2PCE4
/1UyuE5M5zwO6hNGUjz8gcsETsx/YzBOgm7/p05UYG/Apt8WmJVfn1ueK8kFs3WE
zHKPwxFCIW7hzO1tngZ/w3fLBF2/WNcmoRj2Oxw8/i6g3etERfB6ch7cBme211sI
/1a8ndbVgrPCuM3EPDkNYbxAT4Q9FRLoAuNAZY6Yy9GnsSDOIEAwjynFAsMxKkh9
PoPBr1Xp/S4Ae0nMCqcjJxerYIxNaIy9QkUQ6kjKgxgyKEJCNYRcqwWk+u2PKcac
w18NzEnxjArfH3EKBJ2ho/GIa7NpoASV6fhDexSBQ0BCsbC2dzbLA4VNVOmbURdi
y673oIgNk4f6FjyEs7/OLkj3wpvh0RtU+Hwcmqu1yOgM/822VxmEsea4kXSLzB7E
icx6PgASo8UO9RbMvMUU9xJkVmSpISRV3ifApcOM4tueIpOooS1APhU907B0lE8x
W6UHXXWh3pFJhawUQZzTjyasZv2BescRoKieVVYz53lyGHFakbHA/eJyLS8l8Hz8
2bN4gBY9EuFiVfTnp8gncjy3hAHxtZBCVLwKmyRYZ5+h88JDdvFgxtGZ0eqd2nN4
3crUYRXSwCdwxGmtZ2xXAzkuaPjhn1Z4A1Ct2j8OYACcsiRdHy99o0q+QtYu0ywj
3RGVR22mRdw0l/4hzvN4eJM/3hi5rJJORuQBE31t05+qei2LtBAAonhBLDX13h3u
eWzeNClfPllwIEnZfStkCbVPPD+aBsbp+ZmdzlapGjm6589HhW0wk1jqydpKq5LL
cmib7WCfHi3YUrJqeeE2JT3jPAqXkkbGe5w7YAIwWVyWaqZHnEpmYXzNRGk4a2SC
s3FMd60wxcUhvrOMGTV39lezyniw8Imep+/QWEl3GggzGEPu7oZiW4c9b6WT8/d+
xEr/Insyu4eX83LuYv3+RH8/xb5EeTkJ5LOngZ3e+/hQ9IZWBzbGGVqRqjRua01D
J9WBo7vmf7bOH/901r4SVae5tUSkaZCZquYfKn9g/jIEO83FHP4O81QbDz2CTb8X
xJxKa+U743HB4Rdrg3dWqgsyslbfW9nEPDcbxFu3E051ruecdKA82v6DqtZJqMs7
mVzLlOShKwDaFLZdv6BvRvwaijrvbGCX8PH7h8yjzHRFOLgm+yDMZpe/w3+ccgoy
mfsoG3nAQjl5k8yWQ5mbjYpDsSMC4h3dNMMm8dzcygD4098QJrjeFv3ZzBubYPHj
JEMMxF/fHsi2g0/L4XbrSzCJ/t9S04DzPMs6qYlGoCJ+H9I6CJdDcCanm+qasHb1
vfI2teDbOj/LmFfofMa7rKS7aB0Vn0oDLSquwSPHTSxLUIyoWhj2+/S/SU4Ytz/t
5HMubP77DqRB6sMqCI/AaLVn8K7T+0jinNoWfqcHhclvvgH+OLKWVUKHXrIEheZ4
cBTUMZHfFgkRXxGlQvO4+VYqKfN3VVdlbj4PW9kFNkP6d1KAXSS9HLRnYenUY372
VVFkbpAtLJwZhb4H04ugH2QEudGVSajzMUpOoi/7ax+/ekcpaLUyJajXO9E1Qiqk
rCEbek/tubjDKX+z6rug7LF3Y38OILJEV8gRaFXYX0zJ+M/grksKsk4z3sYsgE5I
3j1KZR3PVTQ3UjfDjnDq9s3AHYZkEWXpevD+X+IWvCgIvifR6cYTNrC+9vi6w/Ju
oDOC6RpKl5VC549gbqD3wxKyX/NLsQpFzDYMV/T0fXx1Hhbx0Bd+m9emIkswiOSb
EP7z0nQIrVtzx5Gi5kAqU9qHa3SpDEMwqmtYY8ycz7JY1JZc4ccaI++IszxBcNMb
AdQgxcsvdBrRJeqHPV4D1EnCUSSjIFemz+STVQHoLkyglqlFsD4UZJfxYtXi6S9V
0+6YZn9y/n5tu+lgJ9YVCBbMbIQ9k8ZER4ICUy3bD4ZIjXCPRAiSruHm96jqNL0T
dJsNler5fVEqqO1B4YeMbGFgtrP4s0BLzSZAR74ZfNxz07bZ/vde35vV7a6pQSkr
CWbn+xxmkPHj/T3zTL1JvD5Nw9nBSjZ+PEe+2+X/TNptKen7sazNvMjFjmX8lE3+
nxPADzLOa9A4C3gnCKS5xY0G8Y9VHLk7Uh0ByB8J1kzUXC0y3lYKBUD6vTVZ0nnI
xpbgTHkdmBGigf1VaZ+OpbRi+0nzSzB/HQ71rIbAgnMd6IshEfmHbPBaeTd96A7m
7M23raO0FaP4CFJsgeU1o0Dr9ybJvmcPwKig8Jqci17KP/jnNtmpmIzEn5S7gyxx
oQMUiFHmCFsJDIKB7NZ5LqnUv97b3nqgl21Ubkgw4A0WacHhgEZ8FBJC1goZwW9C
zfuVg3Ex3CH4Zi1yLGJDbWVfCCAHC6AKILXECPXMssuw9sJekhQlRL47LXqzdYT5
sXOYk7McCSQ0q4elX2v6daBjI9WmKKjHE9mr5Ia9puyPjURiTWua+PR/EaNZ8v/L
XrygANIFS9Ttat2XoR2BrsI/Ykh05dhbuSJBKQev2lw1YO8HQG/rlS+XvIK/Eaa6
dSUN3gkXM7o43dOym9ZSRNj2DiXy6tJMQkAw5yp3BtpF6HlL8xGL35q8SxgG52cw
TU3w4fOI9dzXHCWlIgjhses20oGzEZpXZ0TXLKtimKVG1ZSxHqirVpIPUjPquy5h
zBteNNQlVOiQvVbEJeCkrYk/n5KdW81sa9iDPBpugcZ7I2tRS8+cY6KyH9nDSIZm
Wt00ffaaLu8DHibXQo98yTHow8qsQ3VIRSNfpW1BAvxYWMSaSZXsunYK4O0uwVBA
138NJ0bxe5MHFSeIz9iMWpF73o0jF4hbDEIJbu5CRJlMPq/jF9N0jgYjtNaLUjXk
fhBOFf6A7q/H8jTMw/OLiZEHr0gj4j8c8nrNfy2d89rCybIqHh0ywwyUzd3smB/1
PHGWu25L6VnVWFJQePLxf4KHwA3gTZnyhDoXDjLBqUSfwJr2NJwOlFMt9KCYP3V2
OHC2DqhosH4Zt+xO3rItje4F8wvAFW8MlPuwCB99Bv5rntgPXpV4+GmVx8yHDJbF
jb7q+l5SQJ0gCcBjnU38zI8QBMvCeTM24EzvN9gVbqfmJC6AZBbj76gkoHi/3Tz2
tFaZNYBHweT/Ui9aI4AxO/BD8ZbFbMkK8uTJGJ5JI0zY6TahpXCU78ISEj50UcwW
Qz4tSjOrObdjoag/zmHWUHgAZkGOcEM7RBJjODavnkGOI47hooBpiDEecsKw4B2s
Uiawg2NhSx3PvtxFnrevs20JjSx8ESzwSbsc2cf/ks/9IcAVEEgZSo9/38Tbnytt
D0bdnZcRua3hhI91T0QgkA//1aS5MnTmnLPE+pkoD5PV1LwP9vbrEp4B+kM/jbY8
/3x/fbAnbnx1n5x3ZCE+PSjFq4Frq4jCh+JgDluv33HLdUQl4BLd5YfdJH4RMzji
yQBpIIS7aPLhPMazVLrV9V6mGOASpRQIHfZgtLlY+4EndXbZVRHlym6onGXGmnIl
rIOGd78bm4qeT9Zx25442Tn7u5n4qNryQkK77mFohsbYQRBO+eabijonXgcTVHqF
TC9hpY2I4N1wA9c9Lt8/vM/MbYI16+wAdZj+9ig0FndFYydN+ngraPgrlQKUbRgL
QqBorW7UZWcGSRImv8Jprt2LxWFlMSW0JV9hhq7l/PyZqQRUZbHnuM/B94AxXMZ/
QIkntK0d6wDqJyGvz8flwX3G4hBV/ds+0fCHIi8CBS3ZvabrQ6V38VIHeVPzN3hR
uFn+1vmYzmo/zh8qITa64P/HDj3Au0dZiV6BzF+xG+qL4GI7meRDq7SPamiPFZjX
z8WXmmNKnsUaMJGrC7cv6kagCtHMbECF+RFj+pxdZ+f/qGnAzk7YlMgTayNY4ZRv
GfZI7IXD0iKAf3LuEjbveyHq0MqurT9SYL8I0lNiLTYHDb2hczI2fj9puwTBE6pw
YR4GIAfWam2lJWVtUW3MnuIzdoqJ1DJs+LKC76HultRRWjsL2DK1tuY+FMuytC3o
E+bCxz02f60Et1h1+o/USG4Ob74Toqg3mYcXEeLz2n4iuLmHGocnIO+0YCaH/z9m
EF274yB9jH7Gge2IGlPXa3NEcePMpCyPPpTPkhnJQnWNLMvRi10a4ACGc7GnWZl4
fMZvDf+m3dZCnZ3B1zWRsvC4bf3HuFqJAomM1/kl16AxSTMq1lfFXeHtN10QjDKE
PRjQNr0vKQsZKYAc5vtb3sqKhNYvGcCRo477IatEIE0i70mpqmX57cxXwZCwjwlu
8qDMxsdEdju/J3W4Vq8Be4CGm5bdHo6zxIkO5Y/sKJJsFFJ8ytlZaZsyGQj4FuIA
r6HM0coiaF++uvLdO1QMHUKhP8iS3vBfmlxv+kYBZjetTiSAevJCgUQLXnWmtrCf
IX4mDEnXp4c2kKX0fVzITpfPEqwsjCmwRifmhsWvDdp79UJRXbwjwaLbTxL3c1Bm
S58GV4NoEK0mSPsh9qP3aqUDEtjHXGlL3dT+lcpiUJW6ROiK43RLg87PQeKOvft1
rShhw0rNYP77/EbYUoyUGk0ZeMKKIPuOyLDcrZm4eLA76DjUrgOBUmUaZaEQJSKU
+tJk5SMbqEYYNzochrMz2tlCvM8A7Sig2gEG3wth0n7S0M++11c9tclC0aBzDZKL
CECtZhOv+VLliZNtkHBeVCoGTg7IdapWW9v6hTx8+g5kNMxxVqgDsyYoQ+9L27l9
I7hzvNehSOvkYizVF0+wXdb4X6oRf2IHIN7gxZRuIzE5/gY5G1Nkd7qK7ZVEzLo0
jKawlUx4vK7/taU+BN6woZl2HxfBG2QyHjN+7OOvO3OWg1hEhRUMOcOy/b+wZNYy
XpK06t7Au4M32ttR5PFH3lts9Vhl7zFYKLNgK6yk9z+xI8/foeTAxjhgUw8mAv8X
uHAEYg2H7pmRxvhKsCP8gy6AcIHS8sshuRtbcOgLmQ03Hnz0gJt/ii5qAxu1ELoB
s5pWvTKGk8vkRkA3k0uoticJAVr0fL5Wx14gSXTOqwVnxpsXMAYVYVoIShTT7vYl
0y/XkJ2OL0IFavFtc0CmV+f0HqD8LP+wgmTkrwCHQfgw9q0jC+hZIs+eKxC/RPnS
9JAa0R/wVquSG6P90R4nLbi/M14VjtF7EcOkkfwTuYodF8A19nHTtIGMqs+DrJwq
slqJS52EimgsDjaM08CWH/COHVq/F6ennlkktrT3xAAIJD4DuTUyOsV/fPazr3ux
q8HRhSps9U3pSM2o1fXlGFWfl00e70UUHwr4Ul7Kyg4buqTZ30DtWR5oMOlq11I3
S/kC2vlQKChU/yl8SrCRQKFnm9NRxbl2AmgwKMFnzbdzGIZMYba/Hg6doFfW/iOC
XUzhOSfH8XbOcRFNs9xWy0DW4nN+YdY44JtAYqKODP//zhJvMPL6xW4CF/Ks9BYa
918MGYF/4AmIcAAXi9qtF4bX2kTyjHJkIGNHGN4L7Y+sbTqvuknwAM8mHK9vm5rw
d3t+ss5Y2MC61ORtuBL52x/JJjp+qb3kx6L3ImWtpUhF7BF0VF41BmcFUEhK9g08
p7EmMggxst3MpqKqd6n+RhdpNahjdTli+m3YErWf08UxHKc5smXF0w6/g9qIAp4F
LcpwtRw1tnGZdyVm0TZzd/v/IYFRDzCrgzRilMJ9Dgu0ckEd/CdiiZZgUKdZx9/I
DupklnmCHchM44ZdTGT0ACDfJi4d940VgL1xyJiDH1R4MrFCRfkESDBT/zlTs3DY
3zVpzLz6/mtpLVkbUtGENvKmkg/13JpR/2vtg/WecF9SSwZc30hsVyC3nUH31Wpl
Huvm1D0jUjUrY2xmLPb70jzB+6lLth2/IbMVGhtKRu0VWDYAty/DLpSq1JX8IwKq
+vN1T+Z+PYtuGICkpOMxoh7yJZ8sim5gIMMO6l6r4lZE3e6klhs6+Vomdc1sfrq5
c/iQTXYNxG7jkS7LnvBrM+R4tMtOZmibjCMb6idk0nuohk/cZl8zHtPbfaV0qEl3
LTj1UK9g9UvSVRzn4gALJOjFJZrMafWbFi8a8Z/I4Q0G27+oYtK3P7R2UuUoX3L/
X9LiVaW/zA8WBne+OFICiG5/Kz0Dln07NY0iiX2ZDBU9MNgieotoRPDdxCKEsdBz
I0BgBgL1Qbag7mvJ23Obfq9BTs34RZeIBPWoqVI2iJ57cKY8KM2Rc7h08uZ4E2sd
bWoNlt/OSKoTpi7sj4DYtmqXpCc/wFkV+BA8uzQeGSqCqw/AFiheMTLEdX1+1sI9
75GdnKcW8dFvhZPId7VrtjZ3BHYjXAn35Ho71IIJX/JELx600+ZuNefisEObq+x/
G9xc4eu3x+jMln1oy1DTUMBonnPauKTkc8rh2EYutjqZNb+4jYzQvtNhTG9u6jzU
m6Fd6dSge5XE/ffQ17vjNhBRnesTtgEFWoZvFvHC5SewoUtJHnnuccwP5AIx7EwU
C8tqkLwbxa5W91TqtBJsBdloElozCYK+315AjvXQsiL8zasAXD13UMQBfjfYct9Y
ofmeKMGd8nGiO3xwS0so1hfnAbqGP9zn4zluJWwt1+f0fwR3om4EsSTFS9TTpZI7
V+qk1ttKTkmrdeEQCBQawejiL5V+GDjeRGz5TKr3KTJMLblxXnmDieL1Bzrjjcqr
urIe3UZT1FNLdKYPltO3RryYBP/q+IaxAwlVwma7Ixy2sUbpDzg4i+7fm9+aMCnx
8hNLqNQz0xlsDODZO+tZMGmD7pzKvnGPquug1qLkUOvW4RTeSxCHzx0LXYlidSAL
HQa9tkKKU6Hej77hRPr9Gr0dg9mf2ylvQ6JBxx9sje7kft3w1ekGt1BpvPmKlafw
5GDB4IW6bKjdQqlnzEdDgZqYlojX66gazb0mV/JXgzHyTAojm6ivk6FaAkFex/w0
+gg0hTjXxAcghQx/yx8qVksM242/HAi3Fnz0/f+wclTs6+FsHo0lRtVsD3VT/0P0
V5RmDKDwvNY55tXFPnB6tktIn4iAuGEzlgTm6bo+/PLLKWJLBN6e8YxVO3p5O2nV
qGwQxRCZtJrnsAaUjxGwAVKOV6jM12lXB4yO1lL9NT0VYQaG+bW8PhSbPGYi9Usg
OQKumBAAo1JmG6hz87fVcfPtI4TS2fZ7DKjY3/W71UTmR0dEdvTJhEBW6x+VKnfD
sqvhJ9U70U8euioXX90eldQuk5T8AwZNvww/ouqwS/5oJA9Bn2tuHyBI9Nmnnfik
xHvXg0KP9fEJNz6OtEnmUDw7isZOcFfip0Ka0kMZ0uzDrmak8XcWZ7CQfezt7iIX
aAgSQ3706SyUSOW8Tjna0PJWBbzEDlFnBPMWQZzwhWB6ahUCgnNoBAUr+zvPIr9C
IgE/krZadnmnWf2bgumjS52byvrhFNjf0QPT5Ar9MrI8jNFJH+qUiaFkgREVxAE4
6UJEd/UOzihfXGzlSv+DC9u/rNBK4puzDiZCqQGbeege7/fIOMog3nS7q4SUU+r7
WZ4CTyqMrx6MtorUSY9QuV3zVlYxIQ4St2H5vy8fEKhbLzrss58pIrNJtQHHomE1
5Sg6cOu++Hp9qyALsu8mUHYSHoiqQkMi6NcS4FJULX5s6arZrriyvMXe2c2KY/NO
YtzgwO0ucLj6u4pHttpuwNxfT9oPWmvow13m01TEuaV927lGpBxZnJjNEOGN6AMt
h1Okvh5Dxwei2GoiR16GVoAJK3+M60ohjhPF0utvYCRV9z9+nuiJEAA/ZYeCZewr
ZkUdBdrcD4AiNmP8+22Oa2QiMq8Cl0Qm4CPn23HiOU7JaOs/wje1vzF0s4OoNeUF
s1PqW1yhtFc20QMWX8uoUZYeux35HVarsRK9uxbqb7RoTtWDmwOKQ6H0FRNRWgUG
E1fZuCeT/PQ3F1u6plZo2T71hDF64qCOuf4YvDqLJgLJYnEEG/S9gUIvd883csBF
9/9kfa+QnZNHK/dZOxHCM8JT3bYw5s4CUTnnlUjMVrKnNQjqrOUB1hxpTbUso5oI
spqzwKkeWCYBRTP9oH6NlSz7s1VrqY2yYvcFyZ7v4qqlFeMY7nPONzGzpKoaBOW4
OVuJHOeCIR7gJfm4Lqs0+MGbd2z0IDzuX6gx5+uQhC0XQBGfdd52hnH4rUqVRlCY
6V4rhKozLWecTkBVoO5bjoMLWk+1idcHeFeRO5/u74uOdDeTDGfCx8Dk4Kw0b6H7
GJOkxOAhyMn5szsnWyLIqCoMWmW6CYBigpOJc05bK4cKimaQrSjrbm8WQzOqlPMj
NWOk/gP+r6xAwOIbC7gXDFfWyYTXsm6umJFAUeSKDtZO+9vZy1Il4pf5Sz+bMkRb
qYSzM4dbb10abuasPhgyyoJzDNpyvmjuCCDGGNTlu2SZZNd45HHEdICtQvMstMPq
4BDE4dP8pn5kMQP8LgXBEJLkwdeqz8LHdBXkDt6nVqRbaK389q38NRt9f6UWH3sl
0Ik1H+eaa8uz0MyPALY04eevEPmOiz6Vt2Bt5RE+5j9njVjDmWz76jXYgQqkl8KY
M5BDZsmZMdnCvtUYkdZC6yaLI3XmyUKG3UgaPIUkf1oh7vhPiJ0dSqxU4kX+mpHB
XIt2rzgqSe9t8DqzmJ2LCC+K4LQOaX6dY4fOzThUwUGAWMeKOxa7nsTIFPoBegBi
KRdY0XC9YQetvKVNLmWeoG5fa0i5NKSYa+ynDs1z+37CKzBRu/MZ8C6inKC80DSM
v/tt+LT0K2ijGRkJg8+Zz94z7k93N6ZSW/uxkfmZhUoppnr0bAz3sG4Wcyi4gkbT
6yatCVJK/3JY2PkHj/g9NkySKILImCkyZCiZJhYAy1YQoVmPs/jW/i914TO26w0P
lmLGn1mbQFLl3TKStx2SWG6TQTDiCq1ff58aFLgucxhDs2QqTHQcBwgUQQbaHLyO
4FnjYRsamU0YKD1GoGhyq8HluJwaz/vDWCMO14vOa20N/rFTbQqXRByxX5ie5hoB
BKuUiIgkY/IARU30UxJu1aIP+GnGQLmMPGCh0Sm1hOPngv8CC+5PjTvuAQsTvdAq
eexAtDLoPBjHCOktm/IoCeeFNZ/JgjUjOzoYxludgeVapC48TxFUokXiRvoNV0+N
PsurlrXG1aIPerFfJBA9M83GOHLpaD9aqawiAS1wpplVNAcxheySLDrJkskYVzzW
MfiEGJF2bulg5Zf351NNfI6cfoj0Y3oQ45IlRZ/lMd9I4hxdh21ycFWNzYIU9zCe
pweUKB7r0vmQVreeuQpV2Myh404IIM77n/mt8DlyT6qeskK6OuZPNzOt9DXyJ7FV
6c1CcEsuufzTWjsKkISbZt/TtVV2PpovGS95SOIth2E1yg3OwOkVgWm0cW7f1DBc
Ii/QRNtcegva8WObulxMQUIL0QWEkNdGhryJC++Aw2nEqhG28Jfmx6cywaKDvs89
hpOsI+dlbPH/iow/igU4O6hWHX2RIOnnqjuuHnEvhRGml7wn4++GPSRLTHYS4Vjr
Q5CEdooqIOoerffoPx80kURFuKL8I86VZIkWNnAhtOSFj1J4UhZjdLYaAr7RL6el
9H/YcXpiMgfBnuG6fmnOMbkQkw3ecDd1uwxQS+3aBLcx97/R30ujOjth+l3dh/VX
vl1JCbpAZA17X4bdVEdukTg1wse4p/WaLwiyL/M7T2Y6LWK4SBO/FOIvgVChZSai
DTHhT8T/w1RF8qxi/zeMAQ+3KG3efH8zhbtK509uYvpd58b/COONUXdF4VEQTVDi
HVSQbLsIwg+l+C/hF+xSZBPfQ+/mUiMp/K1KmzkRYdeSDRqQB/TSr1ClbAnJ1XDl
cGyTYaLdr56QoSD6nQZ4cr69T9XsqZj81SEwJ9WAHt2nWNf45UZOBDhv0Y0JFSHW
AUpqD3v/gROdjHR6qFHtNWl/hxSG2ShtABD+BUQp+A9Jp/R9Uo28NXBw65m2OqZ1
MrbH+HcL4AeSLgOt33XKnwDr1CABsy3y+pBb+NQcxNVDO4bEhredagCqrCgag0Ua
Cuj5XWFocDG8CRtZCvzHBB/63qV3kAw89j7T9Moio/CRBwYkDora7hiZlDH5+Yxg
wS3InsC72BcWAb5gmSFqjWYtLlju3nW5dueJWuevvlLGcvrqSWvlI1lYFsoTk1V+
fgGJkjClU0IEKM4EsHAgfytEVyBslNVwOtzsOrvY6L5bK0i1vUvoWDKvyhlR8/eG
EmCVmuUm+JdfNwyv8dc9SPNFYU9IEdSwOlNQd0IZY2EPqZTPuSxMCkkO5nd0/SL5
fk1v8LjzaDwT39vIh8Xy4uFV9JOAIm4cNNz7JOjrChOwI8T9yLd8tL1SZpmzBMBw
tyCliBNC3om4eUfE1q884/6Orh67qVDyfiOggqwNRJWejt3n01YY8nt3TA4lblDO
1eOUUZzfGlHDe+spEicbAhnW3bK7fsWL3sn6AH2jt3XteVfGosXDFZAdgWCdpVXk
rVwcO8bz1nQVNsX2A6rdlfKJSxIAIr1VU6Dh4BajwEAGbwpGFWycPyStCPwK74QF
Hmu3uEXtOE3BYtSyKn0GecmAf2a3j6uTBm/DYYlJFNgeUgS30tvJSdfJ2x3V+4xt
Fyn+HjETgecv4vRsFUIZb2FEbWVt4QDTvEkaCvFUYuSjb4Tv2EK/z04o697AmOry
4KVFi/l7hSxWs0mqOxdguupxULHfQudrKb6QklqISBMCXfti6y0LjKDBqYDpPHUN
lGzkBp55hSdw62ufUugqArmNlJ4L1LFh+ZHfqDj2t//3EmjAhtstZVoqzMzHRl27
aggmnOWzVm7yCLzGY+lS+4DKhNZnOKs+0fJ4gHykXkJIcEBVobd5zjUIYImAcJH7
LIbTexWsbm7b1MKaMwk70ur5dbL9wk03IH6HR9xIoZxi2JSDO4+ya3V/E5h1IzJV
l3ex3H3S0kttk+Z2Iaa6Gy1vDmou3rz8T//ZVag/T5Pa1aT2lO6Qoy6CxWwcl+0D
jn7/U+1JdcDRV9pp3/KWBHzHq9x20FuqyhnJNcKwyeQGnKhmueHk7YAmkzKfcAk0
skc/hab/nzMeZSq4r1+FooZNofTKh/tiSmkrNakZ1cGcIiXBHVO+O9k15MUDKVz3
FJbWYw3W4fmZgMpJM6uBvEAM6LHZkzxy9rocgjPOsnUEz8UU23iFsdJjlKoyIOOc
Ta7yc6x/iBSycBgmAizPWEfrrpnpfoH7gjWi2Z311wfzIi01QAZ+1hhsgazmQrz1
pVvOF7zFHrNdIk8wIdADzg8vV99OhRr738j8RyJ1jFcFzhvMz5Ep1BSfvmbOINGa
pnDh8LWr9TWWLDnZUVauKYWBe6lFsj8hhOtvYGDkkOXk351OHwjxJuPPAivBw1Pn
yntj40457FJyd8j0vXDU0alD+QSn26F439nmVK3T4Bro9cnCQoQ1YAPZ3lnzZCb/
P50aplLqgI6gpphucaJS50fCAswbTddrMFiA6gTvTSCKqUiTYAvCGn7w4NEQWyq2
wHh9d36wCKbfgnkLIIxtjywUfxw3a+cLM0tRz5dpRrot4gMyqid1DRm9hzqq6rem
kQVv0xKf6AaL/Uy8rmv7d1PYvkBxDNRWC7ry2mGFhKvXr/f9meSIv9PML4+rtrep
UsHvaIWOWCLuYMs0Pm5PmrXM3gFJPFJyzaugDxDdLyymtPmxSdwtnqvoOfWfq+v5
O73oBAvu7XIfByVYGI0cdBG7SyRiPsadXlAhdB5pX2JaZsMoGjT80K6WkvpXlmBA
n8DJxNJdR91ilDnmtG1dG+1glRgQnty/yutj9XqPF+lLQff3C7B1ifO71ARNfRtb
eGCFBJXDojdbUniTnZhVh4iMmVn0mgdcpoxawXZom5qDDk1ArhDogsh1SP+cwgeD
Iv0nRQ/Yza7CfLkii/+xCuOT1IAvWe+TGSd2fNqiYtp8ERvlnBbt9bu2TpzELd9h
OM0zuCs/lPQeUz2cE1CNi6rlUnR0avc/Y13J8JQoMfCeQrJew+vTRtaOXIhFIZmk
jO9f0Gp1b0KHi/p34VpT8g==
`pragma protect end_protected
