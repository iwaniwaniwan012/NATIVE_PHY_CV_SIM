`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Gp3ZlbqSho4cLOZ9kLlPjFUCKOCQP27ENYWjDwp66t2AfeloycD5mQ0l1QmMVbCb
tyOd8XEgWGFlj5Hveo3lLtGAhGrG+XHiR59NR9rJ3O3W0mi1BApLV+jft2h4MLtt
RdT9PZNKG9l5zY85JYE4qVBUUdg6nBRzMhFqkiKc69w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5664)
ifY5WPoJ/xyb1pXXn/ehCXxJv9BAF/8Yhq8as91qtTOWdYONZif7p34i6RV/uvcX
FUGE7C7qQVPsBW2VaXpZo/0YMpKe9Mz17Vb2jDKBGswy+sXjFWtNkdz0uu6/2Nt2
btm/bt8ijNkfUR2CmAhgKr/KRyyc3vUoSto7qdWpgKX3M9L2Pvrycc0Vsx7PBUUd
F1aDvCqb90BvMXmAQemK32bXPNdG9GyJ2UmyCch9TBOkjGioCWzgovqnrhun8v0k
cB29QohSl6rYCrGWHuaXAOJrDZ7vDwNFDejyXj/BcK9oMDIKVSJ+NYJcaSZ6iZWL
GmLW74CtVa+nEgt0UIcIhU8kHs4wuQ6ZEBlLOLvwVK9OphG7huqSV6PBNDl4nSyn
GzrxKrzLE49Upwm14S0KxVhIDqGPHm2hkwIHg0TiExwFja5DawHXnNzF/n5f07Y9
FsLkmd/aJmdbcf5lSXlarOOuyOnECn663syMref5WpdO4yreMd462NaJuZvjGXBc
bvOft0o56D5uqenJ8YuC82YpKGblT1QA50IILReK55nGGoDbFd6BO1G3vp0DpYuN
iT7cOR0vlfIo1o5A78ZD/eCKSZz+UhF9NqHs0ukHh4JzQsZhmqhV9w6KnpUP79cn
oXX2d9EloechLx/Ui849tT47mMzZ0V4fdQJL8Q0SPukyXnCDywCGUiYK80/VEim1
Q5AUlN5tVt3z0YrUQL/hE4I9m/RzE39NasPyH+psV0hBZoXJ2LpCOpkp/7TywYY0
mPYs5GcLHb6tatMBMjIgfal3fx0fMDHH3e/mBGXC4Njl3dj4BK1gA51BZmxAV4/D
rfFGdu1LUwrN/AcQ2Wz59Wgb8K/Z66Y4p9+ZaziJ8PrS1mFfWtpt3acSmCx+P+Ez
8rGb25lJv5n/TigPAmXfXseAwleva7Y441aawS2MWSyjcLVZYI9XQMdjEV+SWqKm
42B7odAGFUD8v3r92M9x3OwsbMfTFAZxhZ8Tun9cCRWm4XTS2EkLENDh8ayhiZaF
5iKmQTiv1EsAz9GAZmpRvldbrnXdoUptmeTKniW5oVK4u2wIkASBqjKtUdkTTgi2
M3yVahaN0A3JU/GfBVty2m/DBUBlcpdq9gOjeg9Ry8D8d/qcj2iLhs0cxSRGpH6M
LfEpMsmHJQZyR8tdGaekZFg16/cGIWdaLTM61waJo5L6MYmx7DIVYx7oYDqnpsuH
iZzF90m4Cdm8K0AjCL//kplf0zB5m5+TsXR92Xz2FidPqBTZshfB2r1gBDFEhUeW
vWfVYrMVaI2M3KC9m+dY+qerSavsM+1wjPKKHoI8Km9+hS4rnK0fleYLy7WG9QIP
eeSVBB83rudAX47K4J7En1Yq4SClpq2SeCMnY+ckXYJQhPgDZfshz1JcJ8SaAw5L
S+BoeoG1G2GPpNTRRWSjy8aR88HDz9fj06khbdEduJO7e317t7HKWlgoa8oFyPTF
qpIbYeB4Df7kwpu/7QvNHCrEZ3AcXqIxviAddfYCiZdynkia2GFMIltVxftorGEe
VS27SVPFcEym5o9YGVKglGagJv1LvnyvtgRaL2fVZLGjp5ZMf6Nwx807vJ5MgAi/
dkk/hYpLf9etoLbxzbjKbKwUI2V28mzPmsL1SbISuIHrLyCxqQFCVabDwugodZaJ
5AkL0R8G9Pv2GQxGJ3wIjjluLIBQKRID1Jn0BKr0aQU/e1uHbLpcopP0Awu4CfY3
00vCCJgMpbp7Cz4VCH0DEksDV5YkKftt18K/5+SGdoL6m1bDmuHxm20h/GSTtcLN
Qr7figIQ4TBYYvzgK9v7ofV99OaIuLh60K+MlZnK3zD4XTqXXgJ5ha+cUb/rO/gD
G6iZPGf7urv0pX1An7r6SeSEx64CdbfjsMD+iFxVeTzJVzVol7xBmWZVO7LRyUVx
5vnprgfpxsxnj/hixlbQPgGHuLBp4c+nMIixN2BNuUpPTK5+7W8KttSiuJjb8tEU
Rvbny0Knye8md4zoSAdIqxwbTQg2MDp/tTba971qFbqohDiLxOzd9Zw9R7VYiiGW
4WzsLKj6UI+A3JmDFMGz5fjyQ9bC7IVZXZuBwe4cfYUSyR2ytWHZ2bN83u0eXd57
paQSjbFdjs4sfCABLxSaqc9j/QmL/l4qhv8JONDISrV/1Lb250lBRhJHBZ+/OXmT
h+Yly3WFj3hi186fZqd4ypX/5dVFURub2drH5ghwqtpKqHydv7Mr0KASTfH6zKU0
Sj203Rl3APopkmGRo6xEgjCzvfPKIDQOX/1Qglow9dy6WNeiaaxaNKB+oeUYHYIr
gesJJ4deeTqOKOaEq2Gm2pdSVjAtXx2J9bAPRfLGZ4Wd3mAt8xmuR7HrQx1obgc1
IOBB8RdsKjY0sQZkQ1efUHX1VOd1RImHcg3SoixpXcmztmYVcOmYnur6mWxycEqs
ydJ+47Tb2dYQb1zmoSLtGLHwIwiKLHVQePR9PwIrTGKpS7PoUyuQetSA1Ev/Mmx5
37VEepbIRy/M/56wU4IPV+lQLIHtCHgX+FP3zlucRESSfunwfO4ETjIkk+YMvPkf
LdPMNw+95w0TB0RWMjWMmoWy/e47iycP7Ts8CnnqQuIgqDY+lTBXKgWRyf0tkFtX
Uzm8eR+ZFEXXLajE5XXegXw84iDCI+ScBwm0EKaPAvur1pECKNq9whUFkfX5pjM1
ZkU+BmNYKTcG63vNRxmqCDwO4mFxFWmjGU/r0jDp9dW8iWGpDhw8TTurHUk1ABtl
IWCicGezr8EwVYnp+N0u3dJdq0Qxh3ULd5MhE8HAoznulhN4FmFp6br1lNWw2wOZ
zTzVBaVq/evvCMFJNBx3DU2NLCLzdZ3d/1+ljEYOWYozApWpjRaUaK/aNczU2iuk
H/Tagx7ZZPp9Kc5V5ymYHwVQaI3zHkalJ5nGMYszn6zh5tbBGMJ6RQ4BVJM31dhY
zoIghL5sB+B63BvBoG1UmKlq2xOdcH5k4f8GxxUAghut+6deUkgw5BgCEaQRu6wF
pKmf23O3Gmp0J4TBPtQkaIpG+LaLKdnOI6ooZV1Q2dan7Sb89lD0ltt6wIMDNeZU
oYrMpFdX6BOmBRY0PaupVer6+IsZDVJnvyw/xykuCP/hUWd/kCugEhUlOEi+v3Xs
YeEJXEE0sKX63G6FMl0fKBaw188aixzwqEdvzuXyDRo/WNYy39M8VUHFdKexRTao
2CtMTpGz5AdN88GKD4q6jH8OzeEg0+j/tBJV1X9uhIKeIHdKnjQtxM9v+GVnAmgj
eKlrKZ2/f7AuXx92gZcPK73d78fw/1vnxMf5SvIfVoWGT7EhSuoTFOj5HxyCF9R7
Qkw5pdCLuL2UY6R383XH5GcqGZ3Ttum6E+UxQwfOcmri/36MAeUFBMMvkiPXSMVP
5eef8RcrqqL4vShB8Kq7lbcelLFVnkyRDWkjrVp4XIbL/KWje/peLmlgKII+A3y/
zM/VwZl2M1AMlBJ+rjnMtPWh1nmiY65QPBAm77d8Hken893cMG7fY0jKQzleKr8S
/i4IhktZmAFID2gYeyFp8z7qNCs78QsM3PDFWcyu9isJPe0Fmzyx4Nc3nZQDHqzV
vM334kEYfwS8GFWp19sF7TVjTz9jiT624KzLqYurOEOIUkmAmTvKR7D0c0hhqylO
w0yFvxc0/jlI71IbXfFZ3+kHpqYF3dTnH9Mnl8eEngyoF0uJOsLO7wH+khMcn3Ip
iirjE7p5olNnOoxfjg8HYV7+YW0tkRvYqL02RML0c+uyMsBq3ZyctCzHuGgsMsRf
VI7SMd27YmzDA6zefvMVLjoxYdb+bx/KLDxldvafRt+4LUvVUW9Ahp29KiweRUZb
bgzCYwh33qXFRamrXrtmvvDjpcdaW4Zmt2VN+TrA8PvcSndYLsU6k0qDg5W9BrCy
wUdFr/nYBr03nt1Y/N65iBLixLKTTtCqqAI3LbEyqsRZvdBfMygCnPtVmHREUI4E
wgCcCGRPWJYHfHByM5BLQfGsZvd8174m3EHJFpKS5SyLXPco6BCK4GdiN78o6Cz3
GWQzOJKWPldzjDR3upQRcwGqhDrhp5pBvus+dPM0c8+51d2wZzNtKCQ6Dyb6GI8L
DiIPCo7JGWzPb/uaRTq9rlUfPwlwIKATcEE7ERc0ENzpeS7kfF4/pqdU/X82R74B
5qPS0gx82TbzqRB03JxW5OYnVb8gwx+pDTUNNNj8awQBbrPSh3pXv4RmG02EY0x9
RoLEaRIver1aQOCYuhLy/OJhQ6q/xPDE2Ng7CqvlAmXA+U5VAwokP/iaV6s0hudR
BtOid2ZbxrwFwYvITOzsgahffTWRXw8OoeoJVZpLBqJ+hopPicgZGXZGG2bikBo9
N5xyW19orbmPI2ZiZQzYm2J7fsJa9jlBSa8yXyhItpKtl61BEYp6eo0+xgDyUw9V
VMojuhcbT071GM7qs1TFxS5TvOz4FayoFWUrC5NuiVYfPaOSHDNqML4OqBi2zS4Q
LXRPQ/AEVTcrc4lYu5SxseWeAwphhyxBTYupWq7sv8GLUCaiESYYELy28IFPzTly
4kuiFZ0QfAoe8ahLwT08hYiQB0q8y+p96mvIHVE8xvDFEErKRX55XVVvj7Y9SsUj
g4Js0VgEJL58AbH1XX1HmzAmv3x0nYzCSn3kiwXpk9KMayMrHKKuixoIKa1kgkna
tWDKwWQ104U6WkoyN60GAXV2l0mXqVb8W7RuOD6VE/Od8EFY0aHS9qiZR4h2CY5o
7g1CujciZjhOX/ckz9rnZjQp1QTfuq2MkdiG+Id/p+sfgLYdgck2OERFVxQi7J02
ENJ3tGUE055OGGuggE+Xq3g/oLpk/16DEWnxHh16uL1rD1qpaXEXEJ/9Rde4Y41g
Y+8zoLXmzn6qtymnG9RbhfwLuNkCJbF/Vdc4l1435TyqEUrNd0YyO8GUfoZK1tyP
tT3Cq3+THf9DPMkKD8UhS2XbLjYl/RrYjgNwcpC0xrljgmOfGSF1wS8rZN3GKqXq
A4jcX/jJoCGPU7dtDH2cBkQLERw6vQ4OetKtMGHVkdWa57QjqdZHn+FETvCMT1lX
5vO5thSgCQXA7qtJ6u03akGioYtSpDoG7MeLKjnef/v5yjfHLyv0kGsXG55d/UgT
KABQnp+2AFiDTLWpRQlDh2Je/6fAWqQ6frU+PZg8xd6/vopakxKb0oGbFP1cL4rj
fx/6aUi3GKgCpaBq5ft4X/SmzW95GuQQCwlH9OSFDqCiaky+wabKPlWligqGrzfJ
NfWU0bHi6dn+GMjq03bznzn6g9TjoLNIQFQ7Jv7mDho/NDhuEH2h0XpmiDqlHDtj
Ma80oVpfAB1wOe5CSbu1psbswDnVbb4hRsoY1xzGEBBkhXYxpOZwd0UUTxorYZMs
QqHAbsseIdUxrS1o1TaMLc1d5R/Css2nUWkD4qPO9WmwTc9Nr5pJR1hFUHDa2JKa
Kyuu4CYI+7eKDGGkpr7YZ66y2MMq+W9jXDujdeUG+RLYBx8WQq/V8na8UBqJbpan
xHLSsj8pECveLkHiCW4yWG96sSIlzWAvGj9GGfDBogpkqVOW3/sPWPGDgz+ixSnK
x4gDtjLAonZMcjyC3VyHPcCqjv9/lazcqItxARloSyCFszg+0N4s4DZfFxZocSEP
kCHAKyEDCx/1lF25tfwAp4MqA0FkihfNwIAelhzkvl4j7rhChAz97amZoYdSSOYi
6WYg3B82tSAN4dKENtYz0GxdPJHM/ZlVkRzKyNQzOiTCN3haGyhA4LZlzywFcNKr
5kIEII6ZuQRUMsRbKUzQRq5SrFbn8wfPrj7FQQXY3jJ9W/Foq4KLfmyMKsc+NsLB
q+MfEoywLiZfJLW8UeYTlQR6k/AJe4Tr0Ynn7N+u6s3Jtl6nTbXXsbQ9XP3I5hTy
mPK8v6296cs1kZMIGXUl48xR0e4+cdy4esD5p0sfCKlGkYFQYi5h90MI3/ZrRqm7
7PuY3F6uqkhDARvBs+klrgj+uNkG8QYBx7wdPeFVqLFlnlMkjyI82MhLARpXaIzz
Db3FDsf6J5tn87fd3tUiqrmrDVb8hDZod+GekkY/gdFxhiaqoL91UqmNtCJcXdYq
3iN1W6Hft/Epdrf9SjXKplO38pegQoxWPPytD2hja/ctOmS2KIOcMNYzyL99D6XY
b5IICYMe/aIiqd437sJq7qahPTmTddMcm28hGhJXQHMsRlxwTV/ctTETF9AElsEP
Yy7pbkCtcHd87F/T3fw2//BiSU0/1ABM/vVF49nLQDKz+SKpwdBiG0xcRewsHp4x
zYNx7p/+j3APr63NNFvc6zG9trkVAqr6KNLtUK74G1jvFG8h4Nxtkl/2kNic9D/o
P5B7UdTEdgsYnWT1z/rwcD0CJsOXh5tAZZCda95NJBqadh7cSVH2E9bB3VAOF86q
bpAM4xvqlpfFZYxz0U1Yk4GdBNG+GgHdFtMEbkZ9A+DZMfynBD8b0yaozkQBZN4p
fQsNdqGXQJiMSox0oSe3JOfkbrL248M1CslFO8YTOrHkQKSR8vPAAiS8DwRRIjnw
b9MJpXPhWgGoqLUof6cGa+y3KOZgZpz+1oHB3LD5mgC6a8Xf9ZvfPYjcBMZzKXJE
UW0H/ABwgmiKck9JLwKG/Eim2bCMIES1uOqVboCmPkBBt7ZahHfnI6QkXseoM5IX
12Sv1yqZ/0aaqMZ1RNb7IHYr5iEnzZ7rROKv18YlBsErrMhg1pT3kR9BUES12sIB
SY/aSw0Nlzj2WmS7lHWIOI7/om9Ckk1LthCJ6wu1bn2mLDIUXj8xvuIMEunrHYEr
JLDfJMLSE6GehSeZ825uWzPXU7q9fXgRYaa4rQXBPbzVtDIiZ+z2bdvjZy+fDKSI
xd11vwtUiXUdCt/CKpTvzPt6vWQkSE0BSO799+yjYYlC9WiK8X4hsnYCJg6gZKUq
oPGhG3i81bJifSpZ6h7hzE2/ihBRkALz0cOusFLtZuVceM/4UIrXC89OVnOAzAxY
7/a1nzrKuSEtiyKD4i4VwHLhBZLJ9J8IXcDKju1E3H8fS1zjx4Nx/+wMSzLFUtaj
esVoWBiQH0JmzExQhS/yysvN+6padsJNuF5yLe/0glTQmeHJTnJAdKs4s4Wtvlvr
WN8C0wx1VoT8Kh+xMtGTIaDlZSf0peYrPMk3z16M07LxMsS5kq01SqXNiFYN4LDo
tFo+wZNNHRORUuAACUH1YTYwH2dcZii/QLO29bH2PqGtYKqHUQPEnVCeHKJUXTyc
UNNCSAWquu4B4R2bZddz9I8pjIy2Sqc88ZLJc3ck5/XuTV+dpYIPzgf33afjqASQ
vgfNQGibpv1ybB/xO5fNdY7KaXYjtl2Ab9OaQvmNyTZvURslN8lNtSBWPio/cTdi
04vEk2OJKbCsgwoPz+E0gMjw2IblMBKGUmzLQxgjgud5OWwKq9Q9e0Y2dqtb4oaC
Ki2AcpqQxx8v4ZLikWoi4RRd6Q1J78lZ03UvZx3Yu8QhQ5FbVNg/Af6s1FX+uquE
dhQxchP4bAvUXkFVuzTUCwVpLmX81JO2JKYHQmW/o80T80xWLiGJVOHIpXQq/CaW
`pragma protect end_protected
