`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HFUlDiMco3RoXQ2G4wnpOzRj1dW3cPvTt6OPFr3rEi5JAPsCFha/ae7Wq+UsSLxd
maGzVBe5GVMGMvdQbocZTLp+C5d7dZtikAwfOcoL9QgIFMDAGgnpJCOXhV5/0po6
BIICINqVNyklaEhOe36CwGtWXeYSBxDzPHNBlINpAIM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15376)
8uKXwygfqIQw3XWnQs93AK6lTPwmutsAs9FJa57o1RSe6VBuJ2xAZx9NhtFWlcsV
UbmqNp+FetK2qiQ1ken352FBqg4KPQQWIcY+KA8FOl3Ze4ZsrR6wdK0BE/lsfhqT
hpIvAiCHfCcqAzBXL1IO+a3sK5maMk80w+OsTUcQW/m4Ig2ssUsQJgW2NO8l05oD
ePAaJan6ZpU3P3eKzKUDfI22QHyV4KL2IO7a3666QJl2EKNlUMaRi6ykBNc6uZVt
/1jFUnLluUWRxrP1kdLmdfkMvHH/s8arXrKVov4WgpunQltTWEHKpnnSYuU/iT0d
pWMVodXi+qqJYHNHPlH6yiGvatwvKgNPvlpNFVy5AfYVyxwe/JqCckUQ2eCC9w77
wJ5qTH1xy7TbVyPf+BIxnglEFGrnScVg2gQYaEl+7ojBudHY42bgpdSXEfgLwPgx
4vLu0AQJATBPvdl7nOqZn+e9aZcsZiiInRllOFKbmiu1fw0d4F4s5RuVi7NZm6Su
429coYRiC3AQgJgRaDzvp1+jl9/WkxfGyZTDJcde5ArU3aLgseQUFtijxtLk98Vj
lB89V7VzqCHFW/4DgGPOyvLaR6nlaelh6utPrPz80sc/PNgzXZ5R453dAHbr4MmW
1gBL3LKvR695SehHLCM0xmnHXC7rV3cw1dKDhegVAr9xmkrbwwrenXYpoWbquw5x
nHjPifaRWlw/SisEJvJdZFpw1bEhxxdb875WITVhZaRsSOmsYnRam6cBH3iOLSEl
MZTJKOV5fqBIAk2Tz9qD8WxXGTBb3kLTx+KTZel0Hj0cs58/UspdSU98fFh3wlsb
psOzdAoDQ/xGIqUCPN83cYU12nEY6LLw/yI/WNSsEdUnA3O67O2Ia+Ri1iv6ZxC5
HrF1LYkKtgMZu759XJS2E0zkouv+Knq3QyiG8YR+KlB3Az8Hp0BhgjfjwiAWJXq8
Wum6pdJoYMfHdEX3px+bZvJpJ0AnArsvduztv3hoqlhjd2wm4bGxOTTrduyFaJ6e
R8Mod6AHVvacoIu3LYCRjlIwY7HzoxvageOcx6d12knmOcK1N+7Jy6Jxd0StoTNj
lNzZjH+cE3JPdinZ5dyQeQbOg9GUXD/i9U+I/d6N68C5wIN/tpcNIC40t4366u+n
r2gP+WEL4/7V0TPHUp6p6RMZvFLZ7DOIby8Z3i8LSvJfhBl+PUfsg31grNudKZwO
WS+NLgD5hVWFFWVuLo1JZZvuvc02uUoWc/JhwYl+w22F8wfuBDB5FjNPjSxKJiJL
EXS9GSzTLn+ImznTePf527zTtobJOS1Rwm02l07Yxc408YXmNoAFzwNPA1v3yyXJ
KJziMCpJvPEYBLv0kGEwCjDkj07gJDkhgFKhh5oIix5P6SgflTTWVLP79VtxuJBT
fV0RZKn+Ggs7GOmqOoYDC4OALj1k5GJBkV0WcL8UaHqVo3pM8k4c2SeDd9FV4U0U
udg1JvxcSGVigoQYKKfd0DsRnsswLjHU7SCx/nsVPpZjKEK/yRcX/LFbNzT7Yeu+
dsqhAkCzecCdke2HHDNR5EcV+6OQ+K2780kMKlAPHCKDu2qRnTf9083S3P7qMI88
XCrH85h50VVeril8AatMpW95dGWMSexuQGEorD6bEAsyPMV4dBEvg9DSRMECVqX0
u27NOt7SUvwrA/HmJFVLl+DdsrTYbfKbBEC4MIFbz8Uug/pUXkjXTDMyjtMj30+w
ZMak68ivslkzHoW52AM/mQBd6MQFMIb36T6lpEvmww4O/zk5ZnxF/q+p12WFSwFo
ofUfvzm1lQRck28Nkw92JLaHCbvYXpbaK4os937CzGtTYTiRU9JKQhwgwVjaqzVA
LiuWD5AkUkUE57XR1gPF6u8vvZgrzbMt66ItPdaZ18ulIm/onzL6RYfgvI48l02J
VZvC0vUX0/EvbJWkaUChZAFKJ3M11twQriX8s2SVRpBx6vPLP94KBSfPDcymbXWo
XUdky66TV4W0+PM9miV11QcJ5ojM2HejlfbLaa8haepTTI3SbvlDmM9Cuc4Il++i
jzrczJpHG0XdXVFsbBBLWHivQ5NUZ7tDiGfF/n8dq4jla3DyoL3QJ+Ktr/IN3CG+
sstCi4Jv9m8fcEZ0G3do5kuM3k6qdTKl7UDOB7GgYtZFMUiFD9z+HRKz9ZbS0t9C
4bOEwTcANJ8PaCLVCb8DI9cuKwlbQXGK06Ds3hGL3JdPZfHlXCpV4l6DE1jOXzdK
tv4OCvtVmhjTMpeshj2PPLwjgkAWP4xAjo7YTCROQlyN3gRW2jKu5kstMwu6Ffce
8+uofEc7M3lbllZOcgJhCedIP7STpfewEChimOMY9E2XqxJrzO0XOpk1qfqmzDf5
BK0LKa5kHnykL3WdMe4haTvuQgKJPDApZL9HupkyWGUGplHuHPTKYbH0sHecXsqP
QJ0+eYu3mckjQxafJa0pERZXBM2TYLits9LitVf7+Trnr1hcqlEHrxFsTnuQufuv
3cZJ3DuBNpkOTNJM165hkKxrzFCIO1swzVRkOnsbEqIT3ionpPC/Md5p4oKXvtUO
qcL9DqPnbKrhL112vjQF6KCdee1k16lVqYdHduAJ/Y2LthMC450Cf3JUBZgyT+p8
fjPQBb3bNS7q59mFQiDJnfdBeYr1gspE7BduC01C2UxNJq/bMD4gHYXkxb0MRp18
U8lK1z+bD9YHf6IIGlRohAwxigtb8tlQFWZctGVStZKF30wkCDTX1LvL86t+MMFj
tSY8aR/4t/HTTOtCusZe57LzARa3+oJ8/pwCxzxTwpRbPJBaFLEFcqhFq2axIo1q
C9buvv6S8hhlAdIT7gUtSd5zow0xg3yEOvsMu2hO0bk5Q9u1NI+7eacMGXeF20k9
UUCnIP9iUdwP4s+kDNGKiD/Dh8mDBAMpiQWVwlpWQ7H1DFqfwkg5O+61OPfZHzkz
7V2Xboz1vDZbjCyJBBjBADh1LIdI9kWyg+rj1N20qBdiv/J6W21m7sXy66mXl8wt
hivIz49NEDai9pgV56mQp7Eot1keCGr1i4Shi00fKs7zUHl3AmQtugfqYhApGwCB
tYtxK4cL7ExaRiymGdjZQ+mC4tUjoENZkPoiFDq9KimlOGJFRf/9ruyuKOQXaeK6
eIROppeYOwbDK0Va+4WqGW9yveFLFFUl0KyfQtk/KfeByE80t8a5wZUcmGsAyiBQ
0cKVdxtVATfFo+Mc55sb0crFgMSGMLGjsa/n/momx1YsflcENoDFFGF4+TwCseuT
0oHvD6w+V9Yh+9d/urDvY42kX5zHdMkTM7MSdu4tnwWQy7pU/74GAQqFP1UMbKgb
8IzLg3cOfPLGY4FSw426Ef1l1SS/IQ8RY0VvsAWRkg+YHG9QWXomgf+Vs4Roh9rl
bEOfnnSaUMKnKdhJnbuocVdXvz3USgok/vIKROEDIF2YAtXpbHX4uZVyMv+3N6dM
UlWnhcTiYM92Yf49FiZ9Ol0mJYEPDReKjVAS/z6DVjEUGp9ivk3fXGoKgFf4DEWK
s3oVMKcJaLaJyU/whza4E5RIWwR2zt8UVfbcAHKx2vJS1rusO+lLq/qV/QHyXFn5
F7ZRQFFZzBzT7cBXcAiOIUr0T4Qmao22TU8CeUkTv3GK/JcmG00sQGwef2BcRKdd
V5cMiv6g9oZW4NaFRVzgnTGu2N57tPcCLC4RhGs7NjOyMF8gIhymOFT05euPWZ4H
+D2Q4v1JXTVWUocAeo8+Pus7/pczzmeBc2r4pGeOxB5+foyqiV1BUiMbA18yCg4x
2PM6ukOXjcfnp832rNJUJWQ2jX5EssehthLO2iZgkgx8V62XbYJDVjKH4BkNkk86
RfaylifxC8xoAd5vWIPP2Ohhpn2z0ykGESIyMNYBIhnLILqMiw1CUifFIPXF1QTl
TwrCag+lVszOZ2OyAZW5jmqOc4LHpGAcj0gCjrZu1jXMLxcAqVVVauRkfMZhoosr
d5ms3WXnAGm/BxmNhKb5gDGpyYpSPDP9yUauR9JmeMRsqtIzyQ+BpLnz4noMSoqm
oWP7xje1vfAbZiXaCstDHg1jCT+mN5bt3+oRrUtRVbqfS24eodelZPBuf3iP9NVR
mTuNnphjPmDokEcG1uCMOZheVmsGSZm+VluUU77ruhuDubl92Q+5psufTfWtX6Rs
SBEf5eZ62fbmfq85VwR/iqlqr1IHo7UWnWQFy8Ndk0e2+mDt0levljElOK4v1JW8
KQrIV8BaxDt0MQ+9ZE9WLrrwbAUjI1jUM+5mqnEpA+dzHY4ok+Aiqo1jKoVR2PFM
cpmQj9yv8g+0UohRpF6dYnA28XQCGxwyhbCmiQuSEsqIXNYriQ83W+Uutf6Zr55Y
6gShRyoU4F28W5eGnaB/ef2Mcfp/uG9SjCi/QnX/lYyiTH1UY6niWsnteEebMhIc
iIDhytpP0QseqP+oaORFu+YhstgeeOyhSf/vzb0DeAIoZb0ObUdSXjaGoj6gdBoB
4nGJXzEbuaX/RFA/lcFQn1agD2kqRcmPjegf5rox/EnIr7veKym8YYrf1wHh2rHG
xWVRlr1+Lgg7rzo//WJN8BIEyADcQtTjiCsPeCKY8gmxmP5rtVJysEjJL32pxbBx
bL0iU/GJ2+gL117MrhMIlaHyGcNQ4bSGR7LCkjmpnPEOgeGsYFE6IdnLswV142dZ
crOmBaWSjS3ul+DYA2H3Sp1skvW4czwI5zNIVyUXrf7Xhg9nLvuQfFJtOU9RdyGy
fa9vj38bHxjN+Rb3HyYuRQlSBcSZVKcKE9mEIQtMTp1P+9SVF4go0FQJqTXrd/Pp
w7niGFLI1zr3TkuXVKTL+hrzy9RbZLOXYIDsUb6+KL8Kyx7LTWRPLr+3s7P1Kqvg
pWNysLrW5Hou78r+NP+iEX89n+Q9VcOOXBCSP7lZs793Mn43oA5aUWpaLz6ok3HO
yJX1g3N10Qu3ViZZ+O1jovxb634v7FQPa+oc0UWrrp7DKBMN3U0kzPEBb2UnfOAy
o48CuqnuU7vqNVyeB5xDr2Vq11Zv3935EyldHfqYzDwWSQToy8Az0cekM8yROsKf
7V1Ct2TpVw0Wx2FNKI+gPQ9r/SraGeRZnTFQU0wQcvhE98ZDLd1phxn1myJTCH7S
FPZWQyTjJdwkwUsO2kk9ZDziWDKb/7u5VpUALOrgIjkhP8FCUevEmKddgnukhLcX
bZBnEAsF5ntDpuKQl/8Fj7+lnP/OhTIgQ9UywuFWrd3goyY64jwsotJZHk3xsfjv
TJQCCXsf6/a3Ari9Dmq+UELlZLwJjOGZtNwgAaCT+ag5u2zfHTVDgxuJM+ziH2ri
LdAxcvd/QjLqZQ7Uhefj2mTYiI7cka3evQyX5Y1maOwcf/rP4Tey68kskOS4vXjf
wE90AqJZkLfeVmDjqnBjJM2ErkD0rSwvTA2kdwOag5vLSk8Hq+oBD2PdC5CS03Pj
6Klh1WgWo11oe5UJirvDke7BDh3QVl9dXSZuce5rxckfIstpW2VVpyF8mEOaPG6g
a9yPsggp5MnN3N38fXfgA+xGsCVcaFKZ9quFszqRQh/sukdiMF5HMQDyYf/Q0ldk
DUBvdMncp18c6lbFRXcEn8Gfn+pCgCjnD9kFokplmAlC0DnHWLquL4EhyV29+NT1
rpKfqC0EdZmsVa0gIT6WHSNHxhZtWHrFCJzmU62uOt8LVQZGHy5HAraIwjPZEP+r
GP8eMD56M0pIC6nK8MIuGJ99bq8CCfQ+K1oxFxgUWaKPKS1GedghP3uoI59V97yZ
WSs83TmT0yKZtzAiGZO5fCOU0hsCWKEoFZk/3XgoqBIDNUXKFs1xPbhXxf1ENnrf
np0vhxe/40iYezTPO2JRGt39i9q9+e3RHZPta5B39xVjf4d9WitHO8O4GrRHn3IO
Mfd3WbwSEOJVstIZt8ndT2vjJ9VImfQxTEE+jEnL/oqOhNvcg4dVBxrYqR8XfRi4
17PhxH438mOGIUaLc7L2o2DKrCdJxYpNGiKLvMogiwr8bf/MEAy/WsA1wEWSKR9I
Rykh1it5RfZXx1Ypz43Vmw4S13+m4r5tPRDSZttTeRGwKLRvkoBihs7BX6/1ZEvL
4XR848u9+O4rmBHCi3PdnQoW6hPrzMrN8kfIBl6RHxXjkuLxD475WVbyklG/BS3o
ktEchV1WcLme64iBJsSfB8EkVUwhLG/YOhqe00Gf94N+8QKNYAH4TUz2vVX0OkrW
CBKhEsOK+vIPGpFiaamqoFpCluz0bNis0Cd18sjbFiKHYw9glhJ0zAcmLNS58Om6
+Fdjm4AHj4rmfxoa2U4G0HvKLuTdvI42bkEHNjv29W/vxKeHyxqHTeRDapCxeH4A
Cl7Bn6bXJRHnuekUfV+0sdL1hmyLW1loGmhnIzfrgRNoVIen+JK6hNfFgXvJavzR
Qq1yRM/T6pyyGJTp5bK3AZQbpxlO4dRBo7muLWlYMsHEoU3xk7W211fyT3GVhw1+
Cqbfcpzu9B+59n0TNQhZbFxP2/JL/HPppO40SXYfUbTvafyXKiaRGwZAHU6hZw0u
ruYOqqUSPmRdYPQfe+TAQIQTtA+Esm4FEuI0Z8i6VggRW3p1xK7uKqjJlVvJH5zn
PThaN+seDuMdJQFGapbq+oUta4PQmxhP58y1ukjAzTCBDAiZ0Z87gVpdA4Tj5VoI
+c5/QCsLZwYJgMfN/UW0MYyoKK+rFfsAOGQp/2AGqY8AiBJuiow+roAJXsMRb0aD
O1UZwqNdvJG1ErgTO7wjEk5VJHhmy3UPaSYWGremplAnl2VY0rwgheNFoMrXo5Xj
tqyww+xCwzcHg51HKg1KvU5TSe0LoJM8Qvo4pi+Plrl++Q/6sMWiyvASuwpAexFP
bsbIQF4zrmE4swM+nSdYnrEfIoKp98UjTEwdkULY/AZ2/7CqBJxeIRl+uXL41H+C
oCKjcNmsYstqsOXTMhmTnH3x9TSMDY01XykNjL6cu9Fb5CH1wEXquuLaVmrCZlDF
q98IlbUcGxt7AS8NsQwtVaXphavIjdCr12iwtFsw4EqXPeGlRIJaUiLfbeXosU8X
EFiKWyYg4I6yeOsZytUA/iHPllGocfAZbanzchObFhtxu/kw5PGLk8QpG8L8Yf+J
lmrGLWbFH+7RKdoIV5MY+CjbuO+X6sQH500XTvkdcQQQmxwsY2dg/niuD9xX60HC
bHGRUlJ+ruNkDyTha6inc6/VnfyVCt6qNi7H+ZYpCuJf+yACW/hZbJi3JLarx3Y7
O2dbPe55Ua/SCMBlbUSc3KRi1jHVbS41/6FWcEq4sLG1pfhrMHs24Ffylm9xMdOH
o18kGL31R7JFjBske1vMyXq6vq8j5zq/Cp+d8smCvOwl06FsCL30gZ+oLpmU4RIw
y/lYOBu2qY3hdnayyDYMdxl6g2dP+MRk1bIW/qmXIayRbyqWZ32ikDesBrWCZZax
OqWGGXlEucikbHEYsdPdMD0yScyDFXcGibXtzSbspMwciE8IANk2XW7cyDR0GTey
CQQMqCHGxKMYUTFEIQHo+Ngh6kgfW+3Euq3/1oJALbKoAaad2O/8/EHQ4kieAPUU
RIEms7sEZ6lop/hj5zIGmQeVSjnrnNLm0y4+rbXZQKqkgFetPqyvkhO24jMgGTPA
km1A9p7vIAGqTypadiL0fF4QFjeSS3ORnMY3ybEWYjmUo8Xl7G1A6HR0xIABJMSU
hnkVjCheVyWayFoMeTEbgmUWUrMAbed5k9qiBM4kisPzsImgnN4xcmfUG91vw3wo
xc53zi8rx3U+5rO0ydug4Qxd7n9IxaUbDBbhwPzFO1zp6XiJBgfkWsjzu/hiVq9z
GToxDmr7iqHjNqPKbqKBciq4kOJViY6nmnj0UC93PZrNxDMv66zWP5kmRfScXxN5
q1ruSu33tjr1QI83MorwEMiYg9LHZEspBlo0/1r7E/ad8kdcqJJoEvW1GbVPjl80
H8wuj2oIVDtdzWuPUDbjxv/3/x9zY1yISw1m7DoRRK85zsxwgcVNvxvhF9y4U4e+
Kt97lulF5dRbMBhdG1HVdnJjCY/RiA0tnQKCAo53STokzr8FfL0EDtOUVvqV9HxR
NQe58zDWpwKjBhqfMqyqi/N1j0EpvyeuT4eIAqywlNQIseMKEjZI1qW0ZcF84Fec
VFiAiDl/CgUShLRdQ0TSgxg+0qPWhkKRtHYhFa5aqh7mg8SlIijYv3jF0ZxP0D/4
r6wbwzyhy7JFjthr6bCOCp4JP7qwl3vVcu1TIVDGnOHNdaRkeoF4B9f5l0aGstqV
UwVNgNYhSeZXWYeFQuEuL+NnyCGecJFoL+WYcUiDcdu5G51HSgrC1P1rWR+YnLFq
lR9tmi43sQ40nnaUbDpZVwb8JjlT7gxkUQOz2Iu2pnWfrPXQUmDG2XDOFbnsWFfW
nD6OP2ILMYygkKcJkBbnl5tmqnRh+kI8CBBAUWhC7mjTw4JCZ3Yswd1l/aI73J4S
1/w0/rXttG0ASDG3JsEe1rnqNTwurCLBZSzeHw5s2MnyMCGs6QzbBpQDDCqPr/JX
uBt+P2fpwMaHBeMMIi1ck6fIBO2xomwzMnpBnwXWGMzQIqoK4ItkIFyNQ7l8owzu
0Ajsz3tYniJQ4QFVbEoLsxUJAYw3qKp57PRCGA2Vl2oU2gC4YH0z4/TALpfEr0WM
oALlp/b4J2rhywzMzxayYGJ4GqDPFJ8mei493F4aJ/rj7O4uqLrVYyJL2hEx9eG9
ULK3oTaQJzUe1U309Rf8V0jeFSYigJ2w/lhotuZuzL0qXEuzH5/GhVG0MKIfj+/0
dixaLYZhUCLbLG2fKV85ku/u8QjT7NBnbPGJYAXcomg5cpobkxay+3MwFJ718PQf
355jYi1RUVgGejLnWcr1VGwKsBGGkH9Kz/7ektmL1a1NP7gz9C09Hc2FEZmOD0H1
8nuUgeazOEM2ROYZDrmXemf5MiapU17yEQ1GIoodpMk3bfDDIHPcnYu8Ay8zL/Dv
uGYpv95WKGxXtLGYejVKYKN5U4dgbW1qzXTABfBTItCPieMhLypeobO4V0vCZdBn
ZyulmxMBj877IGOXGk+tggtX/U5yI/One0AkYwd93cXzdGlwDgdCX/sxFlxAU1XY
l8BbjuYl3mfTG9tMRy0rD0vr3BLHrTzfPkI3Wl5L0SbGTgvSqiPpElfGGtmdulIQ
O4XsMShUOPJJDW+gYThonS+nyGzYuiSJNEwSvXUWh+r55SZC5p1qZ5mbhcIFwavm
qR+MficYs6QkzUdva2B7DbRYj8k2s/hONy0vxBUKqTwVDRlfmy6oS1hHHUC4dBTY
9mUKoEJszsllsRKactvAEp4M/0eETDTKG5vx+rzbMaLV2W6DHWsGqGvtc6/0UeaT
hlsZOoHjdzJLv+1/TRzu2Kpa0TBTvbSwOipI1EJD1qnv7m+4gF84UjzZu5VU0lJT
zZkoMh1bHtPmCOv4r9Fc0KLSRRoL4uyAJ5T+op8sHN/MGROQfl0ohgHBfBfJxoTG
Q5i7BU3QIQGf/wmwU5f62HrA0K60cZec1YCGE7wCGy6rtYicRNJIjwcUCVStRyx3
tfuMyTuBjqyTYq2yXD/yPVEwV8IpURp1GxdAE+iWS2bkaX5BPRLnIqC6sgDE1EwQ
7bq9vCfDRsMEKZpqL/m3PvxdQ69jYXfzgaSbwzd6yMrpfcvDSGeQSzsT0PTdcakW
J+sWhk0HETjcOmPNQM8a75uiwIISq6M1lHkxkOCMWmJqsBDaqidx3EVpeW9gu3oo
RDvwqcpwcWMAYI37GmiQ4IRr9GFKtrK9koCVOW8d9eWu7xaUQe18iYQH+wJg2nhV
UiyoSAo68igjh+LZaO6Uigqy93/r5POfeMjv1FXWP/3t4uPn6b57jzk4B4nGQHqn
M4TPPZ9agkECVi+q61w43Y0IjwdIu+3ixB5pTWVGJUmoBn3D5+oHk9HQ/ReykM0C
+2E4mtg3BRKB/1yrKEqUfa+MvHFz0ixkvrOxcXBI0VghjeYAAWTkuLWsBYMR3G9t
Ge5js5mTjyrS8B23VezO6SfsHbanfT5tsqUqwqZ65wsTEVIzSJvW01X22CVhH17N
MLBFvXtKirByO0inqWzDGLiG1r7Egdj5VPjSBys65Qn16ghyf7DH+ms9RHn/204u
ThfCUEdtScUS+4s45p9m5JN4loXJ8bts74sbUDuivPx8B+yQsu85mPg2zNqlqtis
bDXPsUF1UvockjSzO9Anx0eyi/Klou11qqvBwkBb/E5GeVRfaj7EmkXNMvvFGBpe
2eyNR7MleEkAQuaIv8YGrDWoRaq9GsKYbn26q50j7RPMDyN5GmZGeHnedavX+HOR
omW7d1OIOaeIylAQnKixS5HmPOqInVS2WhCspT6gxqBdsCBgO5F6hJSu2BY+TFnS
bo8+/h+Hbmnt/opysgonTEPDaZ5uklFauhcyGdRMD+FzvZZ5/2mC5Cnsl3vjnSJE
xtYEDqVAdS2y5s2nj0suh1zfnSDRCa1iCOgkGRJaafHb1DvEIT5eoNL41qI0uFB1
+0xemBZLoM1DWkHWkGPnzF+fuQ7oHfDlbrG9KeTNYRzwJpzcXjj+uuFph3qslqqi
dD9+2d/Yczo8Yj0OtiEdOOXgZVHXpoZt+7Nx76p02gouusxeA29RlzhMuzM6tLfX
NkBwCNk5xVBdmnL7ob3uKgHEDgcNXApU7S3VmCyr+KZyi4UPRzWCScPfj3w1pxB+
wWRcQ0K783saWt2Nxz1VZAvMO7TsFOeyaf3uT6UFLByGOM4XfAqNLw6pf+J904FU
RQ9sQJQLQWq3mITSO0AQJvDOkf0uuRjN2susnn+GvvxexZz6Jjrvc4kGMg+raedc
cPIiIzQcSS7I+He9skBAOuLHm38kRjxt5ccEbU0ulfGNb/WQm/zpgja6HzNKI4fy
PnfiHnqmL7A8WSwNGSF2l0RogtCkjIhHd+OIUezZSxhdS25SDdEPa/x75Tmc0YpK
4I1taDNMXpgh6kelMhwCWk3dDAo49p8u05073d03TdNfIPpmsZKyllxvgST8jqjM
FvpuXWad7YqZuLhHOgcRcU9gAVLl716CF+FCV4Zyaznp0+xKwVoskdDofsqB4YbU
a5xN27QtF9vtYjqN7b+ZXIhmoY5RXaBqr0rRibUBVnaU7CqrAyds6UvG6193l9Ct
/Sh0KnyNG2eQ4bao9hbOS/Bd0rbG8aCnGfuIqwaW38yqRZt4uHHVLPIDAauSBoME
zffPyECC4TPigJQkMG2OQ+fSySKHa5l3lfrz/OfTLSy62PFCjiGlCn1xZokFpUeE
eAOADi0Mo63UYYVf7wNz57UlBXXhnfWaQGHlZXorGDVmITY1PnM/gSd7FQTBDGcJ
nh5O2jxBsYDXBMhJYJ/ObmT720saq2yW05o/FLdPxYYmpuXNzIiK7aGPoODL2Ul3
SrWR5YTFqxMJa8Li3LFHcqOePukXpyuW9Xt3URotVOcFiU+06Bu7a//LtxY7T98Y
FwdGjUH13XORo857LocL+DkiPeCUMG0g7Ynm8OHk0uCJrpYeYPFIazmY5QGvXu3B
htR6sdJ9iEbDyw3Sa6ygNb9znKk9CP36Fy/B46j6TUFEVvoybTZjqqk4qJUviPL7
a4ADMKkNKCbP6kI3AKWQzs8UxgrEojpxzIYXYIoi8c18WZuKlZEFGfjIXImoEWrD
nwnR4CGTVH63M8VP1oEvJuvDHHDWKh1F9+W4KjDGc6aY9NsTnLu065fCzpusg6Di
QMxc0XqV8v4Ue4tGgSemI5xP+PSslUvKEOSD8JE1GX6kI4HXxpfqbV0CrzXriUd4
rFXKJ3DXdM7rSL63HhrgTVJbRmt9qimMG6p/qB5hH89n5mRGbB1bhFcIN7DoLN8f
RwGlZX53IVeuw5IWw3c7/VMkXPSln/49BE9FPTBMxZ4J4jX27/MVsyS5QUaVlZfC
tzMwFSSLALYGIMQCN9j37IZRsIhf8omdO4c3GcPw7VQoD1ZhUq7/cpmiqfPBDsoP
/osEfHiTtVuS4qy62MWM1DlBt84/O9Xeeop6UNeA27d+qHANiW6ymC3GWhCwzztZ
EOWVKrJgO+t7L2Tja0Jw3+Y1eEAmms7rtpTU9vmWjcjvgjWox3SF1kckUUsQVUUy
zszJMDG/5YnZ3lkWEoAzarELXo8UrNIDuZucCJ7H99JpHSrBimtrHmyX/XIWSByK
ildApiTK/fZufEBLOkVC+KJJosJEY6C22Mq/wy1cA+1BRNoXw0MKaG6E0POUuNgz
rO5Fdvoct6N8oV96inMX3kr+ARdK6OBDwI0qHoHNLD5giDGmOKktvtehHP5y6Khm
EyZ+bUWem+Jsp29dC0AxnWytQJXonmw5hPk7WZhzru/k1PeKH/nDZeHRAoZD96xX
OQYCLUnzK1sDm7a26m1Bacqsqu+ytFVLvVCxkZI2v2okCae1hg+0Ol9D1F0TYBmP
ed8nmKki7LPTsI1hQMQvTsW5ol0sK7jJnlc03tz+xn53Ed/W84IqS07D7K2O4m05
izxsH6Gt9e6L0DlofRSt/hayeVpBWbC4/4QAeKEnHxyhq1gCxvYScFa/JgqMPShY
gLWy/7jwfCPkFl7ETC+M+jslE7FzT9ocNca8Th/4S0rjr/pOmKl7IU/1oMizw2nX
PLC8K4fzekf7EzwoJRKPRJE/QdWGjVMi+7jfa3Qy4rZyHLoI7+Rj2x3wLxVf2FbP
uhOMmJUoPCdumE58MYfZCjdV5kdKbAxtP1yl6gZ1ph3lPJopJRaI++oZXdXiirsv
bQIafgDsS1BLXkhB0fXNXGnuL3jSRjDq9JVFSCJEyTddVaAXbfY29cbqVH1OkXSV
jw+2Ene6dOzCcWBce9kudKMt8y3GCbmVST5RB7BBY2C5qg3DZWQJwEB8pdvkVLBn
ih4x0/kf1durf2XvCWOlheEr6AB25HfmRVeOERGU0NLW4C70aMeKFEHeEXgbDAZl
PP7Ik/1DjyHY4gFX2PT6PuljlrUgp/lEgfwQxrH5ict3B1zVmpdQN6RJPZFgT/dr
Su4GhGvGVzv/mc0836nXgUBH32QaMIvcLqr9AzdEoOl3xTiO3yXhp9YcFFZu8EH0
dG3un4sTJAX1My1V9zSJukgZcL+BSFG3MegmwMr0sDrBRUGYdNPw4q7c1obTHEvn
ggh9kToSRTxyQKWGz6u3yyPb8d9DopN7v98eFV9iBvZ2ZVD2YwptkhRViGTGlAze
54rUI7Xpa92M3hJeoCqwqZhFpp7ICg9T6lJCyyBQvgyswqSrcWeDEAuhVfqMU8fz
PqQn98r6OO0JA9naJts+wSQM8YVK8fFa3Y9DALrgx5LEU3/HW+z+zxgT4DW0et2/
rRjWnMYX1rX1pSYzZwgoT7B9xaUlahaxu8wmbTCRreNxj8WaVenX2RyBl50nhmRu
g5qdqTZFVrm/XadI+l6FnNjdKVVtaVDsBWjPZg8EPIS8hgvOByhmAci9UqVtilKK
s5hZCM3XdUsNdnN6vNu2SIRtknFKw3y55ZQf3OfUgfJbekWC3MVVcVW2+jKPaFZY
BF8T4WZIm0R7r6px8TIDPGIGQhMyLmqeORraOF3EJCV7kHpddtPuFG4rYn9gvZav
sGXz4qRmQ8bkI4J15Rg0h+ZbAsqG/oplm/J0Jr1bQYvA7qUpeoqE/4GAfefPRCr5
/SctioM0hM9BNosFkfMOGo2rrbpEoVxVAvKwA6a0rgN02yTY1VhCRc7cCzYJ2ci7
RUGwgv7LET8Ofqa/gM2YN+eisXsgXrsa7esaTZa55zRx1vEQHdZ7uccRF6Rvv92c
w2TYFeFxbx0fFSpQO4IZSfHyQTYZlxfKb6HUcSZ7N+XtFGRcu9wXKQqYc7e/Bqvq
IHwUKnV53iTKTIf39AxM9iWMNJ/YVvEc0jDiA3aTQtHHm8bTtQQvT81NG7mw67my
ytBGUdcx+30k0kjN4nhETtOKpfD+ycRtTJBC6U1wopiepm1sJ09TXKEv6dmY5JBA
cuIqXmcTG53bF6yrUPXhL/ic4WZiz2/j1oQF+6z15UjElausT43QmwhCfsYernO+
P8CBbk11VjqFxm/Nu9peMjaXsgFxL25lk8Irtb/licN0n/ffd4F38tDmvX1O43Bl
tuCFY5RpHOfONuZlfyHznFAv16SouQny1PYcLLKQIBzN3mpP9Qa1VGwqvMs2kRyt
VHpayUrKOCh6HHXfjpYLOapdUYzBPW+n8nkJCkF8/sLp+rl6J60vndtFx++UR82b
P8DulRjl/aFtCsXgVOkzSFAJ2JnYABWXu5o6p9v2eKvmX5pVF+tL8uJMpflpwjqI
qPTVLihpuY7XcHxRGBe+VhpWVgqJ/flATQC2EV2flOdgv2sCYIZEYNaAsOZ654fG
23AxxjJPIngD+7SiXVFFG0u5iNcnS2WpmE7JjyznReP7bFawFMaAjJJok5jkomdX
vnABjO1PccRr7iY5ViRkHFATEbvBYmwmpSbA1fur4v0BxDeVD/cQDY17/ZgILDUh
VdC7j7BqJa0QtXU+wXn8Z1oWdTbVUxRekxnougScQ07EQ0Ch8jjArGOTp6w2jVer
Wwj9GLDW8+dXg1bml7YaAAPxM1Uzv3/LamJjLJ2OPvi2IUHcZfZqplIRAef4O4nI
nIdIMvs/YGLPIV8VrIZbxsmL6E9hus8CZo6XZk9xSlun3UoSIXTXO+bwU0p+gTGw
DLJNaMP91fD6qABa17pgX/nsgA5kQbbCA9wL1hOP1DqCXOlyJVkN8uTtc+nT91o0
rp1EUYGKEn8rEMtUVXslSI/IhqSClABMwAAqVst03YlXN+xWmQWOtaseDlctcCn+
Z1ck4rW84y2yACynVlpwT8x6lcExfDN27vzo6QTP+36QTKVk+ujNL4Z+KU2tZmHu
iSD8/7UCLf1rh4GANkh7O1gquEPmsy2phcilxEVmqzGEYEnVOpcJgKt+EPAApl0u
5kxN1lm7gsNSvIKlwqMXv8Ddznpgdf+ystHrnF4Qg/g7G0/gF6dO68vfVNVJWDCd
d2yo7LecbtEaJk8HZ796oE0DoaNiRw53hjguNvZ3+DM+UDfnL7T3eZ1xrOZLxexJ
4+qxbgX8YxW0nCfhuQQ7TbGZ0dkZurnxqam9/TXFcrSjCKzVRE1mwJurWEFwUlTa
v7He/twGcM1Y4tbvb0fMtl2baL6c6Xz2KcqpWkC9DHnQmmXY4cAtkyp6b34W1PcL
gZ3RHUdv/LNVhuf4pntqGHb2bu34+YM4ksJtkrt1bSav3FH0lA0vzzUNtu6zghve
mogvI3xCaN6j71DuLQAKa9ARdsRdbqHLT0DcvIgdlqYVDh3MgSTsOJ3K1GFW/fq5
Lg+2hLgkh98JqkbtgfQugZZ9lbXMK1rTb9FqPf/aJKmluQJWEmX+1lO7Zlzioydq
aDagS43qEQPcIa2YbHGbmSIQdRIwxc3OxpM9w++RBshM8hOS9HfBrmXnalcpvsZ8
22+8kf0OL72OCX0UlPrBqUXT//nX5y6z3YKrzMmrDopV8zui3cKXBB+3KQka+OEJ
vUppZX5dAGZBUKdk4MupQvcmR2D9ZREC+Vwgk5Lc0e42rJJhAtSJ8RgSCB0dHNcC
D27q8sOdy8ecZiQJhcGJxEuyBsJtxMBpmjzXAF+l0aBSbYpZ7eBC9/6bptj+hXam
/Hzn/x32fXIl+2ouqB6m1xQPz6esqaynGqSp0j2XDxdX/br1OLz/x05d8cVbG8kI
quOLW9ITQKMhnWQSKq3dhQN1JflKJszdg20nk4nC8WmuOrkV30C+VFwS3ulu4j8f
WxdSI/dqPFw4BDU8K8szpyitdpRxZw5cpkoyhMs/BiieR7cnHrR9JW6xp662QLaX
X54HZJACZOjhEaPvskLY4NN9R1ozky7UQC9sqfAQocQzpS1/8jF7W8sYggTHZNOD
KzFlvVPKJXc5LFWUVElD/bq8qpoRJMt9pwEsyJ5kW6xL7l4kU9AlXY5oaB79q1W6
a5O5SR94CxvRWq5ho90vTChEhXLWTKk7k8L+Vab4uF5m1fnUAnIE3OQ6dxXdTmiL
VHmjkNHa1e0W0nTZRzGbFJDABd+ym8R4euL7inCZ+6Sd+uxtUIIbh4rBd5i3V++T
nRJdOH8b4HEedHUUUNF7XvvE3JoXZ/x9Y8n91rFnd9EjPnsLfzO/Arm5pzNUjZ15
xn3lZjU+PAWdKiLBjoPmoAEVWYAjq8vGQ0W9aWXw8iFUUtOt2/7qJGOB8uqltZhX
FzonCOYEfFC3BPa7T4a4bMDDmOqmwxJSLuvRvTP1z3UKQZgkhnrACLxu1Ilp/Utl
m/BPOoHHjbew+1S+2XR6HlFh5RMzNL2b0+Xt6E2FREd6CE07SH6AjmhA7tJ5L6dy
HV+isMJkbOItiPq4SfqzvYgSONEv31vj5Rsr06u+jUcx9w3+r+yCgKllkjejvZCX
pHDV0pEUM+IcZFmWO31vVyfvlMV9A6cxCO8puyqtLXAGvNsVu6AeuW8o/t9bvu6G
diSZfh7NvUjo/PgeNSf3jCl0W4XtDAMWWvfyjoxj+/q2Z0y0uIv0aw1Clypom5aA
1Fm/dJyHZH+aS4071PVQuex7K4RA26+u/qVq1BY1o/whl4JNLsggXc2ewTsVD0jM
mt2xul/5C9Nxcv2PbOebu3gx8jVkQmEkVjOTRN21KHp5Hqbkaigy4i4nwoaacR+J
5yIFUeR9TG3jzfgPGEintm98bK8ddHvKRgOMf8ti5lAdSNTuly5PX/IeKAcqRX+L
fyzh6UZFwT7KkyTRX8vKIUp1zAq0MJHr1RP2TeIW475Pm4+gFS69kSYyw6YlRtOL
ROrenaXEcv9DoR5QJnDu50J5GKjulZnwSzATXDkF24dEVyi7HyjXp7X2umC2vJTs
CzG/t4CdZOBInQJ2UvTl3FnjuA7EG3VpHC5iqiCkmvWGeTzZ6BmQrh/InIrdirAl
OIEqFWGBwGFihb0BAJL1SFRdonrQJEV4C23CmkjoqRvK04m/2FwqmpZfWzzg7KTN
yRrqr2zeQJ36qvEDsSkKu6n5RaHzTlM2Vr+wdPCS2QstiauTEuv9xjtO+dBlMEji
GjWWEOrqmmvx7CfRnnqbFybI/s1qZI8bWWU36UNLJSQ3Pspz2tSAdxPYA+/Z2lRr
73QSm8ggUcKDdYJHi9kSbdrtc4uO3mtt89Frb8pagojtB/mlC1HeP/GTo/+8jBUA
tBZzLMfwWBJCpE7Zwv6NOwWiW6XOmmkYawNQr+KttUumrRlk17k/Xe2X6r9s217W
S+23zu4ufgGmt/2o91FHCHFPixCcB8JUZKDOXeNc68CxYPD4Fzsszg6d3YjZKkf8
DhFYpZLrThOy3hhSfWYDLLspx8J8lBGCeNRv+j/tcHDe8A6SdyhSbHTLawlX6xtd
PzYWXVTnvPO673j+ObQttmEfF9KXiTTyqDkLboA5HD+7lU77bdHIHBK2+1BSiYK7
HKm/werCgOFud9L+gL7l2BmA2RHiTX9JU+Z6aHzorXgXF65PKqvhauj+xJRqqOCX
mNmn3Sg28+8ELveE/ltVzfrWQA7TgeCeCYNAO6DY4FR/y14mEd3Yav/VXQGMIOR2
/2Erkz+2JhCOeD1GtNKv/Gdo0WyDnEQVz4VqEs0K3UnwBK4SU8F6SSNkDVD9xb5G
zYSU3e1xf8zeEjrrcGZG2dpZTqqlN6wKwdWT9LIgQ4corIXV/3s0Vnp+uxE4Mkzp
wZ59r5BNib1UV/vmWfiVZ80mUVEoe4ASkZrvC6RdYcHd2RBPVUjrEXv4YKkhK5b+
FdHu0tJKVLHoYf7YlSlhuYI+rXb9uXl31el5nOibWonzoMi6mQlulruaMMy2TIZp
35+ILl+oY4SHNmpIsJ3derosPbI1kMvOOLsYAc4YPbxqfw1hB5FqH7dnPzNSPiAa
eeh+6P0KbcIqi8cdwx6DPP4TwQKhG//r4Khr3iG+KDo8+CD3NZntz75AsqlMNqLO
u4AvP9u8wESK2VVsyH3wsf6SJBCmUeZmopKKcpGVoKXavYPMOTVSLSvcn0jkAVO4
t80EJ7kgHXRXIDwVuP8pqiSKtlOjnEWo9QDe96jvfs338IBTfnEt2Pj8es3zOhub
ARR6Ecz7PEgb3CJsfjo6nRzkaWFW3QREdEl040F/jf8nw6uJH9dq7VZLXwe2fN4M
qhf9e2RrqVtMk+0lXJK704g6ebOeAXs+JTMTKPPdA+ZkJD7gK4lSVKf/6fE10SFg
PCb5ahd885iTrPHBWsQWVNaqdiRUlp69qCaMcXTVOgAIQLUCehzZLCi1YE2io3pe
yGhGztedOx3IumWIupquYY6HwjqTiDny3EeugCnonIKK8buCbAF7g6lH8cb6keP7
sYJxxG0U3/imKDVZ+UEKqgj5DSEdO/MvCIUfIZW4qFsd8WLP/Uu4TJB7pP3PralT
98pkdtWH9S/UtFMODqGdlxrpk8BUhI8iot12F80xYKu/LFf3Z+op4opxoemWtPVT
Vw1bA5VzpzhtvQJDtATH0R5JKWdahNN1IA0/LVItzgjPKByiBuTcdULgLVp2TEQ9
K9hivlEBtzGsp2J0Frdz2hdIdZTPiBgMToGaBgoPSTvkrG7ZGOcWaTtVrIXX+lEP
Ck5jYSrd975Yb0XN8NSWJuGDBgKtKYUb25HK1a5W39pR0IpfCImqMuvyAAHiGeYy
wa3Yo3QTxog+JcBIuqxbVs8lYz4wwcoOE46uDTfRD7UOcwt+fjH7Lu9lPQIfCdEO
3N+/6IBl39G6GnwwQTIP1fhAA7m+WAdrL2Aa98+qKU3OAa6e0mLOS2NMD7q8X41k
R9qku6zbXbQ3uIAfPVzhBBpBJ5LVN2qE0bdgykV2nKlFLvZUk53n70Vr7+i6GwWC
8WcrW61h+hJHmYx9atGYVWIMWyBwlILCPkyAYxdS+TdRjKaZuuO2r0GyXq+Trmsb
oxFE/Vv2vXUO3DLpR2IIiLqCelsem3sDvIHMfCffX4XZVzCeq7oy5MTBKUKVIvXO
CbFE5496wz82t94qC6t2NbVHyKva+oBy8Fq0Q9Zocgwxpakwyhzd0fzE7PaWOFl3
WZ7h7mQYIfeyRKGFZGgokWjRLyMBYisdccj3yORuOFzRumqJ296rwBgp+I2gapKy
nGAhhcolGq4TkY44mRy7T61j+YW3aDNYLsrzpUBLEgSLTmkYJ0IHlA1K/+dSKhnI
Zpp0jIgz3nMIEcXoa89GwKfQF4EbSFYvwmKpJYsDYaXbiYwjL0sv45aBeNMzIHV7
EcFde+IfdgabMsJi4GfvGc6IWovw4SOgZvyDoNwKA7+PnOO8OAmP/avH3lohPXLD
NZaZ6TcNrjFG4osfKX1ANVCo42+vQzqL4LiXuQtBeFv+Jr85VYMxspH/gjmHTASt
uu3nJnX+rSeGSMlM7kSXmVDRCF+wMRgoiTionwm1F14Ze5Mfoy+lY+4JXI2dhNz4
IiPooYLHCWjWGnAdceRR5UGU2rGquAF0ukCFboqWlXis8F/uMDxxEmgSZxUGLg2S
1ei3eBCAAXGGUKCxJDMEn9WSVyJPVtuoddWOsOfKdCpJI2mUo27D45oJlgOsE/zD
2T9qZXQh+fGF0s/ye6IRT0WvfME5N8jaUjUsmvmLLQiPznzXF5kqbb4zl3DkgG80
VfaqZpyurlGw0vBtnmpxe+R7YT+mIj3ZDhI4+RMCfl5WQp9Mmuy91Pjj9jG0c9BK
61JU7XJPkUaZEqJQVRNomQESeoUs9HChlIObnxt9RYiS2Lh8POsFFIVjrQIXBzqe
K4Nqavpj1IPW8j5la3CZaNIYePwxYmMx40U8dAiyOEVYn0HE9p1uHQddC96QK9zS
OI+hy0cKY+46UB/5gTU6MADuFlkOuz/QbMyUgWGMABfVswEnt1YO8mExrViwOJc+
7tTWMpwPDxkNViKpgPxikFlvL9aOED4xKaB+A3j4Q/oiedrT0I3+xvkOMBbXF1FF
rPzb8fdEKv432N8NlRoRDHh2dSFrpqxLqKFUS65h9DinRKiuC6wq7+f86Wg9hodP
PX/H8l6EFUghVNEMi1nGNrofXhw1qL+EBJOw4L9ftJqDaIOk/u2aLjiBqQSYGqHD
Qv/hqurLtVDXTRK3Do974mXvP8hZmJk4b0jv1P9p/OAMqhVM2mNVrjB8bNUIUBZD
tx2ddLtx9zFw/tmxvJge7oKGgBPmQVYjSeuSDdiikzEnCVNMJYDCHfTyMvFVX/QL
/C+nCugYGZwr4Qdo/28K2lYRKWb81HXID2Eq+teG5gHI3PrsEhEHe7bb/wM2SG2v
imk8SF/vGP44m7RXh879U3Zw2AkW4TfpduY1YAkYS3Yr/RQBO0yOhcLSzzFGmjwG
Nu2oXvwfsMXyz5/tf+VlyyLq28fpyeMEdOJgxWM7UNhtH+qdBb0+P8LoQpcyrA0F
twHlh6Xe3HJw2seY0OCDcLeLm3jsretyiPozmy3UP4VA45ps/fIPkYLFvJC6XgSD
nsBCk7yFI6HqSrx1+YF2vQcKvkqUJNo80Ws04eca5aq6H2Aj0YC7KqQWzJcsCLcy
4O3nkYzghI8tEaFOYFReiw==
`pragma protect end_protected
