`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WQNR0RYcfse/7qSoPFEQ2QZeMu9Sa27+0sDDAuTdB2kbngteFkXRMjedca4c2RLQ
F5WqXA9U6+UUykwuAU7BNBBTryQnkqhdx/YlmtVDTx5ddxpzpba1MkCrxoxfoPUo
PZ65DRErUumdz0VtEi9mXxrGVroPflpbiioiMN23NJE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21984)
O6CSqJt8RQVQw5v00o4sEphh15SatYwmCUhPDsURUp+iuZ8dj5FrUdFf/lU44q8c
i5G0O31+2NTimiw9wahR8QUqaaIA3vSZ+eUYSeyggZmIWMP9411X8qwGsTePMpin
5ujDH1bZJpyRi1QxYbxfIGWpdOsTXbsdghSeo2KTc8c2eKNcSuVLBedg+LZInQcE
U+UurNaahPdJlJYBMe69ZLtjQXSkqv0BBifIwsO3nELlklC4FcIIwxrhdU7P728+
HkXrFMeWaAUfGwvktkfN2mmbpE42uIH6FxUMCzTX5EAMNKtGB6cJ5ShcUK26UcvZ
9UyzRFnUidAGuo1OY83fW4+slhxxfFhbi3hGQa0bNizewKe9wKmvrLV9ziRIgFxy
s6cPudVrETgoCM7FBPOP7wDshyvdXZsywL8PQtjaEYtJ8ztFfi7w6YDp9P+cxKM+
gm5tn8cvXlSR9Gn+0BbFYOSUJk5Ef+IkU1mjgmYMuTW9HZcDkA/4qNW8aUPYVZoI
wOD5N1SI7Vet21+GXgxUUyNZUSP8OeFHbtDMYjg45ryakj+Knp8+6020ZZO1oV77
dTuXb0c7HidxIF0RfenxNMRbPZyB0Lt7CWGJa6Ds5kgHMEyISB8wNqfnHmMlLsdS
j3Cd7uFwLyF4LsDT+sqb/0x+PIbHSw5jAYci6HJGt4e/iKT3ExhnQmkxix063gnY
4IAfzemKNi+jjx92gSxWE9fa+lADybZiya0p+WNR+3mXND1gZmFePpBub7Yd37s7
NOPoj3Ba1g+ZdQBiteSpUAiTdDO0ryUw9+/U9ZiZw6JnK76ZrW1zDYgTPdty4HXO
75BOHn8asIRDxlPoggzXjLuDyHd512J4q/IEnulDpj2EelEhQn1TCQlQtrfplJul
hy1oNO5M52fkXHN+iL7euEuCxIG93sG2jjl0SqErVQ2TnFktmEVgCT/ZOit2Jjho
AptAxpZ29GyQpseQdPrgpao+8o563M7gSx9/W4ciCaKOklKZ6nAgfxPEYRGMt04L
DOjnTYaGLtahdCGJAQQ0zdD7kPsxPkYzJxRE0GZ7vX7iRWWXYOPf2g1PJ4IqGAuM
J2a+kHppQrYSAh8VRBkgyg2RCghkfiFs3glUWKB5BRIwYWR2legaJvEgS8pT4+S5
43To4t/rHOMq8dS2m5aHacJzfqjiXT/6Z0tvIbBWDLKHlMh4SUSw4OFAcvJvuO5Q
koaeBD3o4C7mb4NKZXl3tYjNzc/lWzNjYXm+PFUOm9cEa3ZFQK/z8EGrrxOzsYAE
Qd/cZmTAJ1F6MvlfLRykkK3afJg9JXlE2YVe99YKiI3OyuyjXMJgVDyhGKDu53ap
7fh2gn1SfJXFlgf1IbW03U6WL6JUl3vcsU+N8h44IWpMvFynUgtSL9yVv7OJ43b6
fzeBEsnZG7Mg/a2ZTRyVEbW71RCrVGGoaFBZAT8rE4gWNhGA8CpXj1tsobLkRbfM
LrifhZR0XDJX+JNyqMMMoDSa0eRvCb7unTKOXuuuaPR+1ZrlDBKIhtPMuMCMNjn4
pcqQmN2ANGt+S0qUYXdRJbtsLNrf87fR5d+qE7q77Rqf2YXJE2xzxHqRVhZ3ZtZ6
AYc3NCKvOyu85Ph7AJthKOr+OByPDherrCq2Xsi/vOHeYhzaWNs/ecPPlP5QA/HX
t1aU4Iy+WtwIxLbEHCSZzsPoHUvP3PyqDTsDWnrolvVH6KcmreMVUwLrd1T363d5
XPN6HU1NSnrCemP5ZDHskAVsfA/XEkOSe/G9f9PwC2ajuNVCm7kXQrKW+EBU9Mcw
BhFFXf5222kptiBZ8EQ84JFiniPc4JcWsdQmVfkEi3TX67F5SOyF7PXyWrdvh0Er
zGVFUOF+R7qAUQZ2qd9wA00Kq79QU31BZJohiiSsI0GVVEM/IgIsMyXPXveicPEF
LnXVjME+/Lq/1BnRU3ZL45pyDbW2TE2N+pjOG3Sw53gxQ+x1qfvtfuNYnlJMSs0r
WGj+9PnLE4WItXgcpW8CeBvqEJWkAA3NYSMCTDq5A/ld1lhVGDVDAjCi5pTAuQ6o
c5Dxl6OIB1jKs+XZVOE6iXAMz/B7sQ0dX9n/tjfMuqLTtk7kn95Nks4Ahu0VgQSG
nH2k6qkMt3zTmDuzk+Vx1BWv0u+LMI9NMrKGsikcyL+oG6AxAB3xk+IyjcXxUqoo
uO69J+Q3kHBeSEfcBoXqWa/BZp3wGdwMISuqhgFmK1L/M0f7ZbaT3to+miRwAqBI
+kZ6wFizQcojkpx7Xv5vj4JxUIS4UOUgvOo4tFswVJkRXnWTbIrOUr/0nRYaxjf/
iTKpAU/9wF1B0LgbMmRbpu9i9Co8BFWUNHoPI/1I0C4XT3TyZQq1u3n7MEuz9570
4HA8z3rkAbt1flU6uueFQT9+9dL004YzDcAhxMLIwtJWG5kZ4Spnr14vewhDEedb
at93ux8EgPo3kkIL2Okt7SdocCQXSNKs9wM6vf+2+xhemotVYcACKkK3G0DSj11X
qY4Li42W9O/CFSq/7PCTDPNbp/FQiY90GaG+8zC3lXIfrjoW35iBhCQ1dyB4P9pY
SxRXRqkNRPk3ahDH7Cb4vAc2kYcwT3gRzDz/yYkrlQ/FRD7ICHt3zZ+dIO535N6z
sKmR8vtJRtsZYrVfRF+VoysmCd8FO9J1X/APwV6+M/pfOU9Bj9/umDKOtMslc9Ms
ZphZOi2uvVrOGaxAAPiMuzu97DR7eS7m+UwudyygDeOjb5+4C35w9VDPQu+jmpo+
rMCu87DuxdsHe3M8ga5be0FEpY2c8E4LU6b/jg2Gmu3OWchCSDgiKZAb/IvPRHCj
kghfZv+ncNitG7qUOtf420riQMeXUCI8lTW1SvQ08rU7EhDHk7xDMWEiubHVJj8q
DudqXdUN7N4HauGByjjZMYD8gRI4QwYFT7AmGwNcK4g0ChAR0vkJn+KrIUYZQbMD
mJvFGY4l6Fz7xuKxPMMgQJejTaX5qhBKfJKogvBROdRSB5576YTkKAYWDvojzcbv
ioBqTjHtJ7xd3i/+mzk8HziRPZd9/VW4jLCi/MlnaJRAvq61SlxU9aJLKndv8Npa
BvFuhu68D6RynlcEINzBzOrIMrnOWRldovBy8CTib+b1njyLSOSlLaBx1kAc7Rls
1kynEhtJ3MEBQhdmQxB0MirooUrZ4ycBShSSnTjX++A5lBirxYzAQeYPdYQd4rQG
OeQd33+TYCpOqTP9afJ6sPIAzlmFwjYIOXy2WW18mn3dDm0YFQ9Nn2TtfkLSNHJ5
zOWJ5Qb6/+FUGTasSpLMOWHo1oHNrKHIlsHVpDeg8VnIklF0c+iU4wkAaba14u85
x4gKjb9idrvDgMX+myjFJpPOEE8P4DTAAlUp4ALh31bBTprOSUJTyi3KAqiBeoZd
q/+wuVr+hUvCrCYdGYLQSf7CXpuWXJMj693OfG0jqQA4Oh6p+Me1VMFB0O/Ur526
ROJV4p2UlITvG9jTfD/OM6/2BLQ1e3nAPq3RKv1vp7OzX4I0sHnzjia28Rih8Qo1
YXrR6gihbjDnGZusCL2KmWgOKoCdPRuj24LnTLkWflitwxeA6phH86uNSnwN5TSb
aTSkdpyNBuiG+Q24e5oWIBXX1HVboJW2D3gTtasYce38h2kqmkxTKTkG3dzTMuNN
PI1JbuvPVhG5GJnK3b3UkPbOxWZfZN0rE6M5022rMfzw9k2SFwxRCjW7+20vZbVB
Z4vmY9AB4jTNOJoWW2KhmizfTLflLGTvdWkPepdPGl9+ueMnDYyr5QqyFZ/Hx1oT
rbx7SrmNlngUbrIfqI5pNqgqGAxsjVki8c0Qa6MRFh3W5ZqW2kAeatedbNHmqtQk
vfTiiTjeMAWza8DJUGxLAGiR3Vl429WPws6nH4wk4fQHw3VjvW0cHvrZk0Y4IX/P
TID7GWf7850T5xfI9adHzObq/g2lfGivjxDqK08EAsfJQZjQfMP5UDm7rdsV/flL
fOxTHKyjEYqrt2aCKu1bkS/rQJNPcvQcc44IEarSuNAS40nwAtE2i1+k5f6Jx8mZ
ykq6ZkukrSoefHUxf7L/utE/6oiurktHJbLCVFQ1E4l7F028N5/anBlFDYyV/9Q7
mYgTGaGFcU8GCAU0XVQ98V2iuGF0aTK8HErxdO4eg44fEgxWoXKHbCVzfwXfRi9A
Rk8YozBK+Oz5NpyTGlS+4rlRHWwqxEuMrQ9pmlc12OeZ7Us07+N5qdKU8E5Htpy3
3RTyZv5GTIEbpMckIbDikn3v6xrISNPo49xNRlomAucNo9F38N4YOBnA6ojNocup
3cbMjr8yAgx1o2Rp/mILNhp7dAaAUqK2a7As1zf9X3z75/OlKauG6klBNIMGm2Ge
D408eR1FKR+iG3TDR451xZenziETraqDuJF1gtLfIDS3QcKidBr7QNs50GzGzZa1
yuWLTp9wMtFmFoXUXWyMqwJb9bhBFXLQSwduSmuAzhBWDg1FW3r2dPkKypcGiGyz
VncE2O6BQaGqefmXFCOotr5EQmrINVrS29PrhTbAAgPY+Z6eKCslkxgKdXlOJatj
ExBVNqtX3NaBvlXuyyIR8cbFsgaBxJ2wu9vYlvMgdIFFER8EMMULxz207BvDD1WO
dwSfLXDc6NiXM3q6LBrU8F366G1OIZXqvbP0seAxXlZ9Nu8R5UXPo/CyYCxHKu5s
XI6AWpxD0N1ot73j566CCITWxS+xMHnAxZrZ2qlaVwAQ5dj5fif+Y/K8SWStcw7y
FJCqWlphGwgGcfJ2TGihWSRUnV6aXYvQBtZNtitvCBJUD4g3+r9FQ58GiSm3JHKc
vDzvq6f3hgjXJQiG9g8XFWpZZjkl+Di7pOjuePC16AQIRq4nCyP5dTFM1ehhVVfe
MOaPfCbs6mCuBR3Sdz3Su94Vjy+4hpEHBd+qOsG/uTWjUdEOUbq2A30/UVYg8EL/
ACQSeeQ7q+SdLhl+TNz++uHaDBANM7nlteUcv2TimQpA6VuM4S/3rh98+zdTOf9R
qBZi2UILunZO/Q/FpazhWDaKMeKi1jmNs7Rpx4yDMavy+BmkHlJ63Ag1w+bpqWcL
j56fDeJKFtd+/Ue49/PAbRyVOPa7b8K7VHahXQlAFo2Df9LhKsQZEpOVD6nHrkbk
YkcyeIWOOg0SKrC11mVeea666QehqNQfBZgF+0kuYV0LUO36uOmv9y53nOERiQYx
mW0TvjUafjTomkarSEOzhJo9Rk7NSiM3qga81SuJgVCRsCEuOelvxiBfdq5xyxA1
IjAYBKrtMvVGYtuEKMQtPnO8uO8FIhqltT5zx/xB7R1L0wEovpWP9PgSQEYsR0AI
cOpClymtYjUU6G6rZTn34ZryStxFphuUP27OsYU1ao7pfMUOVbfsWuSw7aJ+j8H2
7zPQCTkuKHUfHByKzHguSFlkhhRQa7mvsq+6NU4XEYm5S3zctC5LECZT7oEvfbgp
0XpQTKnjmIBVUDvutKuCMluopX4x+dPwsKs69L4S04JInphoi8KimUlhK/DxkkH7
+IivRe9yi1oPgFNMlfuvZy7CQOo3zgr4ZWPfU5AOLDKs5X21QdHeVMb6fcPEnWsP
406ZPX2myky99o+YWUTo71MxJhCWoiHJxOWk8taHLoz/DDQxPsxcDxsAOTEus4aH
W2kaPDrIPM3UnMLDpEssBNEM4aYkurzUMk+swTFqfSSVmoOTtyA/uPhdcn+1M6Kb
9DROFmvOqKchrNmncqd8Hemdu/pbNxEW9Pz3mWvYJpJKLwZtfeC5KgDdS0H3RMtt
G9pSNcuJGw32erXif/UsSdhPtJ97aQ80qvDPgzk6pGxlAmm9MLmfzHWNiMDB3Dcz
L/mVTxsxq71yGkAx0JxSzlGyTlPqs1aV44/9AY7mED1oyQhLBhVf7cNVoe6cQjpU
KuHwpoGVfA2RHSMmCK/tPsObKkScYIUGyLeVTS5mwC7UCN0udkIzKGmAMZtY6GGP
FlIC12MQnXL2Czw4AsgM5Gn0xVyLevLJm/AIYrYCjdEI8zrquvFZWbGd4gZms9SR
9vn+HSj5LBuS4zF1zDBhBK6b+8lGVeBf8Rm6Oth/xugllBNJ2ImiZsvvVzz8KWj8
yPBfHmvdc1kDP0hN+pe63lZ7yQTluux9lTchXg4Z0QczxmkN6zzzEidQM0xa7SOl
hSN+hYSIOgWLtOtDCPnezMBUBxbP6arN3D1CXHFpzfBtIhgZ0E5dLv3/vPLZgWhr
Helc/d6jnE66FWNJWvnVODq0Fe78SxY2VkKtJi3AZ5GvZij0v9a/ei1/g2769OiZ
NAWNoQOBi+NMXcJd0L+ON9tiMDVZh9ooFQVqPTs917knqeItAZUHCHEXjDJ5pACi
wMdZRI6GlkZY0H7j0SFQt7HIJb2jjlE1bPTkjmZG9frX/vUJDtVTJy+cK6bCZUEK
7IvD3M1wBYMRaHEU4Wlcg8M/3TDDaDaP4lc3ZvThjo/tFBVm9NhsfHKyuKz6BPmi
otxywlVlXgG8Gpxuq84Q0NAmhbPenlX7PfTrapvmRWl0cv6LHnjpzNi8138v8dr5
LAbR06bqFzUOGCE06+RY6FHyMM5USRYlWinuaNjSNldVI6KQnra0FlotSmYcNKgP
1Y9bKIJBgQJBRVIQ7VtVeN2OKAyCMdqS4FZbxEzTiB67j3PDk0CuY2FkHjnr0Wdh
PN028o5Lki4mRfw3h8HGuX4H6J8XTYKdlnM8sQKGZKDuxVu7JCV2vu2+5cN1eZWr
hprwB5zeJX34m4se5MlyHLg/65Lteghv3+tvrkwTRPJhZORGEWCAV99UwctClbOl
5bhsuYfNe+a3O1gR3UnZB0vdqDYawO0imRLcFIhdpwuk6NgCr3VXhzxjSGcFukP9
aMRQU1WN3iEY4TpzAj+Wwerp8wN4uln3R6Hc59n/mw7QE1IJqOuxYoT0DD7evzCl
iOiW+fcD1VBz6tuhJ4utym3YOBafHNvaNM/IG1kOoQaxhmdEgPkXskLAS2pzXAdD
dZGgqEWxtz838ULjl1hjOkxdsXNWMNwoVbb1QRLkq9OYAkAo05jcV57nPc5b+bhs
LH7Rclt66xBP+1I2tT4nBhkcp9rUTX5waRGRBKq/SwfxtIDJZuFmg1e2gE5ZQgVf
SqUVvQ46J7/u53kVlir0n/0b9OJKbVVmHdPXD6aR6u458UtcJtNH+GGZ2Ln+yGM2
osrbt/rUa3ScEoXd791zo2G5iYOxGWzusVhSdKelaxzDqkBm8Gcw92EkSWbnWk7m
0Syk6jgS2m8jAs2e2weZnhodFd3LY4XC/CXKpTCXR/bYKKp8vFTTw+X1hM47aK7e
KUsODIg2TKxxKwpYXI759q+aUrk+68KKTkyDkAAHhCKJbmX0+s+ly5BZktkMENly
1OKkYGfx9Ai1mX4Cfa1t3Y/1I8DlDPBo0LCLWtoo2MDa6l86HNkyozMUjln1pEjX
YxHpozFY8A+/w7Gp++3EznPvOrGA3lvlNTYyf0+RcsLrCN9vqE3/eoqNeGHQ5Jn0
yLWQuHxFGpLziDyc8hQU0q1WvmxM6PA9zBiz3/nlEGR+3sEPY4SpmNBzxW3QAm45
ZkfdcgntJuG8afFFvG4zObZwcakk8agNqgrqnK1VWzu1NlC2zRHkYjdUAE9mxKg/
xgMhjYDauzqe2+R8QsQMG9a3hvvqmDCX1Gsmf6AmItEXIsX7akD9ncA4kL9Z+srX
d7YPSSYDJXe35vJmjnFVj/802ZusuPnvVzI3+PwNS0iu2gyDAhtNWY5CW7MRvetf
8ypia5ruj4dVTGEIFJWRX6iDEXRyHpz3b/it3FFmzXJdiz6F7dQZX97fuQ/Hm0oT
MYn+AU2qpzu19w8f4KM3ABEVFCorTgL1fUVp15DL7UBHHlkB2H1PEfgG2wNiPQUZ
MAGMhg+COX9HbUAErO8+IzO3PJEuXI0rh8KAP8Q5aWdilqO2Cl90/rYUjVq3dn9U
Gtucm+wYoKzLvYX6LMhXnK7ECySRf7H2yePdKk3uKGgL//eU4Z5AiMKW2WT4TB8j
83vWkrTsYaVF5tV+1FNnwV2YRdYPgsMj7mwMnxEpHPAY4luprgk8pds7e4LLS0fV
sSZZXJ0HvAXZaCpOkymNnFt/JPCXXaj8bOHlqQPC2KFrf/FBpGIIuwmA1NhRW53I
cHq6JMy7ga0KiyCruvVvO0I1VZ473swp5I/ayndIb4/Hlr6Yq86GaYcOZ45RkNYp
MTMAKd2BufYFIFauBmyo11FToJFPj8gXY4ZrZ1T9cGH4pjQxR5jOJbez/09s1uj4
wtchVxnpYQfBIk87tj7AGetEjs3RX5m8tSfBWvSni1qRrrCKBCKKKGZSxwQsw1ur
sKrIC10YAm3DW3gOJBbVQHQX/2PIXBtEcbOoSoOt0lenzxyxEi9CwjT/P+r6bVK/
fvfQBzbs0JazGso6sweG1003je7v13XR3NwD2P/hcQLFsxvWgXkbpaN8m3uedQcg
jEBPbtiR1fA3Kry2bIfHhA/q/4YW6OMQwPbbnb8oKZmCuVjfqxen3c+DpEY36ODd
DhxNcn+U+LB5gZUEB6D9o8XrhGWy7NK61IkLns3JrZXjafZ2aFEOUFZBjsqdw62P
uF+56AUwWVbOD+PbrWKwmL5vFjmhKg4ss9yYwzLLbpsp+v/jnkZkVHCR3Bpv/buE
n9UqNwsnLeCE2h75DtnjNlCK2uWpGqpUjSuhUO5IPRtURlTbO9Z/PYXgN2en8cP4
BTpIVA2WmZ4Fhm+ydlHAI1+BSpkG84oYjmE+qzRFVj/s1X4bKS6W8nHyHbDn+30Z
2m+rDYadQwLgao6cTSo4kPmBSeFuNb+yM3D+irso5Ag87NTR+wk5Fr00ez1gr8gU
WLi0n7YCoexoSbeOu9kVXI1n/acvbLgPk/p/tcbEaaPeLGZRLfFF2niwqnIwzlRX
U6+qPKIwQ9EtGy7BzOB2kVXm2MCiOAB3V+B1QcXcfdy8toah8swDEgKrcTxTDZqA
ViECwd2Q/Ub1YLY1taODh6YhIgL7cdHHMQXIYHQwHEe7fsrlOFagIvZQuiiDSFAj
Du/HHwQc694k+ITYdG39NF8w8ZGgGcSvJxO9FXH7vPi5XyMaraGq6/M1wTqR6ZNa
jSMWelaq130ed5LH3heSzIksKMr+rjxPjKnMcjr4sJjCzsJj8X4WikNRuBy/yAOn
UI4S+0Yb4GJRw6lrwDWtfStrK1Rvmi3b9HVK04UaX//OmpwBKIG/FYRyuWAftD8l
zFKliLoABzTuRl0e4XRaxXTFY5DzV5C/2i8e8h/Jy82hKkOnp2ponlr7Vjq2tqIu
I4e3jxIQ8qmKRgI8ufTzxLJFD5wXcBZLBCsEtGal5IBEXTlrTNDs+SRsEJVHm95R
T51Gdm+aQL2aSqbP7ae8a7ABpbD+fap6kzAEz5CwKumISIiiEkHhmxc3F/U0We6n
RoONAV6kLQYVhzs88ogAQBEIr6ss1fstSKjip0VtDtP91kcxrS1jmw9+s9fY8BMR
/ut0nIvHOhlxsapv7RejrKzakRBmq4YUbwU0OhHSxatQit4IBF+wpAtmynnoTw+k
wDDnre3qMf/MQl7rKOgpykABB2aD2SqdfLQt5qPFOF4yjiP164Ep4WLGM2xhWe74
I7IW060sxh1ojX2PrlPz+QbIfFXIUx5MRXxQunMuLbFlZq8+7S/FM/4gy6HuSK1m
oy32pn9diRozNYJAXTNeqtbUczjzHJtpuHQwGUmxdZi/OjiCyu1fQv9RUBRpIkbh
xBQZoYUI7xavVt0Z+7ZY6ZidFNB0K2Bzs6KBoIcvt/9Yk9LhMF7+aZea9xq+bm7E
JfTGI1mKXOb1kWANSX/F3h1eZ0hnpHWZHNiHiuZJRkwB4+viA+nSjI7P3m8po2/1
ZVaoO9XtlIk9FrKBmaRzZv3w2RjlO53Z1+9oobtsxyW9f8vWfKySO9nITmwL6625
+LVFQRtbMJnQN9ybzTdUR2tJdspjbfwQ7K1AmqwLnUPq7/TAkDQYjURyO+G6z3FA
RAWv+t/vM1HGKHf0J5mHXjgDx2xjkDWkEUsv6588vx3qmLYBLgo7BZCKxxP6rFEg
Ky3s6UXH9kMRXkweH4wNrJwxqiDyT7j3+34OQAI2GftAKGrpRH6q8eE5P6mzlxFf
Xi5OUy5ce7wqEsp62o+c7MxvxoHKI49/JTlKwfUEHBDq64qaIKjkW65n7ASd0vWD
61T21f0mW6qMNMrZqYNJd5DqfrXpNDeuPgOyAqUFHP0mVzcjMPhMuER6Ge9tjcnU
2bznhUvg2zv20ihqVwiDi3z5SESL+XWGUqPDeTmFBZpeajTdjG25Ac0aLJew/H3v
6RQ0B61QzF1F9MHdkcprpTyY3iHUcOXfOhoIsJl28U/D6y0Fu0eP1kGdRsmAPJnR
wMcsiLywFvVEjmPVzKIHsRE/KEExFETG5FZQrppbZJhTgWSAgI9sIW/zKZlHj1ca
F+0GXi/TMzt8+/DuxWD/owa3Sjcr3vkZQb9llGeF3KGddEuIOjdrIWY2V+eLG6kX
5UlNQw0MLMCrRhBVzw/LCq5PAseQjeODcep60nXKwMgrgqbYvHlUUQksP5LgGIWN
5l1Mh7NWlH2gikS+4itNj+hnMKx2+eAU2vx4PoufJdqtQA2MhE0hjjkRtbh+9pyb
w17OJ00e3CXHvhTHrLsNrKOy6xZSmmUKW+LLZgz74zV6QxRIg6xXRZ2IthljuRJd
JG+sEDHzWrOrAMyYI342pnGYPjC78YBOWBxV8g5j92Xy9vexCDbNVPRo5wejOVNJ
1ws6Ugvczi5hxeWPOK1HikhA3FuFTW2mcAuQnZu+emGFD3eYhNYkqLqT8/eFAIlF
AnFfEAqh9IwEbZ1TrmVCh5NF50z+hwPTFZkk9jWK8CecQQpp8y7NsOqoiVg0KISF
KEJA992dlc1N84yc5klgIHbsd2HP1k28+XGlWEamp3O1A5Q5uYU+Hr6MAoQ+WaD0
+878LrQpZPJ9/kFhK9/e7CEqq82W24WpbmuTWW1VWno8lxa+TWp9c1TI585M1/l1
l6nePkP2Q9M+2SZ3ZNBaRTg6cm+iRjPtdJx8403Xva/uUAz8OMeC7zmnb2BZ7Dx7
NaSnlvP79A+GnmIwaZzyd4RsxgmRvRHex4KCSUfLZsN777KGUCpS3CNnF6AAOkDl
aLK/n9M2XJdvb8Tl/eDQLpVg8G16vGz1J8VddIdWI62Jp/5z2NXCYsbJpfzcaWPV
9SbuN14aSIsX2ksqjGjp1PwBoVM8Dmsy4+5nGTR/OENJs92ZlPaUwOsa9gNuYLT4
rHlX3c1Tq1nqzPyIzAn9p9bMkOZ1aUp6hN4KHISSGaiZwQXXCQQ8e2/xAYLcAXyT
ck9T7h4149eBH7r9h5k2OtX8Olfb0WZLh6+3faHJdLFrn9OLjxxwI/ZWWePoiVBg
PWETCczMy3ekmxr2Zlr/ZbuNzE59OIZghptgsu0C93gCdd9f7Bapb6Wuq0g823W7
f9sbPOZGSafy+z6SyO4Hd5JC2+4X0og5DBHxVSMlKA+lLbu71DdI6jTNQrlwBvQf
djdQIfsdX6D6pkfSo1ez2JyL40YjGm83gtRXlztOggzRrg84Cjm+5xzc06H80/zm
FTsTLeoi7HHr0oIBmjAXJBW3yL583TLXjB2oa8cd6iQMY7ACXLMAuq79Ac3jZy+C
u3VTjKqE+naHGQxV3tpvfF5wPYZbfj3vmJjB2r2NHlNhzRc4Fwk9wAnKfzlU59iX
ZdEoVr/LZANB+/uCU/fooOkRFv+Gq8HnIDTb8kBfdSryoX+3bDgAdtdivf8+3/tJ
VmkIoakVafb7zmxchmPasssJXpmQ5KYPbcCv/g/TwJWzgvuiVPa0MTIcTBV/zP0Y
vHP6uhnGe+zjx/MOVVYO+IFJ8x59/e8o/qev70SS2ZDh+b+8CMLBQlDEKkw1vVJO
AN/9I7XQf/kekdm2LUnjK78CSPXa/60NX6wQs7IBYBbAlXdKaGymD6/sYzESWR4h
fOR7TajVCq3aiC/CTr6pl2BOP8jLvEawBZ4oLiQkF9rdYbp1d3mWq0v/Kg/e7pNH
oWKF3cJWr263FUjMJfB7l5Cf+lhTW3ty7Qc4vSrjCRH1zW4zBLWfI1/S9tAnr0Es
WSnERpWC+SOfeaijv3XTDL110MFE2ZZ2Rbo5xYtoIRgQoRCe/IdBNU11ZXpZYpNB
KLuop0CiYK/HgRN+y19rUqY5PTRDuoQMDFUGRboNY2WP/UjRV/4LubXvAQYnRoWe
hYzug2BqYLNdbtyE6U7wK5OLDN+Ut/GEyoel2rWSc681BzWigVQ0mNjxcb9X9ZAW
CrMmuzNbwQ3p4azdfNPuZ7AmYz3XpYvgcjOXabUJ5XgXX0RmZcLZP7GcdV4BlE+c
rcEVnwUWW9SGRHspjTLdFKRlEJbAr5qVwsmRSThi5Es0FTJJTc5knfNRfJGdiOXC
DXJM+s3GqoiOnKjTNuGSiSW1ygPDSwDtlouKIwneCvvHejlqKp0HvEuzS6L/O98B
BIvhkD8sBZEZp4GIhdYVJl4OqxlIcqMbvm9+4zzO863cFU8dwhMTq1qGtutB00KK
CxV3CfW7MJ4W4gX+BTy3zzaDhhWkhvxOn2uKoTconaA6BDOpKFernb9+fvrHilUu
EXTQvKwTYJsV7YivRJQ/QtZyGGGdmJMLZ/Wp7LKZ0zVsP999dkVvGXgwlbmJNtIQ
0S//WKXGBCbQBLtWaobgt60gbm5tb6CLKWMnMmRnUF5Be19KzlStChq2qSl0IuR0
h0dUN3W+TyVY3b82bJ0ntaW2NREwnbTONB1NWcmqZrr7zg+RfCq4yUi/acyKBM35
uKDKGJZT9ZkOSd3OlaCRgMbuM45WqcRv6e/O8SpzgiJQEHAslfbOc+4WHs/LpPcA
9cu5uRUa1DPEDa6SC7KkR2ET0S3XZSl76fME/X1bguuEj10maxsqFgs+PQ+8kp4Q
i0qS3EDl1bDehCH2rrrm6c3NjFjTD4m85rr/F2Eln1W85T8H/MXom3VdMEbgIDPy
L6dW6XYrQ1EBrikbYmggpwGvV7sceF9sNTZ7e11zah95cLxNuejtn2RzCg+IvNTw
nbQlVoe3CV1UE4hYePZNfI0L3aVrmiyhvrmJsoBbbvg7QWz2F3Zs97zfX30R6vEd
oik/7EjH4mrCVr2VQXA0V4DILso8HUz8CCEMDm2LgIwRjaANeD70PwQUuTWPyTEa
GoNbe70mbQ1H7DLpaJE9e4rFjoGtX29En+kAJJXsORKrISCzm2EFhvpfMc+fD7AX
00bSj5OgHbZwg4g4ECoPUPcwlWLhwivMS6N2V3J1nccztFGM+smsh6GRm1nWTHMJ
MjKPNHwHzF9x6HNmrgpoTT49PGiLXIcvU6oHUmfy4skGQSigRO2pzf9ZxuDm6AFh
vNRXhuCAssa5gR4C/jyWimN3B4j5Ems0/FFLpLhgUS2sdKqmULNWNPpovq1gDFuM
HaE7o+WYJMChpqYoDtlSHBuv1ZJ+gugiP66QshnD4zOHg1aIqFdmMr2FLESlTt94
5qTxGGjTNw4wbweqyna3fFBgc5bITsL5oC5HnB8WgJPBzxxYyc3rfq7CYTyomwuC
l/j6+kEXr1W+UbSiSERdEUNSYSG4qW2SsIXjqrcZMfDs6gkWWTigQJ1wEarM2Q6J
meHfWV6ScZ5Lu9JipYvOEyzsgWTLHwsmn6GVEokmIQbKag60OioHfk29yMpEsuWz
j/Gxbn9Ld3RPJnt9pC6l7l9w/PDhwGTnOkHlu6ziwZ6qrkT9+g65eIUWLtd/HGTg
CPuq3QG6eB0+By4dNiBhtCmlvAiRSYSaQgz/35QAznkXtC/u2anz1qXca/M6eEZo
BZ4q/7btbfn2AzDs0cNMcEZwlQkuv6I52XHViq6nu0PTAz9mH/Nwm23IEQOXXR+9
Oz4m1Km2kSzUNnJHyI9K4J/K60y5gtbD8m396FiW+5y0qJHQGeMH0Cgjy//U6PkV
CcsGcoOmCDwXWvKUbD2d18k4YldE53JhJijQqlJAAbUeCzwUO8KM8RuAcl/wTQSr
jfS+rbCU1IgZANiKnqRdcvVAoULCEUio5HMiaIWVLgAruYZEpLJEL6BaATYpEpe7
M6DY1RF+q7roq3xSVz0V/m55vcVMsbTQlclTKpwfcAkRBatlgsMFdNRFdrZfG7Lr
eZ3LyAv8MqOoZbLacD8frqncUVhphIDHPixzpNZ7XGT0VR1u5BGs9Q5jXGoeMFT2
Fi5nlCUluSnIeQrh7b+QStOObfbKajzXn44gkgt9PEvc+7TB1yhntyq1dVzCyz6I
fy6GU/qUtA8fO1DOcmvamwGqeeGzTVxj8Q0HTl+sfiagjgXMUpvtKHoaiwFXvsj0
qK3hU7Ritmwu+AvIg0pkAqOLzPOWSEDUyC2z69Jbm4+V7ZcztYrzA7VATQ/g0tJn
wdydfSR8TfcMKc2vxTDloKVAY7pKQ9S2HZr0+KZM1FVSPjibZmYzELD9lPtNEhjC
Lop5WDxlC6XyWIE33abMr8Az72OjqiPP0F/vVNL7uCbu01TDjT7Iip74cyPjDpVE
Gpy8uSDmRFceXtpkgc2mZ4iL3nmt9WyE7KUAM26HhBbwOWQXipklYUQQv6ztlahr
oUoHAirpCw8D1X8sneo84wHlqdXIiLAFPqda94A7fRy/Bp/wRqswpiY/+ZAsof1l
i5JGlRrJi8M+hNHpqM9K5KKK5kEkIR0HHGowkgczEfAFgEiKht5T47OscGY5z7R8
k4/lOHJSgxgEVb7xjzq5k4gL+zytuFjHdesCjKOirgMNe9LALhaOhu8hZswdfj/e
eVmLU/1AwG2MGZQp5kZsHHZoqiVg3HaTHyK4kwkPe1DrA5foVcxwssTYW/VWwQsi
MWT5r16I9wARAMhwObkVIf79R3ToVsKTdcguimKwK17oTEh0NyrB+j5SLCOEXowx
2qVFuMvKGnMVsIXvnNo8CtwM2pzZ3vHrIemfzeH67NR6AN7mqRNFagbTPGbaqLq6
mK49+8elNsbhjtWfspfOkwvWzq4s5wTGaMSmuMIC/FBz2j5bpf4OvJoMzogwO8Xt
FC7+eMvUSnhhTHJ3Q5JrUT8eh8ya21d198yoKYHzGmrSpgEmKQMiiIaA60T95CnV
ZNxFoivptU1ymREP5I+IzRXiebE3yJMI5wnwarmVyXNr0i5UH0mfs+D3R7EqY2y1
oBjbhROUQtQMAmy7hK8n0ga+KSwrnoleh2hi8DguarZwn+E8dBARQiQLrKls7arq
YHGIUyf4Y0XXuQ86KTsTFt66d9MK8nUj0d31a4DM0k/gLvI6OeexEq1Xjuwd9U8K
iipRsb3Ij6D0pPYjZcew9pr1e7L5PZ2vwVnT3R51i89Gsu8cRL5lIR96DaYKxdqd
BgZ0hlLEv01uJkxDi1ly16M+VaMtF6k2ov53HJYmR7OLH8xY5J7tw9dYveC7SAFj
6BNBk/kM8plOR3WoEU+s/7kEwCxTwLZA3takSOiv8svr1FjH72BgtAEgasXQx39G
JKI1lM8N8RTJFYzihDm+ReBQPArtaUat5YOM3yKP3DwzfJ8VKKb3zTrrN/rqqZ8i
ZBuWvogoCFTcOZmo2ShtlfvwQocmwbY5kVzGK1VSaj7e4gTcpnTITL4ZkP8HMWJ2
Or7l/XoJ/jNKxISlMKcul0qS4Q3pV0XuY7FGWajuxLXKpYGVzzZic0v+d6BV0xvr
BjdZqvRHBoyhT34GbOfvud6IQuk02cS2EWVMrMObjpScqqWa6hP16HXGFEBg8G4Q
I/rbTAb7LxES63agWVsH+aSYJ1ZyNSl1vm8FD9FAJDYCnoHyX0dJW/DQwOdQFl5B
MnGEQCcsD040P6v277Fk+5twqiemSUCqbe8XktCDhWjTyKUdEEqJ1omvGvwuwZ1P
w7x140aNkAGACpm31vVV+F1OUOTas+xJtqH5XUDCeiGzS60q+aODZopHxVw2zwIS
l67vMNwgvP1j/fxd96qYnzXmKTjMnMVn8SauDfG8+LyIP04Q+JJKYodD+BvBLgpJ
VSO8u+ip1Ky9Stb2SX6t6hfYRRreNwntdc5rMM6KSJZfqtvHcpLgZdTyBIJt+teB
ASUFweplU4SUsS0vL8Lsh75QKIstdihxadggKB8ygFCEi/nhjqtDOgziSDxvUT/K
S2wvCu/61eFySlCjtZI2Qelr4TtEwI0EO6p0g9AQ4UjBx1cvgN/ZRIWiOuPwAVvY
cSzdYXrnotg2c/QGGskxwDGYmrbkHGNr3qgseOkHO/QD2wMZSuNnIoHB4bsDIHFy
3Lx1msKB3cdZeVnlfspOWZkoVO/QZRkhO3iCe+H6tsAZAZ5QM1z7gvW4sT6josyD
MEUwoUO812BAxD5cyVt5ivO827Smw84hVvn0VaBIoXCkNrhNnvGOy1BS3sOEAcYd
pzz6yS1FC2r8tBsQd0xIhDjbm+KHfpsTVCWre5PZho5ILJVmdiG9kJTQEIoSTu48
mOZVmtx0Rub00Omp8vHTlFZct2/mr+UG2axEpPgX5Ql7zmj9ahcLgzO7vyK7uKNW
8msPn5o4HAhyKP6ve4fTsFpjgD1S6kA99oUMtbRiRVRVM8039sS5qRGKOL3zapNv
g/8BxP4dYWbtIRJvIpIck/R8kAZaK2gxf7mQTW50cbjANnnrJzviOo14YHXo6+AY
SLrheLbt1OpxriYbS0hCRBCbA3m2vAB1vejXFO4fgezh69hWx5wHiNBi0oqEJ1vg
iRV3b27ttCP3bOwlIAUD4eM6lGxnyrQzKUGxgMcbKNizT4nYaahiRMFME4XLm5RB
Joj5oZyD13zfd7i1d7cBn44pTAO6i9MdvUpKGRJP55h7AKSMlllDVIJL3NV4s5IV
qFtyNABQaMZKI4+uPPf+Lz3JKgl1jkeZCPVQZ08k5rmhG1xOeCDlafk8XWaS5R9j
xhX/mEB9S7V1nSyO2jHvgg+uo5zXNRbjBdHLL6d1UIIPyvRx0CUFXLC+FMm7PHgr
30tt/r86+B09+CcP82rFGpJXjOteiRcQQdfttwacmwwit5progs75yJ8jr0/dAG7
Ht0/Px3kGjCTW0gg6zpTzqhnVkBL6dwRYgQ87O9hnnxRWuyPmvzhhK2/txsd/eFu
I2cuXgiiseer4blKDmS4JCIsYPnhNjjDgYoimYvTsIw+0NAOtMNZCU2KtqBkO2k/
2VrWkjNIwAL4do7JCrWZRBS8uIG0kGco6u2p/ZWeyHkwaiiK2UbHO2C3iPJr1xj2
QosCPv0oo0SYOxMDmIFxmiwmD2KTUuJufnv6fh3KT+UafN3ruilL2YnmRbQYN3fL
ZDrTc8fxRshsp2cECPrWPqrgEL4Q25V4eNiMfgfWNDaLsdh1rsn5hRyau/ozAv5T
szSF5XcrxaJIXTHZNtokM18xfEZk4p0fX1AUeTjyX14wwtVLH6aX0LnuJyGnXC4E
fImOEVVwSU9JlQYXPr8zNLpJuMjodgakcRFodXU9adHPXQhMcMjEhfTv/f6JSGP5
vDXCvdwLEeFWin0/GK4/whoI0FKS9SQXYqgfLqSzMw6jTbZR7gC4ee93l7gcJxWe
wLPnsNyy7m5UBPHPAlP94wGVeQlSajJ+FKdqGQ+oY14NGgJZB4EBWoHU1Q310mDy
RAjnltFa16QJhHSs+vqR1r+v5QMHgnKltFt9/bO81ba/1t/YWfwTl/eDvXILKOVt
/FMUWk0+EbPPO5sz2laB0D9vlVpe42jVMP8ck6w7Jk1cTBHgystRAQIGfXfrFuqh
Fmg+86UCG51/+wqE0avfDdfsRJSDEfmLxdbm3ZOculid5IQIsbR8zF/Xe2ZEkTAk
DsXxpp+cZdEFdRnU94hEf/Vxz79HOVUHr2ECDXILYc3Gta8dWEeiQensqhxzbAdp
FPvbjRivPAaN6r64bmwf58S3vWiJhOgb+h2C1dOJNihZK2MmaHMW2i776hUdGLmO
wt6wAseEQBcUkTPR+PQD5uCK4ebxs4a1lHA8EHGqd+B0MHYdJvQqQcEPMmqgagqe
mseGkuUHPgLidJYoeN4rKQVEZb1pDbZz166a7M/Dxq+V+BxQWWYmsA8jWjFWxFW9
XjmSZ22NG+lMx9oIzLeZXGnMxIfGvaz8+jjB8d9XQRfylkXg4Krxy5J9pozCvnR8
PUkilHuX0Jj6T6Jqk4LsyAghy/HZVmXClWyD394QdxY0xaQfVeLiWa08ClxOVVCe
qyntMf887R4lRN8GkaGw2P+TRvE2L/c0pG1xxQq2X4QdQxCL2NcuYITnGfBJKK1J
UCG9cCMJnZdvp+UdSuA0cID+f/ejBeYjP4c5zQgxVW+wccV1p8YZFrKei6YCoCbB
/7P3dMphqfQ+VZ82qEwApxfAzEzI/A7GylEeX61dT2HMBsuQUj0u5BeYoRGmFpQK
9vKtXTzXGfaRCweUTi5HGi3MwWDbiEvYPDW/i7jAZbpw6Pr1jRx+c6NtZuEXt215
oYLf4A8PMPd6uE52sEUQDq+wjzKDqdGK9j3/5wNwnJUjFc+pOc7fWl5XJA/o4m2C
VgdvIY+gy3Jk/5JTbs3FdqXazGSu9Joil0ZfE+bU5Zk0h1i+4ZAvQw9DRGDxOG1h
b5F4AcNL5HmI4qGbJP9HJc1S22a1nTm7ydJRcHv4vYbam2mryT5EnxY0xG6pBe+X
bJy9bIgUAp7W+3IQupNO+eoUAaFKNBYum0Ap74dJfXbVMGb09aPtRwu6k26KH8Oc
mP4AwddoJQiwq9wr/h4T8vb9pDBs/X/5stvUImmyQgbKrX5tbb0+YP+3SLKyNIhD
Ph8elciyUX7uB8J20fjsZ6WLuMPIPy5a+TyIodaUehol856nWJK2wM01ihfkBHke
iV9G5XLG7hGRBzA6yFdNCr4cRrf2AgtP4jQAJzbCoFbEyIpUtYLZB2C7Auzbswmq
ySk3MbHJFT03CGN7AmSVrj2xGHuD3kWr+XmKoZr4ZQdPFX2Nrex5tMK61w9KhDnE
6EQ4xvMmDTZb+7hWSOm2O8qsbuQEJk8MOKx9SeYx9fKii/VthGq3RzZBHA4L1rJk
S5etIJZ3kiqVHOx7pjzWsPur4315BdHdf7y36gmrLTkKGXbca+B5u0AZtERGOaC/
9cuFLB1Kmc/09RRP1UmXHSE5l9dMLFEf34QfauO2rQSScO26HiUgIpB+4q8FkXiw
PXvaUgZxjRxnIgWPrsy/5FlytDgEu4EwIBHmmvvozEjZAk3bD/Qjb6FiCdQhKDpt
Gxov+DocciKxt/3IrzQsP1p3mvprvQJLTnIqW5n6eErO76XAfUPedEPP3ZbvH1tg
G8mGsRwKn6NeH/XTGloJZ5nd9qnSSJQdbG92jHBC0ARxZCxFJqqeEkYzQ0BQ934N
sJrU1d2rJSmqOhTWXoJC6sa0DRPvH/RNHkIaTKHCkVpxeEj5jPolTzG5l+8RnwA5
o9+KSbLoPAK0k0dBRdzVb4jr8KlPczKbEJWv/CV0LDhOWtgzRzpLsxMWYupZVR+r
EV0bshH34PN81qh3T7YGiXjl80St/xDLln1GXf/2fQKoE+oaZkJiahJsFr57jiGp
mnYp61Vs7n9SVBY9xhIe6in15QuO1AOR1kBwwgDEcBY+k8oDOnYRH/f3DtQ2Ud2m
Zw6LOeYXAdyQk9YgLcavN/RIKsZL2g6OXguUhpqSVCAOdfzM64GZfF+2+HTquFYu
DEiOwdmWFPYxdLyHnZ6WSkThH5dmCQ1Bh4aaVjY21TtQ4qlTZg2F8PCH6+5iP96I
9Od3HqBtEzqm12iYceOlP/agMnpFcaVEMmXZSgAoSbErVCkFrQArQjoK82pmx5k/
/iBWrmjREXNEWUWqCaoT84FIgr1e0nJDMda4+S373C1SxySxS6GPHdCMRbXYE7DA
NJm5c8Hgdlo9akaa9W/a5KvVgFJoBda+cEAeq9NhDJY5YFWXp7xWpAiuBpwxNvbl
8YIgcpYFSM2yrADPmJLorEmcu9U6BPtHV1o+R93gOarMaf6bYGmevMxImrVWHTBs
e9m/HDFMwPT2/PEEs/JdCcWM5fLqJZ/h+8X2fVqrgmL8qmWnDRMmuykf1zezD3zB
JJJA8gTVH2whey7B5WSYHnQ5xREqUzWOZcdqflNTco2cns4mGO0E6sNDy+uE4GB+
eJ9KMeu51Q8uf+Gol5Z+giV64mgYsabwD3ClODqN9Q6VlCf/Th5N2aYxiln5iaZ3
CEDVi3AV4T/9444/fKyPw+siMP8i3oWX4k0MUCuIQ2b5H42RhkFqzdNFaR9XLyo+
3kT5ByfW3M6ZeAgryzBrN70CcAzOyMvUNB4rleJ7H20z6ndUpiSvsztKdZJAKGoi
JW9zWO8mbRRvFj2+nFG4uJFNSz3ymBGLI+Ohvc/Aieu+Sld0zZwZZchIN5y+7Ior
EFHoD3OSQ4ak9Dt/h3PO/aRG+B1Th8e/NCuK4TcqaRLsDn1KMXo9RbW15FIv23BD
72FXRCGJ5DJ8tXF6dwxNdyOmsqUbc1yyPCWqizwQ+fATNwlZAXTWFdsRG9sAQ64i
mWR9lVxyELB/QqD1FQg9zuCzQTDnh3DrI7wkfBHxX7xzXJNEF89bq9e5jAsN3Z4N
Gyh2nTQ9YjEVW1OBr+hQl9cOwjlyR9skJ+GU0bl6zDypjdlcKc2tlplgRj07aBFX
s9c6lrhhA3WNdK+omC99F/gvvOHwdSPBabQyu+vmBMZ045zTrR9vtbrkkJ6HGKPs
piMnvz7rc1hJC8C/tS7P1Vjyp7f+NirmyV/+4BXQanLl5dXpXwD+zJjnmPy/ty3o
8GbuAWWPY2Kd2FjkW19alXG1LTK5S43H5EviHAdlPie007LJDKmA7cTNoqAJJLWl
tqKVr9YGuju/9MP/El6BCDAkjubKqQPEEdutYf7abm5XP9dvAw75hEHaTvPmSRqI
4PfETlRnTPSkVNpXhM3omoEoHkMpDnnls2RTnOlhQPAL/VbMEMLOGAK0Qs4LSWpa
SIKSMnvIWbe8KqEwuEoDfyPP5MghtAciHLZgv584tzwfPzvl8GGTOWxpW+gxAR8t
DNdlHmxgujd2iCJXJeMMl1AyggNgAaphavIMVYK9iPUYTobBSGs5U04TNFk5xXoX
Bcl80Wxb7Qgpfd4ri1L/EUYPXEu5nX+P/BH3K8vU8+zzn6LqRVukierovFts3jbE
UPbi2/uz/06Gebdwm9d8OtlejJcyV+q15Cl37O2XteJbs8DCj7+Dd6GbdyCV6EZH
B3rzdhy2mroTQsELuV1sX9B4kl1mi7c/X9/KNnh87aQPDHROqOIssgnOkZiOCGdV
mxnT5ZprXON8nltqlS1VoAPYCkMsrkCUm6uNW+J0yxpBcK+apO+KBzXaeaI72mPb
W/JtD21FRaFEtLATOOcSbtMiyjiwRzFhCLVnjbHJHSdY9EC6H6kVDaLrDH/sAhTy
0uWNmjv2UtFjQuOgD8R+vbmlILkJnaMNNGk8d7EcfYBRBcxeDhZKVKrpfrvSQ4vi
BeXHQsEtkt9BgJQeNVO/3O6aFHRDt2eaaz/KHvQZHNV+5a4UMWOjrFjsYUhZpgUo
5Z1LKobQk8emCB6WQQM2J/PpANyOPUJhZ13ZJwgVCKwpdHfwVNPhNN2gUUh4hA44
byyPOkOzcWmIfWjYu6Q01tMWj6XFJ7QBWxAbZzFRcKRYt9yERr4VWwDW0Q3NsyCU
xNGka08RugHMd1d02PS1iPmyxPfMJIrQFfRYiol9+wiMv38WVSqf0AAfsG4DBAHd
3eJ3yo/keCTZ9cTyIqxVfCoxwg1cLAJL1fAfaNCL5KzKVGmHU5pJ2IsuU7m5YCN2
x5xFFikkMlzEEwmVzwuKw33kSffm4Enqd1MbA3Q2T+mt8YxBUP9gds4llzaGOIoZ
6qBmxJtGLIDZMSVx2Lmb+359jYnfzh+TSVHZy/BtrQ2ogCEnTnfXPylRmV43vMZu
G48jir84CV0yqQfgy+C8xUdtmSzon5W62fK/V4r1RvnFCZT7kO1iaj/DRqjgLC2p
RvW+CzJEc3cWZqzp4lmFBJfr2bV34I8yihb2+kDRg+QyneK0u0NaLt6aWBtPxFMA
zeM9pKqrVXCnLeupAexj05b07mciagaV/l/IFY0irpOzfg9HsIjHeChPb/PL2koq
W8T4Bt1/lAsb7aW3BVfjl0FX5zYNGNGJubSgjPEuCDV+C0EF4lQTi3IxSPLDp9LA
xAODuPrMoFQ5ioO2J5tmKLRchNENGyaimPSfLYed+Vwpafjf4Q8x4jlDdxRxjgBA
N5Geol0tc8ArHGl5POi1VZ9XsmKDrw2kV/wDKDuNyxVdD+bnN1FE472zubXjE7Vu
slJEll4ZGbDdIVnv6AvL+gVE4MAxnCgkhXlibjG0jw92YVJOHZkrgyTsHc5u8CT8
LEBnr8K2XIbHjhrsqFNS4cZ7QEtj1KPuvs2ghoHjsMJVlPtpJbwDQ3kq2AV0rcii
gnVV1o7YMWJbsconj5ZGVzCI+oPpb5HiPSleTTUkQUbgJlh0aCbfGiDxm1D9oDLQ
TOrQPNkiKLuDRBxRIu/klNpuRull7mcns4GKdQyJTjjLalyWfTnbN84/KcLyl3qO
u1De92J+1fv8KdsHj7mGbIJ9SjRExxK/HSXrO1WYAJFySE/HZAsB9u+mMpVo9dmL
LJvRym5q/uo43jt6FJdTH4SvWWPKTrHtpdVd1a5LdGRoP2hTeawO//N7nQpQJuTC
OBA7kM/ajVjQa495AcCIv5q88UcuX1E1aMZCqaN3av2OFyS/bSgclezG77kKIdpN
+1nBJgr2bOAsaVVuy8G+0/PTOQY3lGK36B7ZNUf2bNgOxJcCodXpQitetLLO+olY
8FOyQbXwm1u/06aS44BKncsLQhHMQ+KDcXFtaYYjnvGVmU3Ec3bywEZRObpZLfsh
pYZHDKw0M+4igygnXxYKVFx4tCyVLx6c1OGkkX/79dgckQw+3O7AHFyoF2XgX5vD
u4dJBp8dy7R2RLcxJ3pJvvbhBaxojdYs+2WV2IFDR1hzPtF02onUp601Dh8FzQ+X
Wwxf4jp4zl20omgLZT4J9qH4azgwWKT6M7TsSZJRq9fzfsR61Mvdb5zKYQ9bstlw
0lLzVOrhGkUgkn1B1HUheBn3yXTiJMoFbOeTAfKj16pIUi04M28jHV5jRcidMbvc
0NnVCADQ5RSv8atcgeF/KU7BQjDuTf2YeIcQWqhrGdJyPPl47ZdB8UCnZF0AvzUo
Sqilbl0jeDqJOQeyI6R04qIsgR2PEYtDvp6YFSbOcU0qKtFaXuQPD2Y/jYCRbq4r
bc/1+BFrAX+29rQPC8AdAiXK6yRerxEGtOQE1A9pz9hGuCFgzf9EIJyaJkMkiXtx
d/yLFCoIyB7Ig3/JmslnqwkrtETt0wVSAEQgcTmwsngbwCLXoEFK6hh9+izGD+FB
Yav/ebQi/zeyrnW0zsITewZ5Ct4wjPrcJqYBATtobSNp/5JAkTWqHckMKrjCEmco
A3LvcICG2+xwNgJzL9FGgUnVqia9hhZ506/tv8U1VTxPuSagzORukchVy0LtJQ8m
y/hbuE+okoUjtx5o3Bg9Ki8GtbUDMlJgWlB/NjKunE/fLg+9JVhn7IDkGa0HOw6W
CHXVzubb5sQXMnCmRdjZPKERTdujxcDlbjlgj+T406q5dx7GzFkRiYjH4iwyCxIS
hiYV7xgoo/nxvnRjSA3YaAlj9JsKrLjmE85+NbvkjTZykS7zrc41V2ptvhTsQ+2X
f6/9aTzcJqzngTZancSoNKdiriYMMJfJlwf3RUeua+wTagwtl2YOUpsDNtsdI2Ha
zzYnrAUi16jutpS+k9YNfgIjv9xHCqXA94X5wJ/bL4VnLaslq9nzP1cHg6SVMGUc
ERr/iaouO54+JrePRUU/67WBVoBQdIG4sLj4lzBL/BSIw9U5e0ue3HQN17cqNA7i
mNobGBy0oYBh0SlTTnPQvIICQ7Z+UotQGDgY+zbz7D5vjEnZfYC6ZSf49D8UZf2u
TzcbmGjM5OEtnZx6Rm+5w4S6gcIpXMgjrKf9IPKcW39NQfHBDtpL1pMFDW/zv9Aq
WbZ9UMAV2ytKbl/reBNoc4AteaQraVvzHtIEoaZslyVjJEWy1OeEW+rUsu3BxRYQ
209+PqR7ymz5iF77mxVGOqvMpZl00UHOTIXCJEU8+0gUvFADRfz2dQeb2ECNom8I
F2FRLcTvBRnJ6eTYujNk4a+/naGTkoZ1Pf8hrEofjcVRUYaZfYcqX39knSX7DlMB
2wC7kRij0DpADNPinwRMxWQ6UJu1zhWXaKzgSm3MgO75YjqrVNgMnmZVEJgirOeL
SF/tVMlcAFPGOqj3pjBiNlRDrUtOlW3aFS2ihuipmT1fHDRb281TryFCCG8xq0Qq
/28Ar/cVXcNttzTn3PU2fJ9vwkRebUUYND8oPdTFXsIAiuhfq79q3NVzTS0BwCyu
PFdbOYKgZAIW0aex4n/xPPF+Xga57jo8jsZaoviXgXN1b3x9xbsrgbFfnZzn1XQq
WNvs0aAC+ndHjXtVT4ldimQon3CSMAXV6uX0VDuxVCT2ZPbns6wBRQrxVf8oJXfo
wWCLJscNDuseph8z5Dn2lwVAdMxwwRsqooslhGyqSOhrk8vXk2qqUz1G2ePgZrZ8
CVflx4JO2v8A389ccAao1PstbjiyCEkv2GqOZvomldN95vIpsJtQsT71Nc1/Qsgk
L1kaK7PZBMDf1h5/haY1TsazZi+zF+/b0whz5zbe5b0swtybA9cH9YPiMPNbleUP
E5oBlY6FWpS3eR63JdhmVzFvRM6qHRqci14HNJbei/9gMkyZjBcfmQDQf/M/2PJF
bMgbfaUYnSaEEQPVep3744vvQc3XKB0kXDujl+5c3RTtaX2EwxuGUZwsoNdyPKDY
mFq3Nn4YAiwSgAKrN8IYfGY8160jaLUspUibQNj7HSfWlmU0oe6CNxgeSkLu+mUX
a9Z3aiUdBH/8LDLWFCd2+5FqpXC5hjhRTZUItQmiugVV2dIMeOG77/52uZvFQ8P5
ducjws6g1ImDmrXrlNo8N+FzMKCY8w8qiDTqSoS28zbXVj6DjbcV9Xme/sbxn5ug
RG0dP212kUQfgNtFxU1xZJHvCwLWhyliPpxPczeJ0oAWSBkyg08anFx8nV/RwvWU
gNteDuKCqCARL+/2Viuit9jNj6EWFaeX0NvH5Wj7cW6nzKDrs8k7Cx0JlKaULcXB
Qxuenz2QEeKSY25pyAXQpZPBufNXcqhMJcw2c9xIrcy0b1FxxR5Mx9DOvvx6SYUn
qEaK7CTU8rR683yHdqKo/UwNwwiwFDdvY/BVjvw/FWHOnKQvXEy/Z7pMXowMgvKw
UTqxIEtvtkXBt/QQiRSvIew9iJEkN6bupDKpLyQ4yXs+BQSAB8NsqLp1LQVCbifH
qKpno0sWHi+ItxuCH7Z4qRri/toSykUZzJSi2CFnb0bNiDn1NhekCOZppdGidnYN
xn2nUUhrMhZxg/N+Mqgxa+N2Ae1rO8zJFASauVct5bTc1TWV6WcLeDy+14+9Rj1a
BtaZmnxg1A15od13qgEkw/iXayf+JfrMulNRTEJqlwpZCgnSncPA9HBtzwyJzIwt
GLlzDj0GAe5+DjSTCF2sw284C5je6EOS1ZzGW9WmQxPR8PZH5SmBPLFvKf2AIRit
z3nQYlZBVOVnzXLUGzUjzTm8U70Q4w2NtJRPcHv2QP58hlmTrsyESwOSg0ge+CdV
MXT9REem0Z+q/sYqbNyrjnZriDYiNq5GlXM7Yb/ASWE+/fW6R9HZaKO6DQ74ZIcU
1l4Ern0lU+x2w03z8Dsq+Nmqc3DlPi4kWpbsWJN4sQR2khZbdIDHnNxPSJZjJBAG
Fmm/ofd2aKF7KGO3wsjHy7CZ/J47vW72ebwheZsekRf6xFDzGBK+SQFmCAJX11XM
zOhOwl6o+9MZ3OW+Mxjqw894GfIdsHfDVwT1NsLFvnashmWu4k6KVQoxuSsbDsuf
GBd3CA0UjU2Tt4WiXQCYIUcdDcMDSPrcWCR6RG9laZTZ9BcFBLUYNRjUWqhwxNGU
9rSgdry+eJlLDykVTS6PDSEQIKwLSaSgLMh7BYZuFDjRvhNvBLOTzZpBEmx2sfhh
AsMDWkY84WOQlCkbVQ89gdq41FLcTmCgDLUNBq7bi4K/J1bhdy13tW8vkqLZtVDZ
ibDBknooVUU1QGpjpA/b1dh8e4J+MqVhc++wdtLDaLnXJaylvk8u8Hnvvatj8JzC
3GmrGgeB7kW8MnY1TME+Z+/SOng6wpnHl6DI2HNWf2vtp3yt/Zgzk/YC2hMGydLW
faE2Q+eTc3UQ7jQdHIj/vFaeuraf78Ae9J2+B2pL63yFSsEE4I86VQaJTwBMqcMv
r+Q0Ho4cBtzT4OE4VEEKoCHY2+c0OrjQmaUT+3M/plwzI6WGFtrt2SVNuSDd1Go+
Ua75J2UA1paliOjz/g2PP5XTUYgCqUZrUhDADBvF+7taLS5Z0b792eg9uFMUjc05
jRzQ59EVnQT5ZiARq8avadPCJ1DIEnYEz+G2yg1Fjzr0HBy2FU2Yq+AzwTZL2OgT
AIfMd3TR/WyguUnCVGPWVOd9xGLM6NV87ixc9K2VFy/Ez9AIW8/cxUf1QPUNmmdo
eqDoNg5buA4Q88Ew9IFfa4cM1Sjk/fvg3bOwibGNNEeZXg7GDneWw8sDig55sAxj
Wf0ztwS3wuw3FbZiy3zvrMxrXyEtcPr8A2JKSzGEhVvc0u/fjdx9zHDu28lkZgpe
p9QlfHORqctPF3yZiYHBI95TwrT4p1tJZ6gWe/cW0UDWkSF88Qt5NfjsKP6bVT64
4GmfEOks59y2DSPuI+HopTZiRNuUGKvAXolOzeqfPEx3wCXfI3VCznDT3qGBWCN1
FD8cXFDpXp3wOqxdHxc/H8cF+iF3PTO9TRooWJrv0nWC3FRVyraYIJcSdQaElR3H
MwHEJtyFCHmJ9KCFWszQ0xxpxgpnrYe6DSbLdK3QborT6f+C4KCzKVxBCmvUFraT
VEffKq3XxAN1WK7eyXKNx7YdyuZUI80jUAaqyP2ePUTwDDuhBXKOJ1MQ0WcLJ0hp
/1JEwZjD+N6PZutdDI7v2qDOCNsG/BHbkySPEqyleW5FTm/oFlZZAgBH2YrD2aEO
VOzCAC0H1ourCInpFFIJmzJw/vPOjQndSvAA6PjeOtGT+aa/o5rR7G3XZceSqnDi
DI8utnGz8TWnFyeynok94nFTYWoTOTO7G5eGG+DlKnkdKGJDB4QrzwmRO9HcVwbf
19mcv7c8DYIr0lMeQiniv7kgb/UFV057CmMGAq7IuruhsbIjZ75ZqJw7gKZBWict
ooCklxyNXkSuxV327VCumEJJrnXjyvl9oiA4X3+j636fACffpstEDslaPR5vStJi
5PZ+W5hBF0C+167Rhon5emVZ6DHBiW29yl3yeO/RFML69nJNXRuDqpyjtpGAPcA3
A5xzv5cP/C5xbkyuGPP6pHsWn8wsVnkqGA3EqwNJWcD55mOuLk9LY/vnXO57hi0Y
z3M/FNu5wFhMX8aHeWVwDVHK4QHn4UUEYGSwhoL94r08miMa7kMi2TfJw/6rWstO
WIwEY+EE3uIPugLXm3gAoLg/tDN49ir11T0sG1j2Zxe0PP/f0FTyNrmcKz25YytX
iRaoA7zY58h139CtYBxtZHNKp/aXXDAZ1p0uArgrjRrPVBb/KmvyfZF+R9NDoCyH
gwbS4AFyYdwhX/gcAj+u3WSDexQl72ygtWoGs162qNcQrb0ovzmL0YsuPjC1tj2W
9BlFP+/DkcxPa8VM70YCaZOvRr7Ox50ViccnwU6zs5U3OkjrR08O6hSEnLEurLyO
U9vWQ/ud81UcLaDyF3Im5CQwYnwzLZ1R1NowlTvgWz3M4DaeLFU21NYYCATYIKJx
nhBa5Fteip++B4nE8TF8LYkc1sZMvjGLWKu9nTtFgmvQe0daof7W92HkNIgR3XeT
tjCfSi8lEzp5WOp0G3AGC9wnEfozQEpkom7krznKViqZlfZW59tWkbI+Yugw95BT
B4rhRvjSpC/sN4F8E8jPWFGkAYUBxagFeKmgzCy0bZNaJk8t1LSC7S33GaP1Qu30
TKF+pfQKt8tBk5xLwKjzU5H7a9HC5o6DWVWQ0BCE5UoL8QRcaQHXuqH0W2x7KEM0
+JMq4cRH9jm0IERYDZrVpo/l9mEL1qqrhR7cuCNXwDUpGq3mURaeh8KDWx5+LOFk
z0NQpE5GYRPLiO1ACQzx3AzJgd52n7SO3vt2dVGRNbiGojqWxPT75aZ5MpYWS26o
bJO38/yvZ0qzCGcpRHp9bemw25ZwdFyg/590TfktqRYNQNnl2WtbnDZYx5FfS82t
u/5FIj6p84fQ5pm3EVcFKi9mBP3b5VVrXtEow5ZtQfKpC9+lhNjjD9kwzcEQQBzg
MB9D/NI9nT9CZ2XqnuF41kW2Qh91aS8/5WzcBFTMYv8h8lK+4o9bJzMm5TO9+4IN
e7UO11XClRVVJxi4Xa9KOYVlPF1sk0is4kJAywC2knMQu4Hrh0RbtV/2ur6qgvN+
5gUAeROF2AbPbZp1b1Fa5BmmfpCwtOYuf1aMV7QZ2yfFljORwsYUVXiREMZZdnSJ
JUtXCpX+59o0EcQBYdCEJt0a/yhgEvW/iHiNOfR1HttV6TKp4bV6RhgzjBaeObMM
STDJz7m2b7Ot4JZZ8bD+jHO8MDt2WyMikrIb/gXDKnwzecr9YZBfN0qmXbU93+6C
NWSAHFMchdmFow/tNFi8d7mo3c4mGKkqCUg/7P1K42VCecaG5MdmzlKAW4Lpi6kp
YSrxbdTaKDHhNwvWwq840bsI8nVQaZkR60C8XwfxJ/KECNJNRQqp7l3FPXyofzbE
292mV4ejT/oFidDTaMWh4Shfozp8Tqkrgfh1jJJT9VtWVOUnW8/c7oIRA7al8sI1
ivdFQvlxmwNwleT4ODx/TP8P4sEh9knfAF69laptABgbe++iu9BMhpIgdlq7ceRw
ebeaC364WoS6U35jFZ8Yzry1MwaS3HNBDqQpChlzmY3tTKrrmbqGFrivpLIvESIp
8JWooTn3oTQoWx2e8YsNve0Z6eKP1hofCqZoHjfqABTT2O8yWCw/b69uA0aPOsJb
2RU/9M4QfRcISA4kWELkFECjrw3yKi+DuH4gz4XzgH6xlM8ZJbONvU3m2DOC0yV8
F8LPw8XCKKo/2HpwucL2k8wBk6a1AHQaU7b0Kt4MaEQI/ZJovOtGDPlv/zxura1w
amSUsTlHCDxnY6bOXltVnTYGX4CdFKXGJvwP6aqg3mw8BmJGYG0tPsLHxDN/BVmD
qwavJZJwiotLxjVHSHAl/lBmhZZgJprY1C6XjSvASG7MEib0EtjdrY37QK7Z5Ued
`pragma protect end_protected
