`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
n+n1HsXd+109G+3JNFuhHHcEqcOjJqP1SEwHh346xh7pwcu0/dnYheAsbyvbVXcy
cQT1dA9Gs983QkQo0cJc8tujs01423Y0eKeAlNLp1MoFm/aSzNjBHXfylQOUrJSh
bB61dbLSfeGx4DoVnPbnZvi1kaKBFWxmFuxnFF6sfzY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6320)
etH4hLwZRQqT0WIXG/u6ZiAfIyt9zuibuyKjK1V8JeYdsU1kzoajYbdX5kzAQcVB
hkiD6yM1itc19lzHlPqRlneSySB0nF8zQqFT4cNfFaR5Hyd1yHMMIORR8bTI3jL5
7k87O8QEXzxNAf/RLXp3appscdF06vTBzJXfydB7RBrf0mE0TT272lp1GZDRuG4d
nlr1q6dIiGVBKEeL2T/JwL5e4zRmySz/WloC1Oyo7MT3N8HKveBVXO7tZeFCKAtr
83xfoMhTNzXGskTLsUri7sWgMmlMf1J5TIjpYv1SWaO4rgZTF5fITEQn1OqK1mMm
IMbftYg95Wee7PvuK2iq/+l9wHMzgXIUkPg3Obe3AtdaH07sO3NO3bPPVgwShQG+
lCjTaURL12ewnPwe5bO2QX5r/EGC8GJd4adTgsRD5kNo2g0t4yJLlXi+jn6F5dtp
A2uJzmkF5kEDpGd2QbjC4QduWs8A0/q4LI1yh/UzQgBuMaFQpT8BdF8UWG0T71n3
wuFK3X8B3+qFCNttBXCgpTPVxtEN9eZ7VaczORBjoDwZgEGzyFWfGq0jOhkyUmpf
Pzv59MT6ZnUsuxbkufrUPJJPcNbtpf1hB9MoToH750Xa4EeBs90i4XlUxO8S9YEN
1BHuIxt7JkcRQWX+n9wcLa7aaVoC/xvsHlQM8v7Hilsdk9Q65kE7pLnv/X2iB4V3
qYfXhe+YueHX7VZQeXMdy/vxebWLUr+F3Tw8d7Tif6SetLS1V0hYuYy6iHVM4aub
p9ggsxnQRmHUZR8ILuxWrl1RC6lJtjsczkfO4POu1oKGkqETxGtApRAp4mAV77Ua
1oDA2xZpQAK1GRzma/UXwmmUwjMNY4KxmSw2tlVO3ATl8PB4P0GE8+/YFNknJDLY
3hLp+bH0rSzGn/FlkcvLxboG17xix9pbTw0wiBpmWmoWvjFdkEwKWBcYrMD4AeS8
mrqKIQiJLL06YXXRO5difWFrR0d4NXOBDTabrAt3/HbXDodwEoTCZzjmemQixGw1
HX62XvtEyvwihudhISptsWKtVunsCGY+vwXN7vpjEj9/FuiW8UONijN1v0SRzLRT
gTyipFhI9A52B/cK2eKuRpdXiit7QO1zVWMVw0nzBatP5+CVWVYkHZx+lr2RwvJF
s1FloS8UjEIHxoly5/zQGqD53lidq2dlvHJeKkxnNTZuj6DNMzzfdoXWVJ/+SXND
Al3T03Y6RTywbfwYx01qyRc1LIbpPSrfosMPCJdOu2RHKaCIEjTBZxI36u655WUx
TJoJ+z+n7mEK1uw4/uXpVCTu0fSCB7ER7Z2sPyqIChRpwjE6/XsQzgrqubo1unUJ
MTtWdVophieLrZRt0OUs6T9/z6eYz5wkSqDQd3b7rnzcoTkeePOJTjxUzW3RzDHC
IAe9JBaFo6ZsOMy8NUlXpSDILZyuRytRo/Ni5zQPGciowoJI2gaZZkDSW61/YEW0
GMnTwVedmniHnPhNRbVNbHKDIW3IVpDy2mJCG0gH+0n4iWsjxLTo0L575MqnI6oi
JO3o53LHPuVd8nwknN4nabonXHLusAnvav1art5IViQvkuvXRV2SOKY3cLadrwDl
2zAguEuXwbsymRrYng492VRUsn+ItfEE1c4UJmGC3WMUVp/0nEzq0dkU7n6ojDS7
nuX5P8bHDK2lEK3kygcHzAOaeWk+1RHRNOAVqJjNiO8s/acLBOo5b0HmaCFN8DNi
6YIuSd2af/YX0yLBqmwcOb6fi+qRIDprc60RdHi1ccn4kpjOw2LF8q3susxka0p9
pePLguH2FtVD2xsPCAn5AXh348+oI8fYkqnqe1FhPX6PDqe8Um285TXykZgMT7cc
G1vaF+vysIDra/6w2SIhKjS+9izLjfbb7Gk82g5wQnyc81sNgvWFpWeWiNAQO3NF
eiGN5X9T4Il3lr5B62rxxyzxcWCQx/A2DbPs6O3/PMb93KlnB5PPLwsz8+V6N6Jr
MJ09nNTwLrc9jj52lheBw7hB9LokZCmJ3IgQTxNeRICw1TjgrNB2FQEOfvXCP4qZ
2CBUS/ZHnhrQFEluE3xH10RqKZvC6ms2DRQH9QhdsgePDyX+tUVHEJghwU+DrV8j
RbVK0ssSAFb/X2Oe84UFta/Y+yM45nIDx1mzAc0l8FmXy4Uf3V48rmNdGxK/QOqk
LO94k0Q/sK92DrG/O/pLLwiyg42glb/kOPwN5SyoN0N1RKij9IBnX2zCiA35q4+/
oZCjXJ+/i9u6v0IvQ5bUFonWhFDRq6wPjyYbmhcQ3PtScpatmjzNESZ6TQOYUm5h
W+JF59O4hzcOFW6eXzPtCbi6sfbYMZA7EHfH7fNGaikchWPpsk1r3FNMv8n1zD7t
td3XtS+P2etfGMkrWBsCY/IPfiiLKiYZAFeDhbDudF1Rg9l+lvdBPObzOMoQUZ05
PW46YQJMiQl5f2GkH7v2XDlKL3Y2Ec7wYMqmhAN0eC3gOzx3GsJe8l4vGVmIHAj+
ftUksYvin6xRuqHVjSao5NM1b1V8lsXFcmZAyoz7a9jAzAckzR5DfC+LCm3h4I0K
6w7tz/mUn/IiFNE9NOlcWsavVa+hRID1OPUMBMnypk5mD4B2EVVu2+SxIOMbRiHQ
0oXcDU7oSHadUn17kfvz6qUXqAHoS/ZqIixLXeUbX3u8+aIORtgTdC9hSca+c7pw
IJZFXpPCGDa88r0N1KQDyMz8LzXyeRKKAROLy3kWAAG2SUzn35I2QSVFylhfgoPV
9mXUjO/Lnms/SdKAb3pS/M+TT4VcinNLIOBOhxQ/sszM/5DcfMccz2IKHbcw3PmJ
B+VDWzDup3DtCHVBuUsDqcbfN4JGDlbj83cDT37owvbWcD5bsrsoLNuF4ZP6FAgm
lskhu7Lr88Yz23QIs+GHDhk5J6OxqwMiNwzahHAtrP4FJ6xkZnbNbVWslp3CQDhb
wy3DU02sbpInVKjthF8dX5osBJzmMip6FVRxtJh1y8sDtw4Ou921k4pRBvhBDJTr
3APlYcoLpCOpwgGco0f+Y/Si0/k5RcMJ4+TYy51whVus3C8y5vTCpbCrym0k5G3c
YyRUEcMnTRl72kM+9CVWYzidYFOpm5TRKl+zcaCS3JdiW63YeeWytvb33GAuQpbd
1ZWWF3NYPOOdgxXlEPWPn1X5UAaOMmivE2yJ4vAxninBK12BRrWZVdb9FGPg9otJ
IZXWj0sV4LRVM6ekRlc1OS1RDqi7zoTn1Gr0NKOBEPjWJfY3sdT2ZCeuLKKBo6/S
fkxK8IQHVMhweAU1wNbS/UlHZqvX/szPeOW/Dp3zon9o6uIewaeGJCstMrAY5vMD
l6L1Yi1uQLwQRInYPuwxVagU7ve7fKLoXkORGZu1LGgPzQa8MY69lEzUBYiFcfuA
uohzsWtNbd/oCPhqG82r5vqdRn6awen73xVNuloO2AXY28KCgxcsWHR9wAbuz3nK
K/pmy0cYZh5UJUVxmwmM3OdWt8n0abVq+fEUB9xVznUeLKeJpok3UejhpYwDRamT
wbMHQJ2KCKGB+FfUEP5Ob+OBSS2RtfC05DR4E+w0yZKRzZUg7E7uKOSIs9mSGzNI
TE64ejlc2huzuqhvBCv7hwSUHuett9GxHzgtKputNQODpxdRxdOdLwMP6YyODkZ/
+sh7JpI7cvljYk4aWMIhlCuyw2Haet3iqnV1CIi4kAuFvrUdpcZcN7ppEnvQovr6
lLALKLG2Z+6bzZ0cNfbN0+R+LqTZeSp2iPRbq4eq/b+zz6XAT/gZz8niTrcV6Qus
p5XTV6T/QP0nv7E/tIQ0vW8OQUQ/sn1GAhGByN6u5R3/q+h1NFmWTPIWHYx7R21J
8oKrulufremkw/VkaDzyZyaRb0YEBNUtyithN8Vzfiav1T5NxlgTyAA6/gNE4+PB
9J76mDWCmifgrLJxIXbPkLD4+ejiFECOAhHFHnvwqBCCxs5xrr+xNEyi9ndYEdWR
4cuOeRdhnOy22fhJqdjkc8AgYVSbrNWW4sXMHERrbZ0kTmElnEts1YOg3/FYSxy3
UX6VhFJmsqEOnIVInZfg7MyZoVjD9laUm4N77R1Hl3zOlGD5PCwMg8b95R/xdSPU
KhAdHe5eFnT1SmbMQZujIRQgjudrhQE/GMG1wxotlLub8iI0njzzTotRFu+NKzUK
QS6X1B3GsGRueAn0blH1GvcCWEg789qOYsnbYxMluJAh1YWUfplJk33KEyPASu3m
QtCNxoXDm9x4dWFvNoPokPTVLsyzxsRqSLh96wsyBMVXf0e7N7BTByEDiihm4Nkr
nrOjCWGm1tfIkSZ+0K5o/EMP1gNsvbQ2xkzNNWWnC6nfXAjHvQ3IdbTWl6Oirql/
MRyc6rsUzriB9fB9q2RBU8WBTdE6XmNuMBZDl1jh/Ppr4VHWKrQuMeEEF0bOtDPS
fQZjIgo1HUyES0lPVDjx8ZGGDqj56/ZhYygYoRfWp6FhuIJJIOP9gg9QGJOU+dbU
xjyTFMEB80Qs2XpfDQWd8ZytoxdXY1XCIA0qQvafQxkrJ+flzN+Rv0nWM+e4mRV7
qgFBw6vEsaASw1omsewcH0JsB270JDTmhFID32S0+42qskIE+damItx6F2VTEilT
ilx9SVq2GKNa4lhjyli0X3gGQaWv9vLWICYlMAmlCPsF0OfuyllcbovYSzn6kOYi
1VdK882h8+F+4xzCOv1JmLeY4h9xnj5f0LHo9TznzViXo7ghTOIOBV3C2cZI/kyR
4XLvoOHQgVg+HvzpTYdgGACPDoYlkFGd2rJJQMWk8dM7gGylwhlfVpodCrtMpeiu
UxRrbG9yzw/eECIQ3ibxhSpC6VvkWS1C4Y23niTRifQDTvK9Fq/F54TEgc7pQWHT
l78eXg9hqBmYR+rF8eeVR/sTUqiArAI2xJuX09fvjhQ5dr3q18tmL9g7NASNVZl1
fpdrtNomnezADZXguCLqovH71qhE147S/hpgBd34E48HYvyy8HuXv7moVX5sdz1M
TIf1KZ/+ARhZFB0CeYPG/j4VrlJmBL+d+3H5/OIKzWN5043G90N57+dZLQ/Qih+o
WW/+JUCEJurYEncF86dHz5yKeHU587fIuBl3oQEM1A/iPlRQmDOBMhdQ4mrjlK6b
44cRoBBpc4ZjhO0SX5/pTYi6vsTjg2xOEVA4t8Me22Khtc+DLoRcv/8aQXFHq+Te
2nmXHAM/PIrGTJR3RfBay372rNDruy2Tl5aDK1Y8xzYBZmtnyFTgfcEALHfdkwPP
ptu6gZHnjkPN77Mx7NcWZYevu0FsvoqeITxOcl0jUie6PK8py8ThHCx3qp1Gxjcb
nwkoKzLlVkoZKu/kCitUIJI30Gfro6lUTpYTBW+5zsrrOaCxiylmUl+q7siC7Sjv
Hjsbk+q8TVy0QBY5xnDIw9POt3ohXkr2fzstq0bYt+h1ou2ifjY35sfv3N2ro87X
zSSSMRXOl7C7EhzE21vELB28hQvp5hQVgjYNg42Iw3SrbjyLI3H8wTf3JywiEZtj
xhHbKoFJeAnbaYOQctlcmpO/dCsBjAhZtP6mK1G1jiCBIfZV+3Yc+fPkp5Vk4Yi0
XUslT3ZEaZmXFWjFKnP/ewwJOgC3jiiqvG6qpOWwUk11r+TD0E+cr/XkMbKTJ/FF
dB+mJNcwh1kT/e35naOQRKtT7SmDVAafZ8vjQQ8IELJentBcCjw3FExdHUToNmmt
56DGWZUioIVnLq6BHeMof8NvAjHV4JxVqrv7bB//msBbZ7JTAygowRht3AHOpB0T
XOUFDfGxLHrQG1VRQuCOglksJOqc01LM8ilbc+f5aI87FpP6pLK9FOo/w4AsPMn+
BUsqcHZ4OkTVeOqh0x4x8vZnEDDZHx+RXLihtH+ROXRijMugTHIivFtwJlgScg+5
biCuVZvMt+XhmGlmXgIz8ux9eHbF+F7YxG4oBcnAOZioQ1+nVdBSgswSasFE//AA
CKNWKfRCHJ9y4F5ow81PRUd7O0rwRrJqZB2Fo8eK/v0liZIO2k2Ki0g02waRBCLi
Ltwzb+kd43D2y47zDdCrD+PGYI5B6OPpQobx+saMAaPQ8bQvzK3rbJT2Mnvofy97
8rGq+TipXOGDW0gwRfSrZ2IVcCMyJSx4iv8FfobKI61sAehR/NWh6/ZqKhqeRAR3
ImPnGak0mN93bEeYgvaXLpuz1AptDuAzTK++VU3aoXb8WIQmr2e/CRXEWQQ7sDC+
Ift7zAeuqzgTMiNJZFit9RvoSjrXMsWbrONtfxAOK4HSKr+YaPMOQDRsWLdjjA4l
IF5lEwnKyBv/u5FH6p4wqYuWrAtPilMb32q4b8sWqJ87n7rfBgTSmZON5CmGBX5S
i3rYP//X1eqxwJo3nmVz4Z1vzrvpm4uCrraXaPgG74q35YfkavrvO3Zv5YdCewsj
iXMUyIuWI6QzOUGECHPh5NKHA/hpc7CiW+eVCF+pAkl3Hi6CK50+O9xOkK+rOdbo
JMCXWRpV+jn8A6XY7s1dYMdFlxHSumSqxG61oIPP8Jij8FFU20ylWDXIkfviRJ0T
HqP6TGAxvBsqhYVwBqdORSajIk2/rIsQfJSj/jK/rGjq4Lp6hxt0vCoOQNKAFJ9f
+2/2lW0Gkh3OWthR1pAxceVjY5Jez1KT9hXQDqDoMkA4jr0bhYtd8kyzodRzYfgP
mEV4/cEKqgcBlRMDD2SnlO3Z2mV6UEpHOuxJnaV0BS+AhNhFPthHNS4+PKL+jdnr
uq+lL+M9xjbJ/OAj1uE7clbLPohl6DFVCcfqyGUxzTETCWu21oDrh0wf1JJILIQj
o2cV1xtYotUyoQeTHpuQDjEcxwj2Zp7YwqeZgSEGcAp4f9Apg0NHPey8zBl8U7Ce
24ro/4aktF5Z4YAK9axFzgAdz075E6n8oS+1DctYrCI+EDjr5/IXL3UzRr5tLlrU
36cXDn1YE3sE2bgiEMuDciLntizRGXLfUUCv6ctZGoMhy3NybwUWiaK7CghQHUl8
8E8TfeU9KbJMy2p9x52MHAUnjCmA2upJMB3t5Et9SwQ/0wuPCQfSm/OT3c76tiMQ
E0yjTFCCp46zpRuc7hTd6cKc50vYXGVr1LpwI00h7rhwVZDFAKgeSLMEORyH+X2R
+YlzhU64MKv2RoXPvey/OcWAhI7z/XkEkqnFo9eHcyaJuziIfzyRJHozrvFpoW9A
5RMQuhs1C3tEornMK+H0RyUUY+LjjNRkVf+fsUAhwlkgAfxYp6LEdEYF1gqubbGv
jG0QU728C/PIfO7ysQvwagL3+Apps3PyvpS2eDI0DGBm0So0tAMBw8hSHtumUiQg
0t0GbNdnn3rUU4UOvbEpVqDs3e6g82xaUWhpQjL4nwdn2+rv5ncstZbJI76wSppv
P4A/d8I46fp8XpuzqeIOxm562yuLF/94/sWjDuyaKDrZRqXgAUkX2FbN31s8BaCn
DvOl8/hWUj8hguSdMXuIAMWNCXlCKk6UxSDVvLD/5dRoj/+s/A6KT8R5TE/eJ7It
JgUa0fDwQKMf+L9ugwz0Jlbnoit4xxCu/qwsbNNnyUK9YdPRaY/Rmc6WlPqv47Ro
JH0ueWv1qKbZ79sD3Na2Z+l2h4MdBM37D7DXSd5k2xp/U3WdieENip7jJ2G22lYS
h+frR7dtp+CHc29ww3m1LuQjRY6aFO8uaLDuNujCxNOZ0vcRlvI1G2zcfa2RnUsO
hlVKhcKjnyunZ0w1ZSg0m8cg5Upas5KFpP80ey7v6g4yTWLQ/eY0COUE8dxHy2nM
Jc5Bf9eKwE/IUylRFOVAQ0rG2AXU3abWZxkFkOSfkNzwpiNTxaaPud++Wx04LQOw
fXtlyXs59EgCtKAS18em2RZl9FRYwGO9dN6iFl9qYG8yPlVU1msgdcm9hBUbrUpo
n+sL93f7Dqn8rF5oib5iWZ7Prtpi5BI6bUqj+Q396cayegeDKIA59wgvYbnQaVc9
a2uz3KwNktk+ZndFMV0Ll7viPfV7yWWLDjTs4uO/ocXvXlIPr2jF35rhY1LATY8/
VNXQ5Ydsk5pANxs5aTGLGsePe3cufu9PrPcuGbL/+dLbmSn6+xmTA5hK/mCQu0V2
rw1dmoJvxkKLO6Z8rprTznH6WgydzChYnd9q77w2X4y3P1xsWLfJDjsrb/qO1v2j
MBfN8p1XaTSVb9PBPuLw2MJ88T1yy+I/NWIFoUpLLPoBf7j5yRYuap6xH+Vb5xLh
SaFWbwRoOQzF7ZK/GLha2/gjMYLgoUAjSbAmkp/xMcxfP7F4RE3iJErivf8sHLb3
w3vSCR76mnSk5ZYvA7pBPL6n9f0V3tk/lf3HNPey+jwHMSSO0VvqAiEiz9ouJX+0
UOClXI8kCZGvwWzPB4R/AniEtunuND0LXeTH3/WIoBeE9R/Q3/Tbdl/8sA6OUCA9
hSGaP4gTj407tMxqmzDHCF9XEOcRtanthsd/bk1eiLI=
`pragma protect end_protected
