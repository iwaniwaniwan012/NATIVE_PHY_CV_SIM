`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mcgS9BZ9Ea4uqsyVEwqkfsJTXQ6XjkqhWBN6q5k66YsNfYnbmguIapyWVlA30HcZ
rhHO/rTYKQ5mbezp+rYL8yg/XQDVpYh6dsi5d6wfVFVzLGWmlL0k7PzOWfa2PENd
lRbDZ554Me27+TY2IO4NevfqwphH29dsfsVq/8oN1s4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4096)
n+AbMmRULBXYkazGYpqujYZxFL/6eotltxw+W8dVfSmJT0MovQzVNptaQbSzzH5C
E++sHfrYOZjhrkSsZPZPGYJ7Ao8dcxsjtZiIvYmpZi1i8y8Grd6EyqpG63tKAC3L
N4hS2Co/MULrud6+10tHIiiLN0nULo02iG2mtphzgmHISAfXEPys36a41rBAuQNy
SNVTjdQwSZEleip2W+xCakBSj9pyexv3N1KYIIyREEJ/6nj2m0JUv8NIQa5WakR2
s+rDuxh3yonuGLkbIy/dRAdx9vp80LIutCaJMjaGKCJXaMSautGNdy6asxI7QLFs
zd4c8X8klqSRqHeLBblj2pNxjx0FtIaN8LIaEKdSPcf3oK1FHVG/0bV7mJRBo4DP
LYUnd5nQLxozV/HfT/6PLZqrAblUunWyWad+Ai7FkXxr92TG4vznovI/Vj/o8FTi
pXgeVBwXvJsuncUmL3b9vou/r83C+SUfSyA9SpF3VwITqWVmQFlI7eTePvQCQcfo
y/RtZP9t03U8fUi5K4saCNlr3cGEq4vFyI9SQMp7H6F+2vb07TsMki7JFf8G8GZE
d4dWp4XMxvDk0aGUjL3hCkkEW/JAy+jiTqBhLuDnhZcFG78XKshL8upWDWzMD4Xf
P7PekKavlLAgQo1RqOrx4y3wocVV8jlELHjH1iU7Fw27lwMcSyrFZ9P0e5kC9F5G
8KmV9FuIUprIyB3AQzNoJ/E/GcsAVr0R6d/B67BcTLgVG/QjV9YNmGXGJwHtzzNz
osKjpaoJNigbB+proVH4u7oTvJUx98QZxGsSSoSA8hfjuXwzt/GwiT2dRiHTksy+
q3k6f3mxxXA++HkS3IzfJosqbDGfPbFBlLrTytowXaIuK7hUhmKHstZAS5flUzDA
Hr1fwzB9nwJGWS/bhpFf7EoKYqXeLo5OqAMQmRVHdCKxvrd61hJm+2WArd1jlJKF
JX9mBX5uDRyITJtlEEE0ZA0MgpHaanjd5XqjHPnaVm6dO1bnfmIfm14yFeWJb7bX
VZ9j9rT54pNSLCAk9eq/N1IiHviaUYomx3rLbWudFx0oRosTy4spCT23iNk26kzB
uWOSVj+1XCJuPtrNyR6NkkzOmjpzwSOtdZrvvLsgVzUi+OufjiUPuByEEJ4PDLLD
/0rbHs+iN34YxEBX36iKt9fY9ty8AuLYLQZ5XzHh1pJUX2f3V79vU/l6SIoLputZ
LojBAUIuJAmNy3ZwDc8tm7aE3JpDtG7mqhK/xLlkIkg9+6qAGcxcPRSamnoQ2hV2
ebwU3R3cuc80vEoj3KkMpP8cJWfkYG4nyQyMZlzwG9WMcfBXLUNzQmaAsGl/eFsR
SzYeix4vcG9XPGberZX5MjqiztFWziVWElkcAGqPSOjigT5LgD5Qzcb6VCnl+OXb
s8JTBI6GujLaKjTKL2n/+zJHXLZ6mkMzwfUf7PD/uKENfKl4FxUv5tf+mMWCWMp7
czpEXLsWCPuUTOO4zsovOHmqqtdHBpi7EUKtpxQNR4ED6A94uX7yD2hcibET9Pzq
NvCnw8nRcmqJ/tqPcXl+EDkgBWKjiA6bHKevJcr0w/lkNTklsRsttjkqHbSxLtL0
v5hpWwrKrngOJ9WD7IKRIcWH6Ev9rftyLAO7+087Xh4N/pYR7IZsXpSVuzKAK/Pr
qoOAlgYR8E5+0omBy9vAEGQLj09fYV3ZMVZnW7YvEAtiAlDG724fUIbvBdxWReld
GJyh5zRvVr/9OaQQO3hyo/0va/jk3/iP4e4XobAKM/WBCrk0QQnxuuR2U3BKHXYN
sQR81r0BfmER61VCCGz6eKltqFNzdnRodeOW38/lgXUGvIXKDoFvHEvVNvRbKGq9
woRsCl/CY+vNT1j0wMs4AbTOdW+SaLjb+sexieFBzKH6Fg8kYtmaFj+PGW5Bcohc
uw2LhKddmGT9QQQmf5m9jrqat+iMTxO0TgJHpRMFqblMwVpm/6MUB3dVQg5hSycY
f/KceHLb0/AZrkr1x6+n8p71lYf6XG/KXSEAb3NSyx7ZnUNZVCz6CszZnvq2Tlf1
pCWOBMP3UTCCfc1JEQRVN5vr6/wPtSOyzgNr1HISkmVt18ig0ZqDSNYLg/pDLt/i
ekh1inkf7EG75f5lUUa7ZXLVgBdECKhiFWT0UVZ4otXmE/H5p514ZMl1AQa4dGpF
hNWEgyNWmDPZyqK2MnvCfFYYPneKN92sxysHfJ891WoA7SVMw4LvHYHLMx9kZNo9
cvLa7U4ti+OFLS/Pl2bFBGJ0RBDfy1HjBzO0gm8pyszr4klWRk4RCZlx3P/3A69V
VDEu8HwnoQDWkFeNJe4UDqdBv2L2YhyF46BCpnehBhy4FiBgt2X0hocF3g1CChSK
7/AGLy/oRmDplYHckxK7UmjtIazIBmyNRWNJS55JWvTeGGM4sWED9BpL8n2FQkyi
jupvCLnvy/24Eub8fAtyJWUFWGHlV2M9TPPYuHLbRq6xprHXF0FOux0uUlp2CY1m
FEUBR1JdQ4F/2LYP370V+768ADbXI1pWXlZo6PfzygalEQXGKAm7ASotwTnKX8OK
67PJmDg2fZ2FSQAuCeXZ1bwGZaWfuDjv1hOKLljwPGyBp1NFRiXeyWsJlBSlVwIl
pr5v/UYti8fuRefsLPy4eS8iEgGdhXErpm49/N1GLUbqtk+51H9Tih258pHJ4kLZ
jHOb/D/Q6nCzBCuVnIkZXSwnfjKyI6vlh4Xad3Plr+sRFcalD0WM1jLL2O/KHRF0
LXsuxBKKqcp4EIoieldbkNRA0crDWSRteD8oSmCKyg3ZczsnFMuwFGo9gKCAcN+r
Cb/IO6T1g60BgtYV4uCpfsOnHFw8UnKIu05lEqorQLC8M4/YfpYRZZPsDnLyNcN2
wZFLX4NawwqE9Drorp1LAY8A1KtBefsBKAC8cU8Y4uulSQrLwVPF5d2XJEE70bxe
ee0Y/3BCfTwUMZi+awChT3y89u4zUQ8MZBD2rRGMES87Swhmbhsoj/hZHXMtVs7d
nkc//h4kaPT95B0b1Fd3H3Jf72n/1nMCTphnFOvJXHMXdwew05mrcKUaGnCqYRFP
pgs8g3YUkv83SmLT0fEDkI+BvqzRCECRAEJjZP2y7pdE6U7nEJ7ujgJr/dD19vkY
su07cdW5Mtq34+UQQImTr9gwvQ5MgXNI4SvMuo5PnEwyZuKpWHdS2KNjl5txc9aO
n89+9jKC50vfQGpcPID2UNebDy5njJnPwe8B80OSh9sHtiC7aP9VECNGcRi+b5M6
+d8jREV/XmIwF6c9EEN9Pl9uXF8o1+/2kaPOK6cja2pVchbX0I05tKXcNyiZs5hF
hUUudznk+yG81iK1jBUSidqUfxfVUt69LDn+KRiK+fItOMYH2SFh3jvVx9Wd/URi
N+avWwvZLBuT06GMVr6owsH0VkoQQQypOUOKK/dZevcMIq83fKqlRLEbgHxO0S3t
FLNmZFCxZV7u2bzLyfdKgvQ2jcuNBnNFAqRtX+KXihnScMIR6rsb9wd7OgB7uW+e
l5p/HNFI/Un7HTCl4WOOnq11wtaW59zWsMkq5hSJTODrhndFGCSyqm1gt0LGO9ux
pXjASEQt/5i6Iu6h/KWb1BLYpiKs3cu6jBxxLJ8Lg4hSH6RHmx4YoisXFPItYdwK
Jkq+ImKKfT458MczKDzZTYg0k7/g1sm9zpinOTZt+sg1e9DeJ1EmAb/F6kKHJaHk
id8XHe3KZzAkl9NfLDXh2z4x3hDUZaE6W19AD2vFlAh5BDlDsHFKy+O0/u2uX8/L
IrhbywKJMLgc5ltq7YuhCP/o5cZYPv3tYWsfcV43zdx2DZAxRfPmZsCJcxNLPuCK
HgFtvyWzmYdjY/q+shBD9Rmd9Fsod0jLsPuoSSQYcDufn7gO5vknL1ZG2w3OK6pj
byazzuq1Z4C3DxGyWZ1wGCIf4pSHa8fcVAjrvoG8DiT5H5Eob4fsLA4Qy666bH4u
vTsvErnoDt872UVkn+pwOJLlJlGC00qQl9sa0Wd3uBTTti7x6GqCfH0UJ+whwOsp
gGgb1GvXGUDfBwMBaKOkd5F0u0IWY1BANBxc93t5yu/fdmzEv9xA0viwpzuW7zIa
jT+gLqGqd7S30iGY7dN7CXb4gl+gQvbJ+ZmgHQ5H/pno4ipHa7DKxK+qaKHVqHPC
qekUbG8L1qBDGyzPG4Rz3jjaf4XkJGjzUnIHuG5VaP3F9YJ6qb+QejuF6VdiwH2i
NZR3fknyYLdmVgXU2GBEygER5Dnic1rLboPRknJPyQ+ez9mmJrZo/sf33CGGF+QC
Pnux3Wt1HXOsQv9Df9i7Xc3ex6tVh07CBcdLtK5EHVoSd5ua6R7411RAJFh0jAJV
LUvvVGeMKyBdOPKVazvG34G1bQbZBN1QoA3N+v8qpR4cNuGU62qSs6OVTx4dGVlz
R36w2M2/D5o82e2MtaBF1MSl5HgRoC/2TX2boWSyS4676y1Hya3zm+nzo0MYil3X
NdSkY1Bm+gxKzk+od51l/f7G8+W7KXt2kCuOB+jliflcKRhO2RRp3ekmOHzHD/TT
BVuHmv43IipI0w2GbLe+6HXQ0t4U2VB/59izYjv0dVncirVzUTI1xKX7rxaL0wBk
ixZ9f6SfM0Iw+BuQkmzdlmeH+CT7IIyeSGVhg8K5fKNW7SFdL10R7cOUn9JZYfJM
OJu9Cy7EaxMlEJ5bSQwv+5COz4aR+dSnIM6RYMorl7QtZJfFxJM4VxIFZl4deLIR
OquUBRt/kWbFrWWgQn+9OtI9bh3N5SX4RiAl5hCnRVm1r2DulhHVcJfWRMTSC9ED
/36JJKNHZLZ51y0TFHrQxnpm3SsGxbnNJuNqXc6TW85SIwsFF77kMD+rFAQeeEWf
hEhbp7TaXAHYE7OwqEUZUNwBeqyEm8keLbBDdl+sMVOKtCyE6M/lXgKfu3vfzzzB
zo7jnh3W0qcSbd/jjrI5qZ75ldL5okaiThQDit+lOHjMb3FMbG9wf37UKq0wQSkv
YRKMVl4qX/cl1xM7/c6GnbsN7LgrI7UGfrSI2t4KAiqN2lPAX3hjl7FYRMK0jgO3
wrxWrLZQ5LoDV5gfzJWith3xSVqqtUe8bI8yCqG+7zAYfnGb46X+iSxLEKKfQtbA
lgvgWa5cF1Vmkc36Ch3rcFXOdZ5y7VsuMaBlxSQhuVPTDzHsbXjcvCJ76n4o+PJH
rWxSm8GcQAgNzEVg0QndnOxXrn/M8s1Z7+6v/r/0ChS/Z292wMjwgGI1gwRok5Yj
hdLDmYE8PJ7bZdN2pWmHBqrTef1kQaBaaO+mi/b7GVLWeArTOBr9Eb7yrMupjcEd
Kk2TEovYM6msx+CrjtfkSDn0/xFGZljuIf3D/V56vI9lsVWQRv6aIi2AumukNTPX
1ft6gcDjXCJbTa/Euo+5QlGTsGYU1b4jAldPLbGCsA6sG6KrqRViIh41r8RP4Ace
j81PPWkk/ZpoUlXn2jopvg==
`pragma protect end_protected
