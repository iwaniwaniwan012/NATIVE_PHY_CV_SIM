`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JLcMKR4A4/ogck3BGpohN5dI7lCySc1ytRzVYKCvqcuy2W6BOx70Kahxdfdc0DTL
CTwED7yQp7PYIuizusu1pHDMyxhKxmkP3BJjsD+WZ6jE4oKiktOlp4PHMo919PU6
lQxRGlorG0fzYjJFPvCe0Py8W/HYKYBzKx37//crrJ0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11376)
yC1v6l+ZSDJShSBO3kjdbDvSb85rdJzEv6bAWrHue1yRhsQJ1bE15gnkku02JiSG
WL61vfJNXksKOfzz8nKHQbVk4SjGUPIpac6hJKuUS5xbUQllDi+YuG/1P4ZcN5vN
h3qXH/aNiHre4E4E5d+dHIBX7CSa6z1WBb6SuQAJDCGa+Gj8Vqnm+F59zmk74WBT
rNXFQcYr0a8ZUSPuuE001quhxNmYDNv6grOqAXpNEZv4g0OB3S7hsN39qb/jSDD0
YKo15rJeCnNIHXCuO1XoZzrK+7O+NhW7fdxkz1i+GUCEtBWWQcBGUtqPcz58LbH5
+yQKun6lNCYoKJoisDjajhgMph3bTj//8Uw53gCPZM65YEVTUNDeykBdrFyMnXY2
0nR6XtXyK1yAjSp5MmzZ7DgnKhIW7ep6mOZuwn2qz+Kp42qDLmCnCsovb2ld9SuI
X9RtI8R5rWJ6K4b6qzBvJ2kILi6A/lSxH0sO5RQd9mbW5/vx8m7riMbthH5/UqTX
JVPToE7x72bkbwQknsaZ8uJYdIGANt3Y62SNpnp/WmL4yTMd/EL+C4+U4Ebh3d2h
w8DDPeLTn2JSHGbObhGj1a3/4mN3da1hKUKmGn5HfgkjWad28vfblpFcz4qmMQXW
kw0ZKN2j4b3BKPBIFg/fjSU2wJsqEY441FVsf18zyeLNftmRQdkevmOJJyFffsAU
ZIeg58hdVOA+/L3/lVvrrV/+qCHIn96Fx1F4SXy/J8bu44WAcSV96giF88X8kry4
Ha+SYLLPmgHhBleLCr2qc2TT6SGKXEcDujMh2BX69zSyjcFude2P6BxlihZkldeS
gfr0/k61NcsdHscehDv4nmf5zyQ5dr3qcBZYbf7R7sf5XBSoujD5Q0TgGuNETT6r
I0RV53iroNDSZlCHmVUQQ+GrSN9R/RDA2C/xh3W9QGPP3hEBFJqMv6gPC+DU3D/F
8Ag9NbaNDYP67JZo+Ne+l/MFIeBZHmAo+KJnzntenYrWgVh9Wvq3uTS0TmIDxuU3
8cczubOkN3z+xPhbAxhpSfwGm8Ssd9lLQttAzVSEZWzGWb3uXC7Scc1DNqTS8aac
L5vVNWMGdzS3kBzhzRljjMZFjblIjy6z1Ys8pV9D/vE57R1iZlyJv1mX1PcRMnb1
MZOTRgOYmmtKKIQ6sSgkjbVZhqbAxW2u/h2fJbTcSAQd/G3MxFT+tx3A4rikK0dq
b864HelgnJMKWfhMO69zT0wRm8YB3gxpRNxyoXMzCicO+3S06x3pjToAVfD0sGzV
M8kCi6hG3n6UP8Sj9ECwyeRzx6MTKc1YRvAojOZ2LECBa7HQKdcca5E+j/7DoRk5
LJ3tiPKlNvBIrbvHKrHMJwtEwt1ggEj6/TNm0VvJpdV8vqMSRh2MM6KaXGHk1VOf
lqmdFZWnys9KtpzXh02K4Zhl/co2GFXcAoaY+18v9I52ARrJ8bwkWKRuFBaj7SgD
0g7el+n8p6YBHTdnqGeQDcslhaOgDqdN9dlW/YIpFTqJWXO2z6heO+EOreVumNxL
Rs2HxSNMHCSyMS94qGneSUtAlG8xtkZwXrxjQr1rsyt3eS+NDhpa4ahLx1N0ZQc8
Zm8s2JFPjPX25/Hr1PbtRSPJVXNJJ2xjRqPc7P44kI8IPDh7R/M8CVtNQGwb0HPV
8x0MyGmUp108mG7oEaM/eQcw8L2ZuJs63THL56jNO8psaHWI4lU6Js90re/vQ/2q
wG/8vrApTkCT6rZc8x+ygLR+wl1wl8gkdRLH17mK1YOBOkSeREU6yX9BIrIQ16/C
oVTuQTYHXDmCyJTYqP2ImZvoT0iry2g29WKXUfnQuW4Xbl+bQSSuhoQKjTUuVFwm
fmZjbP3kFzSBR7HCMqBeuwgSuqUkF6aAMZa8mSwIDC3Flhm9lI2sizbFrexwn/p1
rYOMDGqAPy1EEcSsWyXkP63Pedv3MY7at/V03kiRGtgCsntxnTJwTKUKSeYs+XXm
xnldcvGEwSs2wRvk4q6gwK1tqtu9wPsil6CgkTQGEpl1jeqyrDu5QWiGXEsz8kiK
epmfqfldZEY9aEMOpNZdkG2BTnBG4VzeKHr965iuOGFI6954p18JuDwGsdBw/REZ
Qf34kPiBr9/7ohPNi5SJD+vcH73Y33j31HCwV3ibdqaSMaeFyTcMqqh0PHHbpy1K
RoxtQR1iMqzJwMJVTJgfnVc9cxkZDYKRC7+TPVdkQNaus25qLa/YF5XGjsVAI1xJ
XymMuq6AG50dAN4gB7wBzytNX0EkOCR4wdbdgJDj4IKye2sJUr9XO8fDB8nsMJSh
mJCPr/Fx4beAxn0Q/JpmXrXa9RsOGnY2nUDqa1tCmqMCHI8G1JzJkX2Yy/Kk3dwu
41wnqakBVDaomIX7Au2gIeJ2rDmrk3EbHMcEEk4oqFLswadONKSc/hAaHVU0jXi7
ZjvDXdkTwsUVGc74fD53CCYllYqZ73HmfRIsz7PSGMgrlJ8nog4MsPJEnGarhHm/
gU2ETbCYl7tStj9TCNmEH8brnlBV7KnGHbL0VfQGED/YtnoxH9xnEC9H0qh6/xE3
03e/UIO7fOBdtRARZOj9ysKB9k9f6Zpd/iOfst5QEVciX9Wx/bhO59dyip3x5eGF
Pcfoagxrp77i4Q0rJZ9AoVA1BRzWH+pymhImr+rdwu0Q9NjQhE0JnwgtHzPu4JjB
mC20zpl7mYEU/LnDzg4apqLhpPm73xfN1DmpPkP1CYl1TXH1PMfJAri1w6KzQJSp
UXu95odlIZXArWfb/f+CAWe7aduAbiuu4vbpr5kaSbG/EJC2bketg7zLzPAvz4EL
B7VXhbZjvCTP/8CFpizRXdL6QqD4Wi5aqQtciDBxIWD0oqVSCRAUUCqsTVHOBLU8
AClCxlAgDV0Zcz9QLPIzBNOtsg5Id2LpKQVEb+mfnChFe58QcZx6wvURFPYiFaZw
CVGilcUIT/HlfO4eFasJ36y0FUvMeXYVRNf5O/Zsk0pXMps7/XphTZshSscKK4/H
nrYxNI+Ch8s7DrN97hYypd0smN6Kc8yLqmA9rAumLCyUbmWTa6IQvPTTzN0QibZp
f6l08Ka3Cq91tSAvXkCa85kRCIR7DX5mJMaV+D/vtZBJR8f02bwgzua6Q2Jd/kPD
K5o06fKHrWHk9Dw90p+bS4Cw97kvncSgxWPbnXRAzldwkEtSeuvfZ6qV31X9osJL
QQ0YH6uLZ/nDZPHit92fvC/hfm7/HaZjRvqjKEU7OPl+L+wNJs7sE7rdedSCc35/
wEnNaI6zBYOcGwtsf1J/lZG8jC+/r3asSmYYV3klSWHY5rxJ2e1nnKXczmc/vqKZ
13rVj2mpOGaWcqw2/VcIDSZfZIpFkf+tA6V0+lAaO5zOGb+xZ7DtIkjt0o4qDF/p
N2kJ1wnV0iTJ7vp9XsSX8SO+MTdsgwnNCdIvAI8hqdg1nJodWdiPHkR6P9vTFRuF
q7xndodT/BKWCnbxr4YMnRe1u/cf6r4G5c+XQsIO1Musn25Nw4wbzGG9klOya30C
lmHlWWC/rAG/15q9l5iZ7CePIC96kY8AJLd/NJNMJN09v3yFZv/Kt8xidnAI60DB
1eieP8/GLUdRI/UgEoxgXfk0Nj+nbJdVSCmoUI4K+zwNzOKiuO+vhhE0edHYmsas
lQLRG4ErRTnKD8hDDtUUzOAn8yo2K5wgbC/hn07dXMRNSdHXwXk94CwwDBqzmh+m
wfeag8DCMVgtPoLtf1D3DjfMxSOhsSm9ltR+riPXXDh8IvJsPvE59MlYtP1zyEJU
eQ8c/MwlJkQIP1PvZSunTTOxqM4mocAcpNSE17IARFllOG1q42rTsiHN/HOSzkip
rWlU2usEfstrfLi0Cxj2jnGOV8ldFJdl5MTO4cUKh8rxMdT+NKNOZoD9PONE4kaE
AaUzT4Q/g3Tq5q02Fx/SZQc7ku/40NC+rEE8Jl0lFKZi//82aiPLuNROzHnKMSmH
GU9FKxQKfV4wFDeadjSUGFY406noWn+OPtrpmAnpRB7a8VUm/+XEgYd8a9JxL7BY
CHjK2yHjZw5+mrhD5j57TXDi8X2wI2fb29gNlDo+Aj8xKHvk5uJFANkQ/+uxT63T
YjIXTbP0wRUiiYaFyUf2V/I/VXKze1z4bQ4vQcKEVLtqYFNOzMlOFVWouatpCivN
atsLxaZSbKCSCHbwjOdxRvwolqc9srO//YsLP0mJF7ZE05iTDtOhUZ1rjSLM8xZW
waettfQF/t1/nh0KZavPGaCnnGX5Q1q7EoLx0aWgsXP2cQlG3eB5oayD3uXzWWDw
645BJrIgv4TLi/6otr3mgPZkrKmBzI3KDQ7YRd73C5ojYEKKQWsYCoPyu244OA9w
avQB4lHi8pxjDMypX+Dmw3tKs/e3ofgI4KUgz9GyYNigzAZlYmci2b7jJVR/PNYF
umSGM4nlqSmRwINrQZfbDaLE1H3DQQFUarQHQd8eejr2Bdq0+NYYv+Vw/ap8LbA6
RYNtfju35TCq79UIyQ5p5mNGl6NNggKvJYC1rTXr6odI7S+Mks+e+4lNkPoUVe9I
3AwpA1UB4/hiddOx6aJ2jeHZ8NcQpgHy9sFebbT9d/b8xq6VOvJBqeWY1uwaWlEg
2sPQy3umXGQCDneIIjCLUhNyLKtWCB4ho3UMpdPokdNq7yJ9YhAUUtoaCgT4N7V6
5Fa6RxIUs5doJbIfnG6GOOAsSWGmBCC1nR3+jgKg8ER+LwEAHVZOBE53MD6tEi9O
IPb2aMbASxhGMogdpD+hzqDdh6VC8AWcSh0XQAXkFykxMmbzz8HE7p7Kry1/I0X7
1tvoX6hh7W0qPvgr0AsKk2qIslyObiCI4zS4E77yBWRAeo8ktmZiQqDAYc8tAF1u
mr0U4OqxmQ30uCivhKjUjBMeInTDa1JGE0XcG4uzfh+qXV27ut4S6a6gAoLgASMK
7X+Q4leByYG1aJpPmeEYZwtCTKOKO89LyM5EcVwbGSJRbcNpGii1vl3vtRYcugoJ
brFWX1n/ngTSiIf8HT16CWmKSWO3/MrFx9TpaAkCUzRNfNcZD4KqtPpM1GDhQqnI
wvfsTi2e39o+/lwW2vWKCFhUpFktpnZKRUPISXCt7r667pXXw0JHX7Oo2XIUfSBX
jbc6cT6ZKgYIc7lM5QJckuRYphwLXvePFAJyHk1PQe3137yVN40okrOchPwOk1in
g3NXnTKAHWV7YwH16Y+4WtdCVK3wtx57PK0HLt2bBKC9yEgaKvDGGcc+HC54Wl8F
LM3Z2krOxb/fQaOZfZ4yVRSw/3YPPTzXOR7DWKzYykhKi0e0PGxdB0PXtXx3E4a4
8X8ynh4vjxsXgfFWzSjnWXw4elqyOH0zAaJFzWyecBFXLS+ZUXg3RNwaag7W9TPs
fb4r4L1/M4YT7HRsjPIhTXf2KlvwvEv/LhBn86KxUAZ61AfqFvddTP/uSTLxQXrf
TYQJzuG6OORet2IV1qDH6wyKmMFqvbSzCOu+ZDXBUMjqSsseF4Z5NH8Il8h6Ah+m
MQmexMHOW8G5h6vL7uVBZ0Roa1DsaglwzYmTaBRjd6X9pviq+xUBAKB9SgWn7ccW
ft9Hny9RLd5F6Uj6L3zeH/xSaFpCoYWfaMXTpvNhCXdtlalgTgSm5hVppjowlkNU
HAinb8+RWcVrShUrlzYacqxvTCpZ3j48Aju6PY7+zBLdfEqiRrCdguqedb1iuQzY
786ygiL8KkIFpwhm5zMWDYcUO3i/Zf1DGbXA6s4YXiYZQwrhs+hH8euKoGRZkNRO
IZWa2pa3uZFUZbWVeyQLTxxfoq1i9uwvvVUnu0DQJgyF1hid1aKkUfkIieNBGsTl
axssPhj8vRH4KeGUpuvU5mNEPkYFYwuwbhmspv/VtA6A9UYl5DH3PgmmeoAldsGA
9XxJBUIeoUjgykS2rAMIuBr5FY3VQ+SdCTtpoD0/fzddecU8TZbDqKYpkwq7STuO
2GzokDL0Gp7EyVj565qTfyA8jTCG/2qa9xGPxy8u0e22DU8Q31Mu4Q77cx9fCezm
N3wuXzO5vDXW4dy9dofF93fsKRbq315oZJnpiKiJKzcRgwvahWoDaGteDUBL1YG0
Jifdzpl3kS1h5oPM7k1sio64gb+YHv2PdQA3Q1/dy5/ryU6tdUCEDzY55p67SVz3
YGrzEcvls4ZJoBIhEe6ipwUChmPHM4O0oCWeAEZTGWCOn+N16k43Hrbrqyx1H08h
svV9/f55oJDlsahOu4pLrfun7C64EYHzEI8VBLYny2qMEUBuIJp5iPhJmcOgzJWe
ntWickz3h5flzSqHWqqM9QXghjbo73pHToxbSPVfyLOSqc/gOZyGhhcEh6eY3AzH
h1AiagZPcAirKP8bK6zDHevHQJPHARJctbVKnBQRyt83DFkbEt9tHm2/Ps1m+iEs
zz6ktTB9HcPugK0XVSxVjVnS4D9JCJrvpPpmVbit9dAq97JM8RmtOUfG2zTfesCx
3ln5OcD/s7v6PJIYw78KjSDWkWVxsgTvgvaF/AKkA0OZb6iErRbHEp61r6dKar2K
If8wpmhGECDJ4p7L4yVziWMt/FjMw3EJ2dgFeIboNTviJ1RiVNEgaRzHhX5KBlT/
n+KXtYHX5YZvjB/vR3Rnb6hFshudQ311ztyAdPBDs4Y7LDu8RNWZOtRszH0KFLne
nIHMf9O2HY9Rla0GBZT+aLJyes0uSd72qv3wV/wk9SgAI5XQaTJI2ypgI6/ay98K
tlggqmKfs6TAU5AlKQlig7H1bqKphofCbrM2J/nhLT1nhfpN2IMAXZ8G/fhuuptm
teY5Jr0RWCp8G65F/n1v+gl8xilFQ1qr5pVCA0gVWTPPVcmynevZ4g37+8FqNju9
CWxKzeumKixpS3z/tyZRUAmG7Mld5WQ4qgdBmy+TzCouNzYKp0XkasJ9WzdfDX+o
SpquLWC7fpSu7sg4uKhRLCIQcquyLy0hBD0uGoWrPqvZvo23bRLqJInjKcK8WmyB
TShZ8gq5Rwlizl0iCzJj7W77K+hSQjyl7/7+1s+X24Oa1HEIZD1ZFnATcgttKjIH
r1KzjYu6lpyNepH7KzrcQzHI2z5oAmYiiQ2S/LgKonL+2INbp+6juTHRzIab/Ys4
G2HTRcaZ8QfJoUtbuxkwKOwrsp2uaGQD4bg8k/ruPlHIJxzR0Eglyj9IabxfyKGX
LlqSAMwGrG/aGo1dlvep9fP80InwRIOB8TyRGojvoKd7AD/t3BXKnAskAXYVyRL/
vEOb4kHhaygimn9uL9pLltis3oozcu8jLs9JRbzUjmRikDPM7b0fxICeu9hMpb2D
LGVP4KFBEVn29igcfJGWKJfMr6aHduapPcLNLUI2/JS7lmZ7wGiIO6fiTmoJi1aN
j3ZM/T992PUqj3gy7RZ7kUjkByiVeCTNWDnBgQvBjC7qkPq0FXMsF9kHBu0+X6sp
QkwvWQGeVqdIoBT9fVuaeXBmp/SRv2NmUuucksgAA3DOt+F5gtu6GO2e/xJYpG+A
9LR514BCdLBWTOW9vY0xcxPl2zu1RYxot4mDh+WF/hNA3Apn5Bx6T2LMCsQreLR+
oRXSQMbs4dIZEy6wW3lygTld2VMesZAADkRoBg5Mym3sj4gYSwmRy/PEzIIO0dOV
0xyk1z0jBZQQCmv83DhKoSwTcWPEUoUSaPtItVVjg1lwx/GiV2eGplHLZhPLFYzk
91f74ai2lVE1/kSKihPYcTWbHtG6LKaeT6T/Y2EOlGzovAYbZqi5gJIwhL6BK9an
ED3w2DpyOdcvvykbc34ESmLIaXHIpckxlvSEixh/6KK4QupAKfl1oj8C6wHCoh64
oMyqphYyF5dUd44JpK6sDkhOUpYTegZay1hMIXHhzkuWjFx3qaH6yyZVA+8uDm9P
vMDfVx48YfMkyZT1Fhvq+eKxSIspnX/2kJyzgZsfVdvq2j+fi902+nqVwpfS1eiL
u8h7sJ+qTkPMhFprvR+8K3N9384CROcW4oO+v+Eb7bhxtDwMB4tP87quOblYF7Hf
RYb58cty6yVMwioqBsz9Uu3rMOydVA4oGhQvGFq1VD47LdDqM2OlyaIItxdMIOJP
NsL/o3LGiyZ20ExkKs4JW2dFtJqUg5/rOHKEstIhbdNw+xReg5zOfBsEK2j47Bh3
4vTEQwhhdoVXXsKlUqmqPD2t6lPV6dQKfN1potQ7SMe4otW9v7VBpCifynw0TKPb
HQOmgOV03AWhJPJmYxMfShbGZWY9CL6VR1k53v5pvbwN/G7K13PBqTbr+IVjT0WE
+1c0y2gghGEWKnvsA7gjbRSH5xuxPTxtREA7EpHNKzeFLBRJ100yoBTUpGJzC7O2
+hrnsrYlAdXcI3Ea0gsGD0H7mMN4PvwUyeE0HAVxo5N9R1iphNJf40X+YWU+xjg3
1v6RNHxJu56UYZCeNIufxQu9D5ilwAxm+Sos9zHugofXSV9oNDai/R6gKn1z+Sj0
ks8MSnSng1z4jNm4A7nLwXH9+W+CqjMrmLgbnJX4v1lQwYbI3HZszD7rreG7LQ+E
a869lGum3OUoh9SFHN4oNXLKg2Qx1y/RGaCLhjURiwf5qa5euBCQ3HUanFV4/cgD
sY7G3WbVEHRF7fuDcZFOih7I31znHywDOc3VSzh9bpKO+yn37ScKv4Y7Pgj23KIr
TSXGGbp5F8TXw3Gohv8S9P3LvHbdmYGmg6I3nOsxwUmFPmMeePlu0uqUzErRJXuz
GFpJwygCaVi7aHiEIaZAHGf6B4UxcTy5M5rPsdaBaIcWKQEwRzRwpNQZVeP1iaef
uv6fsnFWM+HjCnt5248Ri+RVMzorQ8P8ejSsbv5iROTPqlIB09I3LVsfb/b9N/Lh
J5fO6MIejrRNGfsu35tnNmzUqQ1WDQvnMhm4nhh4B2jEiJcvzawj6coagve6Dpgg
1RvLcT9fCUVXRnvveZ8Rs6sFT2J9NbnzXEOyAn74xd8BI9qTDudgwY6+m6+xqsaM
hFhDxsLL38hFfP8e3G7fJbnfQ1hfqLp/HZGVtZx6IOGR8sOR7SsHv8NLTu9OVuFU
ikEgJqWKqKRjP+fKZtg/V9ZPzIhy9a48P93HOTs8Lw1htRNO8kMnTayWIJ0R4HwO
YabaWN/AOci2AEGJFlGy0RHPKXXdzrRHLVCXemUZ0EMi2jKEwkL3Vxh2LwAfE88E
9gInMhV3fZos1O5be+Q/6fLoiYKAsVuNsD2UVS6z+msASkix/qO4r/imn82/d1ER
tYZtoYrWUV/3JI8JtJl0luEWw00Ln72hLEZHAoFjmLipkcfxaOLN4S+qedx7ZxBN
JXZtEoLY/DIaa7eAGqltsswC9hmrFzz8R+dT1lCkhE70Wm9kmZhCI6Xemp5yClYu
LGC40a3EIbZDNpH284z7zj1sy5qUIhFwK8lx/Ui/+RUDuXPF6an0oehC/RlrwCaz
/wBXLCaxREsiVun4qMvFfeWKFVJkKRJJG15WvGrcEkUXaaSXLlHavlPHmacdjRVU
cQThmk6HkmlbM3jXVPZe+7fYFz6I5e4RXSZkis/N1+KpGr240HxkMAZzmB3ZAFEZ
ZeHKsyfzmIYBG+wOEpkuks2egN6/FdeFhB/lq4xlnh23P9Z+cj97WhXxYVGgeiRL
dv2fFR+vhvaxBdAPNUULh0PA4Afmkx5G2bPgM6on5Puqan1cE8iB1iVzLODithrM
P2CQJwdTaScCOs9ZPtbQCX+2H1iLnw3ZdeYP2o/6J1xK37PmCysLX0D4rKGF76A7
Ho25+Zd6zzQN5r5qRX/dPh/0OPpRCZ3qp2zTW+2oi4XufmubhfoUjLd/qK4K0QYK
Svf+V9Y+TcHsDgXBWyiUDRU5tLwErJB3mvlU0Bdcxhk9g4iZDo7kBEnu6+F9IV2Q
ngh1BVWf6WEl0+m6AfGgeseK1hl1nI4rWlvwNe7Qztrbk1s/yJjKlO0JAH2VMJoA
IyZXMyflsjfeqDkzHiYKKZzTi1lC+VHa5BBl21XbBg9g49G87Vh8mX2fGPhreKpL
ByWCTU/Ub7CvXwpFauZIM6ot1CZkN9wM+fCE3M/n++6MWBkQG6kG3M00BtRF0Q2Z
0Gdh+wj4E44v40IPpf9sVtvmZhtlQlwpPaCWCn2F3XFo2ayKaUee+pEvQWiM4mxq
LZCyLuxjBWFSBzPJP7WWtfLMyczdxdMwYHJTi4/SMg/GQPJ/pspAC1zQghnwqHtL
kDqQkNxMGySQCKsqLF3sFAjjrhJNsvxyj6qY8NK7X3nqCUlK2d8YT3jXEXxNCVN1
LnhEvpzCFvz4rBL1KJ3FUFVja/yVXtkXEHvaiFYwaJL1D5nAac8hcMTTFGJsZVst
e9BbeBzxI0dRU8YUqEwf1y3JAFo6iTF6WS3mhgWtj891sYyULna2MpPkP0YtkgFg
my7KXnSWVHHL37h5Ccei9nSrWYcycfUkvPgtXKL9CBx98oMLVn04TfwS3wc+iJ0/
loP7SvXII4hfu9wMEkmiuHjdymp3hHXUbUSzVGeZ7TSmNM9aWNDsPVRujrVhcd+V
BY7JbWB6tRsnbAiTIknHQoNPRyq/5fgtqx9xaOP6bcpOgmbIwfuqykHt2xJBFoHl
M6MgpYWYytq+i4mjh74HwREWlf7v13yk5voe7HlwgfuzhBJHb06vSt1x2qs4idaq
AeW0LhbGocWI9ZQyhiaJGvJoy13mTv7zIMxIU6zVC/RCf0xQqFXIiOBwYWNX+Awf
nRy8YQIhsvJnLsPZR5THDvqlYHeFSaENmC8CkxnxRWCj2cltDzxvniEA42msreg+
Jar4zp9D5meVORShK/y0PJ7yBsli8SWn6FZL1SJ+LAmTqa0ec+lKEGmK3lnBRsyT
7Qjq5gJWI/RjocZ0AwfkIGlN0AiXa2IuTlj45+56jU/HnIZyz1C7ftRSRG6BHtEm
2NXvAT751DnlxMnNb+83kLKBzBYIARyJR1rWrBKqXkF54zQDLSyfTKwMKmJ4bigX
5JWZxRnbSBsdd/EremUj0DIVGtfAP0VolVliOf0IFxadpU0td6url+3zMWn20eDT
3SSD77sLUyb6NFcSUz08U/KA0FEF1w6OrlWnA7VnwuwEDp7pmRx4QaQ0rYXivYlE
IfefaJJh94IO2A2r66/hcyRhhOODwqvgnuRcl4wJzMoRx4G6lL25jGoCW/qkYE8p
hj6ULz1jBONDfUti1qAE3Skuwe/iX8LuYjLtEpKhaol21MRs0Bww3ruN47CUnrJf
VMEtUoxBQwg6s1FKHY2tCepk4hG1TDPlhX+3AcYpOB856O5d+oz+yQRsRc7QcBeP
EmwlTIo8baxZnRlEhxxwXgys40L5/R2diiK/Bt+ToteK1B79WPWHZZlA2OB6/fDk
OrtvpZ4OOXLB6X5ZBIpBDkeKem1gDIoOeLCioRGZxzPlk2huLJzKobWTfBoiJ1Xi
8xSSoDRLMH9YZJrFEg7FbTWGX4ibBuN8l4p5ENKzGGxDrjomMDU18WXHASaAje0p
4zAxXf5/760Pox8FiyzNqFG42bSsd2Vbksp2Y/ZzyoMEaQDCR1h7llKP9hDxWY6G
TG18TpfP0MCAD3KwzVZeqspLQTylz2aV7EUhRikeM4kNCgc8tpyfnEkMR4GTF3I6
cVvJ9RcLqm6eJKWfsitrdkxLMeDVWqixDGgnWJdLl7/tXUZqTjouncW1UU3EUFwo
kH/cEh9sXRiTPNYwfF3KqM8lSDzM3VMNChy2EjnIRJO5u9GMC+37o7DbSWv8ITHi
6DZjSlZcm296Y37vPpRnNpb29AIAQtniZUoMa2eQRM4NxbjQ+PUZo0DK4KQ2t1gP
sbBYZWlfUgZf/5VfvrTCo+mIYPOwqLVIpKyhHDjlma2VoufceEuU5UHEgwSRr+8J
ePpokutKYC94jdrph2F1Kap6JKORcea5JL5IWRDOnyXZmh9JlEo4by5EEysus3nc
zcnUrvCK2aB4Fo1XtYTd2bOYdDgiNJh3OAwhwF8DBlaX08mrqzuBESV7pg74NqGl
1oEdOD4eQKbiAeulr8SibtyVJBJj4zM4B3V7OcdhTD2tt0etqbBKpyYbjZYd74Qd
OL4VN8be3WGSVzLgypZ69dqTJnOMBjtvShmsR9W/HAAXx/LH3tDN7gOljCf7+k72
rQCG2aJuOmG1Z2Sil+FKXEFKYArfi403Ec+cLkfzvLZXW1BYMjiv+7OjDS8CkwxQ
5E4YwUNPN1ZZJ2KohLLdgRTLdmElisnm8S/BUdoZTt8QFIq7LD2k08kcsWWFXd8b
3zVLfd4qoUu9BvFRWtjJ0xZyNaFLt2R76ruJavu7AUeeuTs59HJhSGtMpwbTrSj1
ojevfgmszdEwgZJyCdm0ZL+PWcqnNOrOd9aYl1TCvqA1lsTrAEwRXU98dVUQ1zJX
bRTUqEjIAAQRiPuTHE9FiVv98IiEbGiw/6pTxLfNEYLK5awvA7BxcunZOJWVtQjw
czsCy8xQC63JZq+QMEXRlqqWHCHX/h1ws52qd+xFHD/SJMmwmvX5Y/Yf4HBnJLAH
Qi2fE6yJ83RxSstt2tHNsism4QzqwnstxBlzIv3lvcL9P5R3XHOCMdg0abJfB4uq
3w7k4io8MuKijmK4ItzJyz4QTQs6tUi8QRGoFNh5LTWOWEvMHFJi8S6XgYg3bY/V
qi6b7FwY+AcZgjhTkPJ3Fj4wVJqGbyBVCsGkvVwmTOvTnsKg87aYCYrhxzyFtx7y
sxvdeb97PYUZTPDLqBZGOZ80fwOtcYzY2J2Z7gqLiEs+/K8gZi4Ao9IltIJL/q9O
NktqfkPpYMvhYKHQreeEBPnn4bDDIYUb8aYGWZtKpVd/udw2LfWn+FhO8UOsr2FI
XN+2V6sx4BGrRPNVl8lvqRvD7TSyNykPnWznW42RauEaKN+et6VPpbfj7Ijn2LCK
hm2YViO7EEv0qpXoltNxzHbP5ALY22KIwljtWXoNuQ/KeaE7Dj68ZE/H/fvP+nbO
oHtbnOPYW77XfaH0oIyyJoulDLrAikYyIfArRGbqc5ZnmvHq7pNdWJ5araUIzIpw
mH/+xJqi1ysQB5s7wKC15fynwqc9O2Ww7iXXsenRneIK3nEyYTVqReY6hbzdB7gU
cIIPvaNdcUuQd4HxHx29S0iSvgKaq8pV2w6d2EAU9O1/BREl31mwODDM/79N1lGl
LL4GphMD96uU9QK3r9uvK/FieSJn1+ufuGgJvAtCpl85h7/iZm5/MZagpnMI31Dq
hgu5SlTyBHnuOQpHDIWWoJQ0MV48y0w2lxjUOx+B+szRrVtWkH3UyLJ+NFvGzKPy
jxkWB+pdkjKVfN3wf4kPqlmQpHer7iBQf9zHwE3PevC2/8zjwrSzQQzYize/cO1h
GYsd6gNDixm46e/hRReKfdAhTpKkoKNXHh8oatJ6Ed4RsODs907NL0BoXjMS2fP9
pzTptq7aiveF+JoM3mUfjAsRldtdiGYqu2aYiFMZn/owWW632YUc8FuyuWBqCYn9
XYEwqE0PkDpZg/yU8yRrAp8VKgHOlVnRhm0bVI+CknDTPaga1vggN7pRk44Ur3o1
s6PinMbtxfMBqyMIt5pM/v41Ey/Qh+/SVj9CthJcqAH8vD5e1M8JNHyzr1IeOL3i
y9Lj/cfJhdtbyRZhWnL6J3DrzZQEm3iaYLBJuD1ugdpmXYoerPssSBiwsZWstwP7
wq8bXeVStzBFPCDxnekF8KySV/6gpZPMmIxj0PMpYk00pwz2b6wx4hwyhUJvtwQF
4W1QT7pqI0pJSB9cC3Y5ELfo1nKaBEfHC6Jro9HSSSMNvvY4cFmtl7CyRIx/MKmo
MtCCJS+ljT0Oi4Bu29geLUM+D6vjflrWF92a8fc5y5SVKYvg+wJhUxN98zzzi8Xx
hJMnoqy1cSpv4U+6XiCn/xJGASCtyxjmqMyN2v8iYXQJq2rZACn3t926MrlyywKP
eNIugOuquTIf1P5w3Tl4T0vftqN6xsW+C0CGMjVwap2LQFdQ5sAxAYP0Aru94GmZ
dmPvM4XYY+sfrDrjQ24VTh0/cjaTiGTiKPTaNoX3G1Mz61fSk+nhhqW8/nvkH1rm
s+WbvK30UNqkedRFvYcCQkW9YPWgGEmuQaEvIGsefA9hJUPF2jfTU909CZ7Qtrk9
0frqXD6cIQBPbQuymHBpknXEUAF/pG6wfcT4TfrF1c7efm9RpqZ63VR6ZQ9HL90D
sIGNl01OHBcMjaeoH9XN9niNRaBI4G+cZGMFKo01S3faSAFmTMUIlRfKe310B78r
Ub7Lhd8dBg38qaSen/Ge9iaeg+GiqJKIYytkpSlIgdHh2/OPnlTaSW+TVbNs4/75
x+YI/QC1Ds2OCr1OtNGgLgiYD1iSQNVds1p4REh6CQDZDg7/NlXZ3Tb3bjcnNwk+
GILwd4++ulqXIgW+O4adShYrWyeVALI9h2rDETlAR3+eR7gyuXRjqLM3VIN/yQbs
wbwda05wO7QPcVkXGy4FzpYWp4AATZjFoM1ucKbpkeeMxqyzXlRJtZa79cLObc/s
bIUllQJVW2aKNYgBkCqoZnDjIDpFrS4q4TmFFWs+NXk46PY99O4TaHyOETPREhTi
lJvYEVvmeKKC4Y7H3a9EUZECaJG/O85osECQHE7SMdvXKA12EGoJyWjfMBOBapsz
a6zBY78q7AewSp/So6nytxVow28wsWfRD9L0f612qb2u4mimW873WmoQsBAkJgqH
3GH+zJtaj8wpZcXiTAuDO31QrTJvf1L+HO9nGajhoPDANuhXi0c6c9oGIXa4KBTm
DVynOqkXAvM6FcoMmmZRKOK1m1XTeDVaPH94j+JMn1zUpbjqcy+gykU+8Ba/vq1U
HFqv3On4Piu5a7PjgJFIg8S6O3iqnANEBPrF9dFbi0yPYDF6v51i6o+ZO6CE5A5u
QhWX1DTOuhtDFXNNrgJSrqu53OwoSyyHXmN6qeH1NGourvYRbHvm15T7jyXY837J
deoGtwrO+aQMtJFXvSjtME6nJL+QWb6HwluN4L71rbZpGhaYRTBKKaq0ffCuYezf
RFu7i7A39DY7rVZUoX6VAv3kWDjuep0wwbBYtJy3JSokZCImYZv5Lj/Y2iyJaKA8
l3SonYtNVwnl9GjPhQYUCBPMzt0Pg+9NE3minI+S2lm24I5rvRUPPH8boRt5v8Dq
JMKaIzHQ7kfbZG+jbazhua47BDrmnMo+SVUlRiA/U69OD9iEqWIkDHqyNnytqKre
`pragma protect end_protected
