`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BNetlG0AJjW1MtlDYcnRn2QCE3T3ApfXQLGtU4SOexFslwkqVy8VozDcNQCik+ob
dbtn/9PsJYgo0fxHCf+5vGJFymIHgM9cJ5NMJ7acLz+8ekEbFLNTxIxmLbtHUdsZ
AAB5FB+9k8ebgL5VFddBSjArlDykhLMcnd2BjCc2Cgw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24992)
msUH0RyMDquQwvnH4UYVWI/ssH/t15jUQnqaUD8vK3AgMmCth6bTMbr61jQyYSAh
AFVO8/Ji9oV5CsUdqwkXged6H8nkJCJZ+8z5ZDKmg7rALatdCXnx4FkkvAnvc99C
98b2E4aJAcqTDkx06FvUqBGVzsuIPlLRRaWzq+OTdl3owEhbWEV0DorswrQSj8/9
/ws2IuMxOg+KnnyS77HspSa7+RYVuohey0rm8eWkrx/k4BExJY4ZLtDCJu/XBkAp
8ZSI5TZWX6WQQXR3qZoIRHEK94o/8qxEuBPqeeuUvqQb6o8V/Es2dFzizr331+cT
hdwVijMZhVRN5ygVmLOHXRteHUh1/ZitcqplADyNsoq/dc7UmdVufjXWoXnyA6NK
tigPxXlb2kCwNE181NvRlThr91r6GvuhkZWqYdBHm6auCqySf9ElhaAlizm68K99
3rWOPBFyfxL77WGcAEXHzvze3UhVY2Uro0HvLfFdC4oVlVa6Vx7xlS7Hwf8XnTxo
l7fyBv7phCugOb80xs/Qfqw+zL9GiTTXz9hciGoPmlC1D/rVM1Fs/1GMNgjNe2h5
nlrg3TluIc/L+PG53NawxWnGmnVs2n8vIz4V+0s+2n/7fekeGTfpm8Ahg7D/8zv9
JWUzEk9V3NqOsG0sz105thHEn+vDHSdsC4Ab7y2mTNInFfrLEntoVjoSA2DSOvfO
S3o6kQBPj3C2MYLZ4eYqxrty8UNscdSxUYwfLsIFCYJTuSToacl+/LHZLpy06mHN
kmcAUcm9xpL/0JhP3juZl4ASAq0LY0u4ibmOEkVr7qJngqbjqK5cMKUaJwY8mk2z
EUD6JhiYA21drD1E+vmN8sBDQ0FF8zMJH7n1GFgSY32RTB6jpZZxXcLSTWwEmEaA
TAQK/QF+0u5oZjwFV4YaEoEp8JXIqEs24MEutdmQNUD1iReAZZ4r1HqGnH7Z6c0U
MsMzDnSDMwBh3jNZyPaYXT4GHSyG0w33Ec4zTQRNinpgua2ZxZQ5o0SwvROHHEcP
xQnQgXgjSCuM+1Ur0Ge/UUIVLV6sRBvULI9om4ioVBcyWEfK+zuGf4jU3DVPkJ5x
Lay5Eg5A4Tc0Mxjii3rd6kN27GhSiIVCLum/IuEGHoe+pfYTeo5Knh4Duya8LeYt
h1PRNm789j5QGRToEJoS6m0Xfg2nBeou3IjYx3W8K8D4xkshGmTjIt1fciaUq2MS
Wtjnogu8O0itA5baCa1j4uQJeDhMPJ0ShSjQHrSrk65L0LdB/DoJ/Ktj07SsiVpW
zz/q+M6hW+IOxCcukxCRiGxqqBFq2rrpsyVtP9z2tYv9w+HjZcfN69K4npA0Wa0F
bJL00Joiy7XhAliUKHkNLrffoCNPNCJYynnI/KmRlkFdUKcv5ObB29utDiU2aMxp
es9YQm17pGYtSilug1pEWiVAvPrtmL/H5GQUV2RBrTr/lV4Kuxhg25d6z4IfkhUE
j9s3a66t4XNZTNYLs83VjGZ5A36Y2uXOfAgEeMjy0CTITcSNX+D2DL6x0E7sTboc
pgSjUbkTn5ejy/ZHXmkjSyIwwIIHo9GMEJEUyFEXd09m2G9mFg2cgAiwjXG1QVWn
dx8iSuo0sU2R2MgP+yohvrRAws8zFd4WnGcF5mf2+saHKWd2OWcfxWNYjtZYm649
vAAgddIffJK5y0KkPAfPL+NMMuVonzHwuhqIfCW31AMvUCglVq8CUT9bmzCp/Mcj
E+Sl4x7IULcmcAfoaIp+jCHCO+dn0hrPzWf+0fUksmmppwmClrWL1oTDZRgCui9D
KCoPBd3bTDWr/0LLzFydiyFlTNBcMnVScpLjdPyoj2XslCLdgcfLFsrM9C8DAMUr
SLu2oXdA0GTrPW9M+lo9y/YJFPiFAgsBOeu+dPTcfc0c84iSn3+qFzb9jQI/Ad4J
ar4/PL7AWt7vFYD1ExrjmfPa4YW37RMbhA7dUCbYZe/taRVbnfWw6TdREs2G/I93
MpCSPLNFpnPl2w+1d8L+KqI0kuARCzdRmv3yCQQpJFBvScV4ZyhPLnQirpdcQxlU
xRHYBFpK60r/I67yZmBxq4zGIq3+wUbIjz6bFjAIAuNBmD7+3xfGZlxI8QugpSyu
vOozm9eu4qQZRN526oVRHaZPXj9Xewbf68PWWY4ueysEXh33ajfNJt/YG8VkYoZ1
tOul2MaOsgHvjtt2+RxIj12LQb9HqyltNzfH3fnPTlfO1Z9P/a9LlXkygWrKjeZn
xhGZdLE9MGf0F6FBQJd9dtK3O8y4Apb9Rhv5Z3haoEdVxB6kDNk+uCFuMDIBSuMv
0bc1tpKjLjysz1gfPJcDb559UzagWTvS8Ldn3XRdWb2GScYNX9CfSvM2YVUmT0AB
v9qlAVcoK0fQ3QZVqOskhtnjGkHz2UhjbIwMNp9WktAuARwGxSPvL/p2u5ZBRsvI
PmSOHH9o+PseJRkzivR8JOTC5bYOIu7zIDeqyKQNGuSwHnaAoAKqskDClY41hPDr
cEJFIaj7oTIh9rnWizp9rYe0mbRovJyjiLg1eoGTs7P572H5AK8CJl+NL9kEeNcN
YfOXtiOd0KkKP8TDhpQlOX0z9deKLFnoRvv33LhMHiGqSuhnW3QzfPJ0Dw1g+OhT
SeFfFpNBBSDTQakM5qMNe8q1KGVXWBCyVLL9U+lSzRGrkmUgBPkMHLrgEWCnuUyr
6y7nF/X21WSzW4adByTI7AfdcMnyJ+hcaJNCnxqervPowTkROwNkcsathJvR1I4I
++WRxL8ERx/2fxqtfY5Bbb+k50pGOHi+5NYI7yMZyJ+K7Mav/0xofz+2ScvsX4X/
zzMyYerZW04SEdZs+XSIIHl0M71t7tfJX+fuWXi2WDFMcId2hAmfzLF2dV3WnZvc
93DGvE+EtW4D93LyiaY9aAj1QGu334WrHMmav767DyEOrE6xQ68DfTSow1/i/rc7
4gEcgmVOUqmzX8tZfdJWpyH1A7VgajRf/X+G+HxcuW9A+UhWJou6PfkTM5jQA8nb
5cGdmMwR/zryZ96o0QEXLYhfwcA2uRjKe6YnOm3S3Y+9cJl3f56akeH0mjCYNq2x
rrd7c5FCw2MbNAzx1We/VkQzZIMUpgJWktuqmtIcc8w1c9VprvI8mtElxCqrOp4i
y1vRAohLwOOt2FkhRio8bGnE/fGMpjLhTJhrmlt7+PPe3faCTKG8dW6HmDKYTOiv
Do+MKw4gyNbZymifWCNor54b+dh5CHPzAfw+FPXuDCoeL146Ku+ugv6xgQicysCp
mFfhil80Ous099G09HziMjGlhKfl0zPXGL/Yt84fUi3nB9WgIMekR2rxuNFD2ieO
dUUJoew3OnStn/2jYd+evqLltEZNP+qxBpycoS00kjykhc32UWyYPHAbQyfE/ZwM
AOFDIQSvL6+eZEyHZmAN4QyQQu+NGdEv1eDW20joYCywWJCgLI5qSCHwnkjSLsyj
mTBUcs19YfthU6he6/ldXEakvMN2Mpsg2Le/dzW1DsT/5DkM7aqP4O085a+FDpcz
AsdX6/poi/Cz704UVIXvoauBRgPfK9Ihi3F4MbwleujGUjyYgHoXFju6tVvwhADn
8QBDkBrsVTgplxSwzpZQsG4tKy4NglGWgid5iuFUnL55oix+1hu4SJceDIpp0mSf
LMlervrmlQwM7KzYeYn8HLvKThMqOlR39TYbd9rW4vb5eRLnVU0f2bPwjfRKB0pP
di7byszmnO/XNNaaiYczVmDkbCBW3SUrZ3P3YGD6TfspL4I7tnM4A9J1ZbwIYxfV
kdCyV2VtIa6jsfuchmSP3qifqPqhfqkomREPKPGvFWU3tQUFrvMST0sFVP9nKb5u
9isRbc752+2zYeLtdl9m54ERT4wClEhr76bAXEuo82uf1xsNDjoi1afUk5rcV8lf
flvftYPsqgVKWbT2yFUA03zd86B6ql6dDizyBZZ35qhXbVPKcopRhe2PeMC3wufN
lTG1vxClYLOcrAeeTDlyIzSVAGLzdqYYJJZh2g92xClZfRS+N5kFS7vC0m6x9lzu
hKU/PJwXQNp+wH8mdY+vD7IDYLjroWQ6mpNUqCpgmpikzt+gN6rSitdssGXei0Cx
BS2618NMgC4ZuwjP14XrSmuvHJ6pJGsM7CAYLHbvmAgPRQNSN55lB0SbdBYA9K3v
BpGLpk9ow0QUuK1Zn+z7FS3yp9VENeOpu0MbqMs0x/LkYYnActmM8NBRsi/9W0J8
RC0GRF4x8uQf0Fnj8zXaEwoaCn7t5qhY7BXUCc/uo1O9lkv2y576ZEa+FcKDXu7h
8+qd+4RPYq1KnP/uU7s7HZbBbkoKgrXG/wlkBqzVGkHM54yzlAt1z2nxQf+93Bso
uuRqiBSgDE6gdLt6o+1PAi/5ORau2OBIwkwoKA2ktGk7gnWw3WJLpE66rTHmwp9S
bZCoS0eF9Fki/GJuWIz4jdQtyKtp/6KCtcfz0uEtAHwczYfwgq5FT5Zof44Zpptj
jw2UVgth4HgSd5Y8dDgNRd+illLFBwipr6hISgvIxsDm8uHXy7QUhBrfI4bDpzd1
B6Fx4RVA01Dmw+l0i30WYdBV+2XTwK2xweOliI56+VtNqhq+/R4zwLHTny7DJZ8o
AgCZyHSmhViv/x+et8wJBU5XB5j3t+4X45ffeZ2VFCNk9IRFQo+CrfQ+ZJj4wUbV
YyBysiAxL7PcQj0p0wxtPHBd9MIplNWf/A808+rxAO+XZo4zdtNKSn7mXPXukSLL
0/SROM6E+LFIBHpkXjMvAVUAG3aXq9RLsl349TJgFWWihq+Xk4TjeAIoCGJHwhAr
XH5gzaEfIrtGnugb/3mjT5TrS8LWOW+ucCiEEcaaVhJD/faYRL4PR3X1b/sSnqZ3
rdR8liR0BZZANi2qdTk4Vj4DaEmTA07qcnT/k+tiIhmGxbqEOcfsr564jD4v3nj6
qE8bDf040zGS0d/GByPvVQEUjiz3/l1ADukUeabhPhQ2lcymaayXFQys+izEhawC
u/aHNMHumyPKvt7wyvBbgxscAdfzfjr/irXkssl2AU+IIVI8Jd89XJatLKFJC2hV
nfY1z8PfVH1yTS7o2MtJXZHJO/wQPvRHG//6BWpxfRH33kGEuOjP4oAiLvlg82dz
jeKnSs4oatjj89dw0eWV/G6vdBLvPuQqZbnNlA5fkXRE+if+h8xrTN62rGa54L7e
Asq33ILVvdYl1j20iMiwq4B4QFO0s/HPk6lE899l9tyXkgxhfO68wGXuh+5KQDlB
1UrcRr9R8kjBbdLPkgnHeklo8+V8gyfML20k5dkAWD5yPPNHU3sXKozJvSBgbj8u
r2zYQZmfx6GFeEdXcXeNVAIRpwncLzAnvEt1SbuCVUdqrAsGU1vcVh+1V7FIMSUe
uOVLYJ1y6VqCevXVc2nh7/6u8DKasdnQmyEvJ8Sx2PQL+me2746HmpzWka3vd+Wk
RiTQ0rwl27gcPrFg+DsUJ91t8EBMbErVFWXkeYstUBnfpULlCechfzwaefSIaVV8
GsMR8qPCLvHrLLOABgzHuevuW/QdQgh5w+JJ1e9hsBCoa2m1QFBvuwG8mL+YM/YI
g7O8sTXVc+EE7uTSZUylG7k+VcvmgjRPskDjkYFPUhpROAOwpqpqEopctmtJJ+sp
/mKxpJ4LO9hu3pYRtQ1cf0330+/ODFsJxiKzgffI4XJsJ3qmNU+7rjBaU8U6Ukug
0teao5zg0ogWbkItSHDR8lcHh8k4D5Q0MiFd3bfVMGGb4ykd+lVYp/zJVl0CLaxg
vOcfTTxwK2fnG6QzCeYfDOsC+wzFfYOnMEnyTLugaoaQqma3JImzhFIAewhrhsBf
FafQKaoMIkfJrKVwmv7/HoaQ3vDcF2s07XK4NPNx3YTSun4YlU7SPjyB+LPUn4C8
v7D+Z2f9MDBwFFTzQA5YdhKNhm4OJr/cbtIRHUYx41OXulQXTT8jjJ9eOuTJzy0Q
WuYJmm6b/jbXsWLBVIicaKVm4MKg9+jO8cd2VjrwNxX9kzQdyn7uw5rhAgRdKT9E
k8EHKqxP+HGQn9j6hSm5ZTysaOeToTc84k22/xJSjwmiAsvaYjG8i5VIh52D1fka
g9bxoL8hNxxlPNl7H9puGHPILxLyk7OVRvMJrNEB8KsBAqeM1ryTMLi30WXK43nh
+NKv32lvS6MEPD9jDt3aBQQRubqeM0bW4d6s4c1C2IqCjjgc4M0TBk28Sqft9ZZW
74Hl6bd4kGlhbkFmJ2lQURcslZ2bcXkt8ZADDMI1o788SfDW/pT3feMBkKuU0b3V
QZIPjk1HNcxFUHtX2ICBcw5pXeExmYL51l8vuvQRiAUSD6gxBafApLmQ3MB+mq+L
e47Pfk6hSprzKafbZVTe8ZG1N0aiYyHzf+XOYS6A8e3J/I7T38LjvtFDmuvGtv1w
wy7IkiqrvYfnthOHOq84yIj3DdDqJmaGvLeZYTaWzzoxrw3Qaj+lQvJ91j/Acbf4
gkY1SmamER9y8FTsKkEyxVVrBHXCsVUBff1Ow0YG3tK3/MXWutLXz0ksUut3UFeK
u2dQlQ13pFd2DBzSDeV4k4KAQgu6067cqSGC6wnZpFxubv6w15bGk/QC+aGt8MY9
Npw7Pst9aX4kM1u7tlpZ418UWfiUdHRyNGoPjfIbydlYBQ5kSnhPJpTDDn/5DWq0
5R1eJ0P4EVwEI3TBEqfILwUJ/65pbFobThM+CJGK1Of9/j/XveFuKxNN5xlZYJD4
aCk5gkPzITtJb+PW7NrHO22Bt9mN+oGP3HzYFTY8D7I2AP7OblPHJnVNoylGM25j
0n0kjEJPp5B94ECsj7CpjcuLa3Pm+oVhIATJom+rv9armgyRkC9oPQ/XikqoYSUQ
JEMFsN34uZNHnBK/mGeaAyVeDdq3AbWiXGGfhhyLidQsb8CA5oC2UeT9foLW6ylC
A3gyugbIFl5ChiiYvVMyENgJGM+smvQ30DO+j7mugDXszewx8wKM8vvny9NsHe/F
rQA1JR7PuBqIaQZmg4LedMGwXJyqQTIdGLECQS1pLcS/8XEbb8O+LDpLcUCXRjti
Q/DdfgMxYXizmSmnSwFvMB5DDYN71fgbpNZxr2zxt45YmVlpQVzRFxRMvidHGFLH
lYdUrkSYSQFTjhBwlkumD4zm755QntYgGRM7K5HDQ633kPLIxzMAe1vcYTO9hPJo
8a4+9gNYrmlJH1cHfIjv7HAS3fK65G58SqNdhp/Rggfk5uifkX/UR79qlw8ytNjk
u5j1D1qJ5HuGkQKUouCob+dbv55prgtaxqhbCwLel9xuK74C0DZarBp6dTuTcI5E
LbPcbkPrB8YcTbWolmV8ARdw9dJ+rEYwCMTpInvdpA8NrnNa747BW/s06/H5oU71
rBu/8dsco+YnOlNcgVUBeJY1gMT1R9n7tQjWNwtOa+g1IVwRxt2hIYKk0iG98tQH
li98BT/CUuFSgoDc5YhRMUJPnyfoCsm/3X63zXC2yNpTRrWS8LaClVSt2i2jP4a9
asGIWyhwjvoeDd1qzDojklN8+UdcmkKZV1u7/MKhb6h5lGDANv3ZzZLkXdcRSS3W
C/QaveqVO7FqJ7l+6sKhIyhVsmM+6RxmpPWxf0JnDLWJxRnp/Wt/XBFIlg4KuEuG
WnM2nNIYtL80WvH03fJ5Em6S+0Ma4kTzmDLR7OLx68LJiV/fTen7XShnX1UG2axw
Og8rFMekNkyBmXSiRz7WlOOYZB12uAMvFuwy5NXsQP1TAVwh0PCNNag5KueMzc5R
z1bsi1F2YuS4kBBiV+XHjlPNF1PTaUM0N59vLK0zDr/qk5Jlk3WScNA9YFo2GeGE
cN4Yhi6OB4G5FwJntJqPC3aRacOUG24/oKPUGehpycs1sC4OZdWHvXZ/kUdRSnao
7CUYf9mOY7Mtan8dKR667AiBpTS5hoRizE+jB5Ca/+Yon92Y2yLU7gdjmP1uOUJT
HGFGBaYfxn0Xmuy/zwWO0rvwBR7OxwrpWP9Zx7XWDbBsXuFBlX3XEZIKzeIU+GqM
x0Ra9U+S0DXN8nZ8rpwZBtSv1BAmZ9N7wzz4LQf75I/OhLkKw3DDofWn3ksOCpmC
XSWkyLJ5/yCh8ggz8XLdiOUtbA0E4i53WutUDWnHaYoW8w7OPaxL2LN0YGa4bl/y
bqDXygTEpubjnzHLUojCiy7D1b0FaN7Qjayui9hL/HSXpcrawLH7F/bD+Zf7z8YU
ahXYAPtMG6/J/v49AXDffcIWA3m73HvKb/MzbiQNF+q7YrDlzgu6CtX2d8OTwGrl
onS56+hAM4Qynxc/Qgar+7n32rexalhlg0lOuqGZjCodp1ZCmABNfP6TK3bescLx
K0L8Udx1NgPcpAx2r3S02x9CR5fSnSH3mkGUpPZnGEwn3t+IPBiib7qzu0eoNEn7
8EtMvBDxthbhE3krPF5CgX84hSJAyBQDbnRSRer2PY35Lcm4w3BHLVIznPk88r5t
8uOgC1USz0yP6/3RwP/tety453Z2cRIu1YIR2oG52aC4WAeWrAKc+B63iA4i2OSr
ypB76ncK5LoDEI/d/d9WVmu4eSzF1WkTyqEOC+cj7s1DWIubtW+giOAM0lKyjT0g
DjcQlStBLr3cJJB4wtl+Ib5bT+pIS94d2j3wmXEKba1EiwY+4q1JMsBO7wegrfds
Vw17WT1sO2I6d+JB6y8XkQVYfU5GlHn2lCwmLsJ7r47BXROasD4g9fe4pEcnqziZ
lc49gGmLYPpgQfIsplO0rv2dnA/PXPwWuNnXFqFIbpVW6fYyEModUJHRg1Z71Ukb
hJnjFkmsLvdbboZh1um2uR1DHjdM1T85OzHmpyEB1zf5Gxb32DupA+XkbrFQS6X/
H0Pgw2Q+n5J6ZxNLOsgRR+qhvGb8bxsokIl23db0VvBBHKjdKwLYqkEl9ay0hJ0G
8mFByp2kJEwGD7tPjKKGcKOWCzavsbPVaOE6AsGKSLdO1ncHCcEYx5NJjJUQuoPn
41elfly3vN1PT1pQ9BRlXpNR0wj6WiWj0j5O+iyfsJkcWUX7THxTkjiBYW2sOmNN
tQpKAhP8lC0HNL7k7fAUER5cKW6deFFlxwWS4XgTNvSv8jluFfX0cN2cKBueSbIa
nj0btrEG+r3PKfv7UGPJb9BnIsFW/RynZ2WLEAsTTXbwYbFhqg/HOUWM6Ei/1K1d
c/8QKrlyhX6QVE8WvFprE6KqDZRydmeCZMJ2kpheCrPZF1C7op8GEue77QKCR9CQ
+z1iDUjplHkS4mMoG6AsomY5JfeTUgiY1Q1pCqbiWdCnnMIOttrw76/1Xjdty89x
hrEMfJRMyikzKTCVk7sTt22tJgUc1iYRyr0eXQmkCFI7QQ93DH0awnrkd9XxlmV5
/xZI0uKk7GNrL9oALz0wfYX1cIcEsO4c7K+U1Ub2CUDbCZDUdIF2TyMQIOX+4L+k
dvqLFYep6VLmPNDS/0bYiWgiUlWWcSFwgCuhcwvth0yopifFXxYWcIPfmmWeEU27
6WY6SmdbwYbD+2D+O9XHx4EYJ8YbMekLC/MR9KsEqPWoluapI9ozuDuPJqA6X40g
dYFDlcwcw9Q/3bArapHLw0hGDm1IKsEPqozJhnXhPUBIG/6xegiuCy6Eb5cuswa+
QHYP5RvnK1ZwXExpU0hmIgn25EMZuiiSHBvppblt9I5O9Kz6+EF/zpPJzsejdt1O
bUaqhvv/F7nMyEhc9CbdIggPL0mxW0XMb47RI5MdiAZOBvZOxQvp9dl3pJM7bQuZ
eyuHXYT/tp95a6SOQwd+r7OUQkBa1ZGdS0QtKLtD7V6PD9n0N54YoqDsKw4Y/l8/
z/EmjkWqNlYYIxjj7fl2LzRH7WrQN1NAlQBi3548WKvb18QFozWgZO5YfhFPUcVj
ehpK5HSXhPrEdSQhdQL0C9Bjd1pK109NRDbu/iDFsHdHc3uRc3O90+9hHC9+UuiT
hOekHTkd0WRVs7VXNU2Q/BVMQ6GmWqhjciV38o1JJ0jVi3vxjrbd1mHUK8u5nY4I
RICk16+XJr8mEdcsSOAvQALeOPDBq/KX022aUT8R6G9QlkQyup2ha+GVFsbcTw8R
kgV6X25sfvj+kz65KrAo2l7vWFEA41dT9Mssf8H93D5BWPNSjpbCzNm48CUtdkjE
heIuUDHPpMjkVs6iO6uLAV4dI7XTI4MAjA8K1Ky8Clsz2T+/1SIV211SHkakcf0R
Aem84H8rl7dHMbKexXgy0IB8VBvd4ZX/e4rMAsGfEUWcAbHYNlSUPMGuCNc/vw5k
CW/01GOr9s5e21q/w5i8QQdHO2RucB37nAHK1sdn2rqtH14eJEOk9ggUtpAlAelE
3ocsvGer8R7Fgb/lLOqgY12jT0C+ULTV4hjfDc1/wBEQpdNIjTXcuGExwtvr/i6m
SBKaQAuEOu8iw7EVcdoBgbBybgz4eD+IRQdqJSApaSASQpoKf14QfSZ1DrWQOwbN
Xetfi3XSeu806nvCg0lFEi7vL8E0nRJgZ+j4TKN/idGQNMqry09uSQFJqqBRnkDl
qeoeuDku8doU86gYTPhrZQYJrCFALnO5huLhRfX/91fZ1BGf1afMNG2tkA7xjNtb
j2n41mjf2FWYJ5rroaAyErqjNOqQqfxCrhXlxXDZZghzWJ/ZCwN84VfJxuOlqkid
6idSM3FR2oQkzSISL57+aeEh3J0qInOY3k5eCTVTqAjUoLJd5WmVJeqGqTiJWH0S
ZaHjhv4CXwme9tk+DoI2mk494knCOgqPBQw17hMVomZ4D47DmNIuaLozRyzyKRsK
z0MEXlZm6CeYWC57f4qH0ExudyFjHBi5aIxBN6Rb1WWhvgv1zVRxx7bVLT15HemF
RLcK/sU0nODbmShXYjdxFCyZnd4Nzh1YFY4MoKurTLz6Q5r90DPpAqDxrgNVrC0v
QOAv7syFIYPuAZEDkSYXFi6UQl921JcM2ysKeH5jHLNZHUSNhUYjJNeJpVs1pkbZ
aTqx6k6mRUtHee88CGaBax4iHvqBfGV8MFr9/Somi6dhYNxf50EmDp6GcPDIo11i
FaTINH/hHAIASKS8S/5s51FUxokrpM/RAX45wvKTIjDgfZVP+1lRgOA6vMieR8xy
Agz8LO+dhObygrq9gRXRpPVgULnmq1J8Biw/ul090NEI+o6PGEvqnwUjIgTtXYfW
u52H9F/9i+RCSmCPrc/XI8acq+WaUePjZuZXIedf79cXCaHfRzeMsU1+0jsUrRUI
0zxgr25xInG1EnCOD8TcWZxNshqD1EiRcBaaZyRzwVdV9XBASRXeqZi8ZsyIjcZg
XL1kux9s3QmXtOnhuhI7GKEZdThwI0VMxllKvUcSVFFe6Go0/nEN9zWMCce8ZRcd
u9D/Ty22nEs/Ib5xMTbtTlrZ986APau5YI+S7KcHj1dWGgqzM7X2x3ba2ritLRhz
VvaDzFNp0I68lcAHrkVkRBj9+lIMgBUGGNc6qlXCjRlRSBOzpTZwM41WsTuhuFE3
1A00rTF693QxinvMf/DtuOedIipIR1r9nGhNQU8VRd9TZNvYvIGPoxX08omgfZZ6
1CqRAO9hSyx+tBYkUp8pG+Q42VNyAmRm+x3g4a4BRj/m3i7GNtnBIC5DisRZlYRD
Z1sQyj4qsN9pdpyGf9DaHVOwpI1/XCZQAYrc+Ckkr7G1/LkCkAXgF4dSQgmkK8PJ
UZfycdD/ZKl2bLuzSMV7EU9Ylf8019Y8cBVOMe7Ky0KjXy8XAhOb1GsH9YWhxWaf
Ua3eKF3e0hv1gjZk5ncw5GhXbhiEKE3SHDmBKfEtPWEj0hSu2Q0FjmCKtBm0/PgF
2u9eIJG1cYQvZruaKeZWwC0a3OStgslaQ6j0mePae+TBdgsS9VZHXYPrgyPd50/U
+DKQUew+8MVoqmI4so4IbkJVZfMWDwDQ+qA6NVyAfTTpn8SvPTAj2tFTwbYb82JU
hPYJXErWLYfhq52K6wgAoCfhdojeSHoRzMiy38iV5WEIYnMhq0EYcoFYUELWPgaZ
/4soG5Es2XD0xdNFf7QD59lE/F/9Om5jYdwt9OXk03ZC5k+ummPr/Wr2J7KHqnzP
DWRd1MZXqY7zQLr13etG2BsjbE7Ms2mG33Rb5xiN0T+aujHKXHEOkhDanAJBPVWs
N6vaD0cRnYCX/pGs/f3FOG/AyqKMDNNM7/b7NZagX2nlWgI+Rgc6Oi+YsdDreg/j
jY9VHK73/tlEMzHIn/2YHw+vW/20TectuU/JAydnNhFQDqWuRoEdteoACM/ZB/FX
2u688K7YtjTG8fjoRHgpB0bZAOjp74RKWlELsjAe4AAUqiO4sQ3jateQtMiH2t53
1vamh43Xw7QqCthdCh02BzaZ2+Nu1wy94Xh6ZMAqOZvLvcGWxmbLQ1jiUXG53F+J
KQkAPVhJj+Okyu5lEBCgz++OmI/W/9WDuBcaNpyAB3lVjkVuNJ5xGAT7yKP31c7O
CYxi5MB21z9kMnZFgE5ULz7yWDSVf09nqsZAyjCYVuiE6x0AaoMrGZpGXp2f1ESa
rgsRNxr/4I1YpWhUFz2hYxmCE2Pg0Xoh+jqVkC1WNEeXRdFSXaThzbAusEtddaFv
lHiTqLAP1qhi5vXuv2heLCpRLOEayTbSJ6Gv8ObK/qkJ3CMrbolCjO2ekM50ZbsB
hyv3h3GyYdJYVm+4xcKr/3te5iRXK3VgIWsLpa2hcrsNYMdUsFuoVkxn6JYbi6zD
CQx5f+yl/wFn02Lj+H+4DoY14aB+KfQ7QSY+zJoDcRRlG4PgGRrX5T5L/g+/RN9C
bx0tts0HwTuIDXfDtJEUk4fhUvdOjiJ3xlO0t4tHNmvVitw8kDCpBaJxlIzGtCLT
oyfuxH4OUI0VBahyPuVFuxdpz7cYpoaFrPGk6ltN7F4CY2sngwX75XF11WTq8ZSd
M03wPIjIKos7pTlmX2q4sZbCR0/9e8OX0T8YNlNI9OWyiTbRddWNEsE2YWtRDsx+
F+d+BFftmTrlw/Hfego+Bv/sd2V/T3/VFQP6iE/NrM86L/auqJIIXa42r4JR69yV
XkV80gGm1ZxeiTq6Bfjo7jYplWj2G/IlSmoesuFoFLqNQz/xrmcbo79DrZUPuK2P
a/2EWwmgqgJrzZpObjMeLN0t5B86YDvFhLsS5jdFBNYPZvPFx8hlPx6sTTtf0h0W
YvRSTW4JkpIAPxcfzE9UNUNiauB7sPwRwNS+a0ZOH9zcfRuBvppe/BB2uq1pqWPV
Qb/odStwf7EBT+oqcBfp8fhlz8MJL5VBO+kTTIj2Fj0F3t0BIbO4tL2EyrCdwZ6T
PMoCJf//UGA/6IuiFWJUUe4ZS3NB0m0fkRNHAQT6vHR7W49+AXIDzsDUtm+L41BH
FiW+UfR0zy9LVVl8O8gPZwf9u9UGE+XNMvdz5yX/xmGljI+JxVztb452rHhw2d8w
gpif2gcvU8GgjbpXD9UlyZCAuSB/KiGB5sBl1FcYvRIxngx2sN8FqjTbzLwWGN2A
CRXAFq+fYbFyfsy6Lqr7BlMMzOtvWGrrnfYJJwzHuiNuII03w/sJ/0M1qBRkEFES
7nrU4MIf2H1A8/jJonAcEeS6fLs/+EA2GHlA1LzzwXJlHukf2Axyuh8W4UacGLin
sin3wGkt/jgJ7flLNThl8zAR2S69a7neY9/FP5O4x8tQA/ukHYnY2avz/vWI7qd1
MBz6u5lAmQ1YzEqUF1kWTLpWP9lXeJueFJSHC6bquRRAJRWD9Q1McXeHvqmkYKAE
OVY3av/2gqkKMQjTSjMuuMmtrdoKbM/Fs7IAtVZbN8o4tcsPPSjabmvTKL6Z65uY
D4EtMXtDraMFK+LSdK5v2Xq6OWLB5BW+rTg4vphDNjHFY56/GhJFEp+UgwGzcaLy
IEdis6zdlruX7d5iZN7taem6lvjReTEspBOb9OrbGgsMk2R4WYwHt6ICZhy7/c7T
EvVYb143QT1uIn6X/FE3jcI0Iku3EZuSdOegzpliPcqWkTIAImz1OKvLrc8hfKEV
JM/ZXZfQHOlb/hYSL08HNzgPWRzYiVB0E2uCpC+7p2ampFBsVXSZKy3Z5VTMaaBf
tkiZH5UndyrLGqcd65FIN8wODJOPcPiejpuJWyqaDMP1y3rry4Vu+jzbFhK2B0Rg
XrCfQlp488jWM2Q5mctjOrnwDKLDyR3ZhOaZRfi2hf3WlmzU+GmdO35pp3jAw3eu
KHjyBHU6YpV605MiD5TO3WUxojBBubtmwVNwaFvPwUlC2OPnyfPyXBDQmASd/foW
njvH1vMcXYFr5odXvb7nTjKfUxfe20IKnzP2kSXyvWDPlm3F4gtZ6clnjrEqLc5W
gSYd2NJiXUmTkN6mp36h7YXzGfGEMQPwIlUAN1RfixcgrdvR4D4fFYEV4fgsYNTS
nL5MfG6/VFtmGiCSHz8BJVM+WpY0h6kgVLPIG0/s2Tr9wzHSIejegUyKMHkhlgyh
LPmiIyKlMfw6Nwy0UjR8IhbY1GYjM6tVl66IQvDuvklG5DHkbCuZFKAKRbNgc31C
AmZDF66UaAnjVBmupZhPEyw83Wtee8hbcEiSUnJjbYs03OlLaFx679pU6X78+JHz
4rseGesh/BV6vRaVG4qANJxguYWXUO+EJjyw+iC8Mafykz4xxAodLV0VtooH+xBh
feMO2NXfa7p7iPZbXglWB/y7qJe/h8tIT68H8udguF1d1Rp9hSF+qke1f3UZ8mo3
cLnVcfL7bJvxK22K59xEptB/H6YlsY9zqFvaykmDGQQJwqvws9lIObOR1WjcWMyO
AiVE4AMo22A8dY62xLg6Jno3bKqVQirl1E/jhIMSb4LNxO0IqA75y7nlHS+dX8B6
f40vfkBIQ4g0Pz/8TXMoxwANUY8aKUEP9yqAHsROhbETDDx8Xw/gU7KuWMkPd2J4
+h280ebExZ8gOQZS9XquSnAvzikfMQRYupgmFtekJShQLGP+z1qMjztQnSxfAPc1
NTDyWxmd3LfT1TwVlUzfBJmmHT39pUQ9rKcq7GwIMngJJPpciotINg/SaIEWL8Zo
CIp2bhtVoIUBGHIuM30l3Gda+K0c0rlH+jUKSudGZ+bpWNy1/MSy3BjETrc/327e
Gl9MwIDoq0lMAiBVfdFmjOzBhjSijjEQwHN14XGR8+cnxnVH7FksBElua8KB1iGU
uuVAUgPx6GoRLwnN/aMgn60nng8cVFR+awaQK9N7289so9e4MbCvDMuk/hzSnhUz
ImqHs+Yi8RXfeV+/ucVIAzjmIoonJyGsGziu24Mvcz7jLFb/1e/tCwSWVh10Vxj2
gLeEL6XPieHZX37GSgpgcG/tPbpmeQ0/PhAJADdFX+R0PsNFOhEL3X8AwW49iH7j
GcbQCCQiSdh9R7g+r/7islAzOHVqd+UVU17edjzUx8whzfKk05MpUL5Z6VZo8BeY
2M9qA4pCrMSMgvqduHpK2btFueuS5hk0xxPkMBWIffBK/Jj733kWcEiJHJ4H8oj9
lOe6DGefsYpYrr+kbT7QggYaL6/L2ABmguouheWBE2vymnVGOIKlrzKSCveAQSkT
VG0QwJ6CcqzgBXnMMJio28iXZHrBNmp+2c2oUDQwsyWzQ9g4BCbL6XlVsgJHa15y
3Y+N8mOl9lECd9N6QjyTtu3PAs1/QOwoYrUn2+eINa5cSt8yGzAUXzZQ5TX5Z++q
ZVco3N2pNVJLMDN0/Pl4SaTRl5bHzr16YvqBYWbC+xwob3dZp9zZ90cL2OD3mvBd
4Jg3f27jHoeTnKap1AMp9slo5cq+LSSEjmOgl6rzdnNlza83EdXKMaj/G4T8NLxH
RcG5NDf5xwhgHzYvj8t5Kid/R4NOJh6eSruvUYtAfw6L88et1DFVkiYjEkm8ttFJ
fiPmWrijR86H9bAmqkl6+N3Ldr8Kh93XrfrLEl20Kpj/ChUN0K/qLHyCaklERYTJ
awzcPobe6vh2VUWAEMYxU/vZO9m2ko0weqn/dNmy22RDTrxq5pLYCcWRMH+gMixY
rsvY3AZRPIDVNGBjn4HoUfgZTbFg8zEyNG3o5FbcuJIoWcRyzXV94gaTQ9h4Ab7/
XwS1T15N81gYTa2IS56EOzV14CMYWyirS7/aMa+JgI6VQ6o1M2FbXcumn0+An9+S
C1/sZQP7FthT4yGOC9jn9rv6AbFKiSSz4iyE3hSficawRfM5gTMrYN84D7iTXDOw
Sb4GGIjjBDcjKya9D4Vn9vn5xF18G+ns47SWB3deJHD706qBhzx8T/t/Qxmq1IDo
h6nXRwsSbgwdaILnRqCeKZ8tTQZxAx8CzXcIlzhQqv62ZMPxZT5Pe8QU5EPR8VFk
MDukUcITm013icybG8jdlfU6jw3tI3OkFdcC6jA/T/3AtpZaUTsIcUd46WVlicXF
lY30Cp3XFwHGYyspT88M5+7ESYF1ZjdQtlvflC6JsbAG3Y1cZJ97E903Vmp/iynF
jmXa0MjM/dQF/sa+buTob8wrBUegfMHJ1pTFrv/tanvtiPgwzzgN9RZEiqwPlYK/
ztugh6hmSapNVGwS22bc4aBDS3m9VkKjxbnK4+dIlW//GacOJXAfgePCqJo3a1Ln
hKjMkZOPOOJvIwj/b5fmKYWGMo4Xs5h5RwAZnAz2NjETIaktsHMlCPkfb9gz1qdq
RatBq/FYrTBBoql3GexFFem1ELO/8MusII7KeidSUJLZN3mgIKh8hjDUZ4yKJ4Zp
ZfSxz4qwUtGjmZKL06gOwrnX3HrogATPWgohY5rx263RsXh3frZuvIPcQR11rLYQ
vpqLMOLtmhCVznC0s3ZJA1Rumi61ysOUNer11YbwanAKaDZq4qYixWX2IEpIm0fb
Tblg4u8j36XSWmX3RBjZMvI4lvtsBhu6iSYCpagPl/YUV72t93YEapQucApfa6YY
gjW2qTaPxJPSMlLSRUvi3ZFAH1HYCX5XBCR1UDzTZh6bk7oUP8uB8iZI09FSlHCK
QiZTRcT8aFqktTIVkSgdcyR+G0NBu/MMER72rsx0U/agRXEen4WeqAYrq7eFrYSH
Xa68nHb8oIZqL6wnMmloG3DXnQRsR5uhUJ3/T0E6/rCJ3EAK/GNdY6ju40ZG2pYR
sSwOxkaXIm4177Tj5YJbPYJ+9159QFNB+M/+cJpu21y53Fd3zCAL7DNsALNdv49L
YvntSbzzJjs1iscpV9iryBXikqxurXyQ0Y0DuqN2Hgoh1s9VmELt/yKxkKpx5Kfv
SghcD1bA7stvKVtbwhI3iCVrbCqWXfGMSX1zsnx88U+PAwxAdg7a43+iyjWj1PEG
adLlQNPc2ctFdmoT77PsgyeeGYy3TwnFQ+4yfTjNdpas/wjrgbljH/3CqyQjko3j
hbq1mbakemlTwt7uitAI8m4KQ1MwP6Lu9tOl3mihwXjHmxzio0WWYeVGfPeJWoAV
1BsgSHxA4Fbi7nqNU84Jz5gplCH9YSb9XSzZReRWejOoFRiZxuSyG317RtIt8Dq9
IwJJpBet8Bkf32vh/Hpfek/w6Av9W+EWKD9eF9CxjxU7WtJa5Jbi5iKUrQ69cfFM
n23cGopI3BY/Ww/8N7z3LT3vfBtvflMqXy8N5Z45Fh8aR3nfK+vudAmNC7S/pbvb
kFuWmr27GendQ/pnC7+utuaKYVppMdE4kvhknPKI7TQd2UA49MdBstIwprXj9hDg
UTKxmsgCEPi2upiNyxBdKc2DMNAMd5eQVJj09xX7Wqd9Yqq8GtQBJqZZxM+eQotV
lqH54SrefxJ+tetN39dx4SmwjESO9ckVvdEuYTd60cHzpIbFgYp1mvNEyeLubTIB
1wMo/Ns3sc09LZwBFP4a+3M3G83QL9geHCkJHuVkXA2+Whu3BMSwF+gPUIidree2
etF/7w4Z1+etIJku2Rpj7Wee2hft3Dj4kSAxNyv/7C8PdyXoru9pnElX3girrVQ2
KVZT27PXnEVE4i1H/HMzadCmKFd3ZNfPyq7eP1EgIxiR6siw5iUIQ/C4I5vZ3UYC
rbq7wAT4OeVwupVZivsobI3SCEcfnnEn5EoycGZIBFZSL5u5Ow5kBmbq50l80Kou
WJXuQMVgdT+hGk6VcpPfhAzyiFtIFKScClDCNchlYtScI+gyeifn7ZJkDJDFmAsb
l+H7rIh58lrVnH16fpotogQaBLqE5vNamI0M9u7ud1gj3LykYO86OWqMfmYOZ3WI
1GKjdSpc6hT4mrqjFuiaMdiudM7T7d1WY9YN4Y92fv2rNflOf7Aws3Pl/LwlLETW
NCbdUeIaNUDjrofh3/QWQyAjM6tH9u4/bTK6Y6iRZoRqkTYZTGUWGxPYSppZOBqA
AO17XHVpiriDzUuOUPETkHzlPSgmNJA99t53lpQDacKKYfKG/3eTT3mVojH4EjwE
cjdaApizTYC9SR5GdTXUR4kLNzw7LpYTX/oKCNySisLHqSjP7P4KXaKBCIYdEz64
ZkdAQTo7FzzNZIxzgjUpw3PRrCKpRLSb3oARM9TR6C6n+H7vxlF5+K463YzwDXvf
VynDluENrVw3o+ZqYtYL+YUOXvebynwcOGkEeEUPtVSPRokKarR5pLKVYEZ5w44q
2Pw6QoCLL6m0zJ84Di80e2W6hWkaTrbfIRne7PbtxHXPk4sAO9C1hNiA6MGFg8zB
zLnN2LJDPJVW8icLdKCE9tVX+hBEZlQZDYpQ13/ijbKPedZPKbXwTbmTaNcLKrJ/
AF1x7wlSeYMGxtvoDf9anVYhoKMMzMA6+R68ESwjx3Hu2R2nRwezNN/wra9sqrE9
BFM8gP7xCp4TPkUqI5QQEvJMnVw0neKi+WRvC37FOxes/N3K9GiDF77yJFu1gc7k
gRpz6lveX/LkM2droCHeB6V5tYDfXfs9qDRa4qpJulbGLUcDISBRLyHK+x1hUwkW
IzLozg9OqbrzqTPI6ePcarE6Nkl7wj4EIYAOmKZPokU0p3b3RKhkU1zBvT2Fatos
QxPmdiLFHqzB5PbKXP+5WHUV6oto6ekSiCXJrmR1nccQrNewyy3azH4ldRhpJC/u
Nrk7jS++O0RjAUiqtoVyE2mmhxBYLPl8KbJ5N9g4Yw/hMlnTcWL+EXF3eFozFtpc
Y3wV60QZJjMm7kV3QGvr3WFfovff6dsyuTZppovJ0YVrMdFTjQZCKUqnOKc1q5tD
tqZbfUgtFibfgDgoIqbwlOkl4GjFrNEXd/1ICs5SMC2BteGQhXgHYJyu2xeGk2KQ
4bBV4zZAh3FqItdhYvJH/OlA6QqwWo7AHaEV7+sehx1+LhevQ/2xtW3uayWHFgAj
InB9DcAxGCwIqhNCvel8ArVBsFAb8crbFMV5J2kSzZWuUDnmUeHRmYbggExHAJFn
xRaWG6uHsBnkIWcYX3WlE5tkisMG99Wa9VlcqF0JYU7kLVorjwFmSWQXJjI8mqH/
IjnB7GfJk/TeeWv5q+lvIpB5iwnryxhmELMeC71aH+tWPgVhDMscrFFNii+Lf5Ab
fzK70vc+cyfZYvsNremPEUUN2ZcFqJFepdvPhBEcg4H0MLdppaZ6cuk0pQKhaS2D
Qtkyuil+rAMrVem0XmbU3OSCwmuO6XDxnd5n3ftxfuptJMcVO6KgAXWqXQr6DSXR
tGCriI5ob8Ue0Kt/78ueA+/FPDjMaKGZNAO5TOkF+zh2KTxWVKdSBwDKaymTPUPJ
D8/qAZk/YTDvUCOgvfv26k6n/2X+w87c022RpHQkgW93RaUxJCnbwJG4EUu2eEca
URhRXnOYCCJ/86H84cTRD3iqW1GBUcgNvMv9AmrxdqWBqbkJodcJg4cPq21YD+fP
5wQD1g1TO3PHR0qPGhzqzlGbjM9rmBwmUrPR5rh6aAOV0o/E5hjIbkqakI8/ldYW
Xr8CgLbTudq7/EJoY1YFZKZX29649oT4zG8PMFk5INfdIKC0LM3FkzSYTmZ+iajC
7h18twgMj+30SZSRnCI5Dfim4awKY+RElQLH/pXgDJ7T/wPvNSk1GjzFJV7YKXUt
XVK1fjpZ93MArtBQk6AgiWpxxSHcziyiI7krkrXYZUi7SrQ0vxQz5TyCWPZQy4KA
woMB0hPkoI4mwpcMJBY2YpLVCMLWKFZScrbI/q2neEuLk3/qp2FMMtd1y0BOrsma
MiqFYE1Q2ySyUGbwjSnFCH6VPVSQy4Xfz4ZRxuvHkKcahaodWZDFdo4ve904xPxI
knmNGy5LOGiPyN8ErgTDcjW6fi/8n3zz5GCZnpUHg83RwKjQehr+bn2QHSq2qlY0
fhYP4oySrR0mwAneiHsJFrnc6Gh7k0gUszGkpqBMnQpcKQgpkqb/9MeOpd0uKTED
Dc1fV5q8z42dosC38S7BN6/Eo9PR+0qvnJg4Gp9+KUPFmeBWDd4FfTv5cXribtVK
pRB9MdHVgrfVOWVH+RQ8Gygrvb/pN/4TbCqwe2mgP7OVUGfTSVtRawDgy6wHPt7L
0mP2KQCWT8HAT91OFvzjhILF76jkwuRLk6Wdlsj92I4rLjftR+XLoO+NWVIZvw9C
J7Mvhu09IBX6b2omVbA6P+isdT/ckT5aKqDZT6ZKEjjE29OJ5zYNFHu497ztj4wE
7QvAkYNHvMDaez1lZlXtKdZYVb+wWP5Ay+x6ZVA+KC2rJv330DkNujv0NFG28LZQ
mx8UYNJQrs7Rf6PUTn4yu2EcsdKwwHVaUj05zZN6DE3hzI+V7U0YAj916YWrmH2n
O/B0xHt3Vixztf4F95lAEKHpP/sC13+qOMKYYPfJo2EUi11s8bavMLqy1/2DMxR2
lSa8iCtU8Ksr9oCrydRyysEsdrwG3VVhWPcQOzpNUN4b8eNybcaeN3d5T2lVCkjZ
R9ZziwaWSHSNZZISKBkgGV3OPGDKM1xVUH6ZEH6JD0AG0HJGyxFed/1y4ve3NV1e
TG+LZ5JdrkSbwZ+flE11k0HxZNVvZa04Pd2WQtYgXK8AVwpJ+GPIsNioQYMTmUen
wXaL9TnfISr/p1SNMJ+ozVIbVJd1L39JZsTaLf0QSiscU/nKxtzZm8f4HaPSLv4m
ps3j81PpVhDpaJ/dcER43c9EeuHvNHlADec3CVT6ir8EXdq3YLXEK4DvsEB6RjDw
eGyllJ9A4QBHDQQt5sJkS+HH1/7l0JMqCsKn/mziHR8iRQy60xsUFiHx2yE8eFmI
W1kLkqRd6KdvjkUHibnFPRLaLcujRwIuFUPqDx95VWMgDlsYBwpVLc5Nelenq3TO
nenUoavT/RVE/HtxjAuOFBJwUVWIVFYfnN8wfa50RxnfrCKGK6A1GxXj6wdMdtZj
waMPywlZYPMZ2adNg5af2TrOdolDSkycuu9sfQB0V63/ieeU4WwBeE6vBdRYd38U
S8eYFzGw8z3q+89jokOTAiyBXCWhbuo1XYLtWX8WzrQEL/dOhPfj0kvtKe/NTUbf
JQdTyHbx5QmtLdFSMhKP9YJIUaMbBYXdFiByXo9GkqoKhmck7xiPiWcXom/1hJq9
F4wixLVLznMoFg1dDzPb0h/wak6sGI9JyfH4qTw5t2B8P8NZ8cXz2yuQkGBlYYbv
leL46nluDuUmcrQ3YpGlVLDeCbRB8v0fEdbMBYKHsg+LrLCN8sqbJXzD3hrbzu9J
jKUXXEA0UCEtVIO1LngZbK5fMsh91e11IGoVIN42YUrmyKavDEgSTKS2BnbFDvjo
j51uYgWq+4BKMB0REpS2gnIsHOjdH4PsYRlMu0k+pFH8t7YTi9JC/EuhrKFxH66u
M6MeeuLh+RMo0c/1i6nwputqsQCYsk9YkDqkQIHz+VgkcCmkpFu9ReriPwerRvYe
j98pZYzy+BO3w7y44gt13JVpEcnzyQabhTdWNaTTn/1hFGk6La+q2sb7xlKTYeDS
4IGwHFpO8VMJfc8SF/OR1eGQE342KRmiz+c3iaUshng8NgO0jio+7frXPGiw8m8y
UWT94sLeCHi822v5fvRArB1HLKRAgmy8z1/Sk+xyvzffy+i5l6VZUSgqoIObZ6a3
CniEzcgxLqcdEqyGsRw6mfD1j7hDQ/JO19w1DyJOAuP3yYeGfwD3BDF5kUCG0fit
0MgngH60gWQ9upgq4p7NWJJe1Ezgx+BX5bopDo24MCMyXQ5EEqbLJEJWm/Q+uTVh
gkcptN+hLZCPJR+9Q7BeahU6yOJRRzPrcKLAwZc3LuRTNQ2sCr9Z6yTSRgM4Q9rn
mpMQI8uJHIYYtcImdN25lwdRW8RG505m8LvJUhbPpWAtT17HQSFwSdyfptor+0/4
O3Wp9yFISkNNE36MW92mLA5TifRwe+dFeNkLmMI8smasd2J7soWqTCaIcJVyYgTx
oFlMQ9JsHtsJD6CdswK6waFQmx8EKjAIA6BALHI8qrjBnoAePQvSUxzW9qhKWxsm
pJ/p1w8ZcmK7ivPUPMNvm9Skj/bi3xJ20TBp26jRvAe1IwVNxfm5I/hfhrsY4w1O
LKv/hip2pboh96o0jybjB0QkXA3RrUrslbiGmzRiOTfxB3i9Jfo6apl0c2Usm/+e
dYgFYwzgyZCUX0pOzVRpQdzTeRXZQjDnHbZ4A0r0dIWH14kqgjwlfbxu/QUx13Hi
0e87QgDbVezlDmoqPFBfAfYtLbESLcuSmRGbrCFy+1OgBkYxSuQOetUc1U+0jli8
u2/OrQe9YHXUJU0wT5eGsiLGWLYBIBsTGqHpSIsQB3BvLd4hUzGUmZzKTpDHlDbH
O74u4iLMRmkl+Pn6l7SlvIWLilRY7iX34zqpmzukAZFaOm+FQ8QrzDEFEJAj8FGc
6Xe8miC+cijIp93je1KOW511+N4Bifj36U4tnZoMwmAHOYg0lQ+nG3eC65xSZztJ
u7ijIreWaWoiMOBOIuuflnD0xhO2RB4yXzoCUPgKB7k1G5K3V/RgYpsALD4YfmqD
XWoCZamXAjmo1ZURSPx1R+ahiShsOYaJb4hg3b4Eqi2Lv9KShQTI87RWq+QpdzUY
azzZtuguEo4vkFA3lMj/8FgYBXRLdno/X3Ik23Jdp73sD827Kru5cu7LPRiC6cfN
k/mWaSwk97RWsoYS5Dv66b/5eD5BN5kLWnIihDedUyej9LZQwG/X5qVVsxtIVo12
g5wT6IGPNfm4hPsRHsT59+ztkC5YU4e/PgOZKSzdQ42EV2DTlkHabk/hhcLfB6QE
mKU5U29k7SsqrT3jSm0xCKKeL+tDr2aVhDNAy69jbxXhFym6ekh8SrrIGVBG/9so
YIyQJU4AjcqZ3GBi0UUN1R9Lv3JV8mmqfIn1gTfi0eM1g49dvZwviIBRD8NVtsh+
r7xb/1KWriKOcN7C7bCOs0vBnMvsFr3fqmCYQBCGeMRl8LmUyj+mIlT145wXEqT4
uJX4R+w3KBWB8dvWn6omUbtJWvxvpUJDnON5AYqbC0FzQuYrzCl4D9E+6OvBVZX2
T20bauVZvE7L8RF3ZKVEhXK2BhStmfwzUW2WEZ8YP9GzgniqJ3oPifAnBp7puwyU
CRyePHOb34fLhzXeX66M27X75FKnC+DGnLwLS1vd8gP8YwscM3qQSlRX8N8/dmTY
8aPeJ84S0ScLGSyxQnfGpgIJeUd9B8xRAMmd1CCkW2f41i+tD7tRYhuZs6jipHRR
NhcgpkQGGIUtwzksCl4GpxR+gsjQ4bhfh1bpogVjMb+G72h9txU64jBizllLFuGi
nVMuACGd0LG6U6vflOyZwdmC2VBXuaKqAnr573ORsDI3GmAbWyHmD8n1RfdAuCFA
+eQEccY34w2cW9fchitGbrlvNRJsAPzcwxt6Cm+O6ikJ7frnGjhm3ZgDUJFjKVyc
MKmRIEU+F7GqT5tUhlSIZJO88hTHMhb10BW4MqHGkcuDTejhcqNo94aXh4oMF5pa
9RYpEl5eClcQLJoxdh2UrUZ+NmBeOmRoqOnG7XdpKheN4XMblLh8HugaS6cJURYD
ON8laxd/YWeRZ2dhBB0m2MBWidC3TwCSUUteJ0/2mnLKMrXvuqFgGEuu1CrF2frl
2NihOWDihtE9Li8bDDTOQKs3Ac3VU4cHiY3XkholLfFILEa/ZnPTltlbAZZDsZaO
DmKo+jDX7SAu8sx++etNnsuqNOJqXB0AOaD13UTafXXRHvsENvLDI5L+jCZA7zBf
kF0dGP13YFJRkoq25vyhsizvMFgEMyK/9cy3VNSXH7EHLhiREsfVnt831s45Beb/
IZoohnrQ9exw9+HEBOrFrsEyqpI70q0GOxQSpiV7d5hCRQg2sEKHwlsaIdqShicU
MFNiC9fS5NFYq8VA4h31hS7iFB2sAUZuvJlijNdMnTYbyuHhgec3ZtSHfydN1o7K
nKyExjubf0wycwKwQ1iNFfeYlqoPiaO6kJ3hbp/EF0BBxTfkgJTjEp5pR+fvIgrd
+0BPhV0adUl2XK4HY603eAgePU8VuFVmWX4GtVbTC27MvqvtjEK4ZlG/1V01lHmV
KiBLN3ieE/Df0qWBowGV3URYfBD+IdIytHAuRHOg9T2r0oguOYgg3MRZvj5X8aaJ
M+6gbrgblyKlY6WIO5DfU8B6MgnXvbfAzQS0ZHMzqryx8q3kE2wOHraOO/XuAXtS
VLOwY9fqBcbyQraZ8pWTFbODL0wuvvKMe7vYRL9/8ztvZz982+6dgnQ7piWjOZG4
8PmZ/P4ybDV7/aV8P1gckO7cswLwikDlNmX+58jVbqxmgxP4SDA0q0SB/C++/vaR
yJZZy8ucmd40ae9hHexcYMjdupW2d6iYxbByFD7qqmT9jS84NzGQIA9HyMtlIB/F
A53eVd23n/FtHsb20IJ3pd8GBSTTrEkOtxZOdFefwWoOYaYXhfRZ/kjjODiQ/ASV
Smgb6tFPU3WETmj8F7LuIcPfw+HOC+MqTqCABQQBZaBVnU4kdoC8Yu2CW+G5m+Wo
MN1x+VvcgLDEI3TCkXS6NfN6tQehHDisgeSXj7nBPkpM56U9V2AWO+oHrq6pxyaQ
OEj/KMfxT6Y61ni2D/5TDM+WnCKf5FqacXbIb7vm/bNoxyJOiQN0+QF05bdIx0pz
NVyN+/fWSa5Dl2GKGd97x0fjKoUkwC+YNZeR2XXg0BPCRqIEwyQ4GWSgcSHzV2ki
8ZgjLsXu65EdzZWOXQMJ54iEb6vcvoyCe/yWCu+bth21kJ75aobZ8m2uM0Hwv+Ho
z5LOgEsgco/QvyRYdhQnTy55f+Ze59fWLD08DG/YzjAPTgbukZad0SBgagZLzSay
KPSFi3k+CpZhzdXVhITfCEYAXDzUSEtCNkNqyamjvKYviutRscm+w4LD1+PTGKsG
gXN9VmFWWjETKrV4lGMBqUJFw49yzxApV20JNak/qPDb3DI9MQk1uyi6nVR89C8C
5lPmPTDI3C3WCQzLb98b9I8LCEU0W8OQssKyByxvYXrM4dIc8YSgWAkjFYGJwJjr
NWDHgjXPL3nODrx87RHF+Fk1M/brryhyn+4hspQJ88bcrO1sfMaQ562vrRcpLqmI
+w3uZbC/+rcxKAuY71XAfW5V3JUyskipA70FmLsPhmihxogiUBlmt+EnavGoBVxx
nkBl1jZA/9mcNVdHzpHieqRaDpJsQB1xSN30HA/gF38op8PYCrN1yjXahWKtN6J5
hn3HwE6FSOsAzJvp7lH82CslGZZS3TqXTw7OShenKQ/jh1dXXkI+iOSf8OCu0eIB
d8Zf66lbh4mAKbmG5H+Vi2dtjbrc9uvfWCJRh7aJvBbfUZbPxFoVEUQwd6OFRHmp
5NxpmV/b0NdZtP2bf4hszIJQT+1dmVFk8sLzvzj4/bVUQQU+PEBJrh4ByPP1sPn2
J4pVXdBlHHw2GQpIHTiTfg3GgrxFyEclrrQXjaXtqcLujeL3htyNblXJRhUJzLlq
fHK/u37SjMX091JNQAdJ4kq9Z1bEUpHJ5RvDrYwbkOCy5Ebor4KaNPxPNILQdeCa
OBylTQCWClKAl1NJJxLZKkVMKpdeE/5ZuhoTcfVGRnSkf5aILp6pyTfWubsIUebQ
JSM8lM8RWwHmEAud3ATp5e5mtJC8Ucbwh9e38Mu0lu9oombkWsmMNzOsNSyoRjQA
zQiGcLYNCngO7ryF5wdyfDr+xc1KGg/pZXhtQPPGnTp1hGGtZSZ+YUS2ndFdrOAw
WmMhXPWbUCp5lHsfVJ5PzdzCwN+8rHhxPLxRGUnaqsBuID3IUkpKkqGL2++udxZV
HsckiSlPnhDEph2H9Mnur6E+qyI5mctlsOQV6KOMwoDET7HbHq75imYvcb9JrA2m
qV222yExtc9l+Byyd8RlgioklZZuP0nkQ6ad1DvfEm1nUjaMGOHmj+5xGuiqc720
90V08K6DD4+BFbaUFBauOmyhikP78z4zc+IAGVx5Lm05NrWGttDqIpTw6pWmV/VU
GW2jGLVR+WhfvDVBlcBnqF5bphm83gdqf+ibF8ANJaRJWH77JvPkpNoXHwF+L7dy
DiHGVMrUBuDvCX4+KIJNdmnecuI+LzlWMvS2QD0wWiLpxriNlqGtO3ADEvEHqUND
4dfFu4VVHVsM12cqKzsgACMdysQxSSGHzTMMGqCyXduZr1xmoLk4TTaJ2VbjCERW
QXPokCbtRbthGsJHi/e8EblmYq9y5xfIHMGuSuwxENGKN0tAGLltebs/mZLh8rcn
ZUDnOB0QBG94m1NS+V0ZM8dyAya24nqouVOT+bq09tFUgmleJZ6eS4HxiNQ3Sa9p
r5qCDQ1H7OIqQrTiCGrP40maqzvsNu1FDpyOf1dO9ANIFspwR0QRz6jU1hFBPejT
YxRwmQ+kSXYrJbVef1OGPvK/wRNYB6aZrDdmcy2dV1x4zipaVVZ2gDixwAHfY2lq
bkYKtSUUlKWuVXU6wV/XTLKU+qu/4SraINtNMdCnVy390VAXHCrX0Al6peyR8pCB
tfm25L4Yly5zxUSyOE/bsGXTdd4/zsC6tBeeI3Uh1hu1lsu7DSKXV8Sjdae98rEJ
t2OeRBkM9OqF3+pukdeD9gfPVe/mr88esiNom87KDTvfytpb+cBm/bqnVPAr4QCL
QkLhTAPY2E3GEvdjDdFiozMIEFeh47X0C1cvFCJ6FE0CLCwKEZan7Xk5bHhYO6V8
/lWtzFFSQl6rrhmFEznDBkgqD2MrqMuYBfs5tjuzmfhJATdwrnKSkIu6ILHzrkq3
rBNVeJFmLlTeaFfw5jAP8cKDD9C+R50OsOD4yTn46f++vmHWCwSZEWUWm5iOKJDF
06jshdAoLhnG6X3WeMGk/Y6kDINF0iyHuOiTdEbSwz68WUKQo1Pvt5jw5U7Z5EdQ
OFTFzOtN4lUxM+MXMvi0U+JBHxxWSZfvriuxoVI63ZSVx1jsqGdEdofj7XxIW9fC
MB6apyoLl3DBqzAsw1jT69iP28t5cXIxcC7wTL/rfFZuI97zQrLKVzbLj4le31Ho
w2l+Aa1TCaLy4fH5f2fp05h3xfBNW2vmhRjKZ7VKDjh8Ganeku3qadWeJADdjjUR
GBLLoDOz82obQsAV8fpF8A49SoyFccpq8209iSFR7W/yfn4HWxivSXfZZP5E6ccr
0NpNcGw/deiffLJ2j4ohHfBVAUCGOU5G7QouWAMdz1oNZCqe95WSvT8lQ3xnKypT
vTAgQPhuLGowgIPCp6YAppM58y/j5ZmXgDxasGed0AUkvV8xZU+wAQGN59HDh/rC
q9i8Ru8z8pWced2jSYubzPZ2Vk3kS9hxHJzlG+sdQ76GvmbULB1bzY3pM0tejgXX
j+zYTy5PdTrP0BclwmcBjOXuufpAkas/fCtX12wZAxTa640lnzME7LLwW2ppVr+z
tlfh/b0IbTR86FW7jmQ1CdyU3dLzwNkr307FwdAUfv9eJwD/B4/zlT/YghJ1hQm5
OghKWEcJEQsPTXeyrtJuQxDIQVIXpZjWO0PeceT9Yz3aO9u54DYZeSIBpRNOaUyD
Hclgb8lyS+ESo1d9w7x/w3d2hksU2Zz+zSrVH3cJOR+uXicTkFrSeRwWPLV+qE+E
tV/2i3HMWXSF1wxfiiUE7IsvfsJNpVP703dINGDiaRXGCKf2KWgmpqxwKxwCLEKd
8Etjc0DwLojpi1lw75vtUP/5GVLB63FEtmB6wCi42rRPX+KrZA2C7/gmtLZARShZ
tNPXmdwAvIRig2epka05A3QtHtOoye4hnfKHhwj5WeFscdNV051othnYOFxmSN1V
EdkFdvtJD7ARbJC5Q/bVbB9SgzB8c1/lEQ9AP5fuIkp0y7p3IDD+HLbs+8tm7Y2r
Wk6ekXwudScBh4nFB1Zp5KMRaBW7aLIdEGrp1+fB8ks64drOHEvD2khTehDq1dFo
t8ehRDQsdi2TgQi9ya0Q6UkjvLSD1wMz+HHfaiPizDZ+2ymgFGG42FGmsMHtRTD0
Lmnm0em4Joes0o2PpbT+115nH6LyydFq+xqqEtazJrNTs7KXqCOxJuNlCL+ZAhhU
ONJN6kUF+6BsZ2LHOxBrhMhHzaENg+ERZxZ6bHpP19COSysd5FtNx99GiR/RcWhV
duv3Sm5nlcZF4CPh/2H/4GzAhDMPMxYFijQiuO5rwU0nTd7E7LIX5O802m0cU2Q5
rafoI1aYI8HZWP32GuUVLzHjGTvu0nFp3eLfkL7OsBacNs5N6af21ZhvevcW4Gkt
UtvV78oTYx4ySLYVzQ0LF0MtHWfbLqHLQ6NWekMcsLjz/znX4QbIb5MqgxXIp4e2
0iiCBgjwwksUOW4OhkZNwY2acGodqJKu8V+sa65akq4vsvHcefCnUc/VW4cIaqxu
xaCuchkTZTXhFfBJaqHoj+UJq0D7bwnqi8k4ta/Gmmw9NkAdO4oXFVKBYiy6zIul
poZJp7ffp6o7tsFHQlQAtMHnBywKdZkWL/s16r0CDVKL2oaUC6nBR0Fg0jx2r/Mu
IqnbylPVQEYUGrPd0zHGEAUgEd9rnUK4xIepqmM6Le72nPeBBHeQoDBQJefh5mH4
Wd3CqSUdG4EgcTDI18wMqP7I/XzynnatNkob4vRi9aZaAv+UdziqkjuNDE+bpko5
gFK8OAJmdZMLeJ6i0AyqtwEfjWZsLn49ohbvDPaEm9Jqjtx0wPPVc4rS+0xII3NK
FharAY/DTTib0auBpkyZIA4rv3MpTWwynuhUl7Ndpcjq9YjQXybJYQCXnwCsJsRH
hwBsbBGQi09bcaBxUSzbT1oG0JwQsgsLPpd/ODx8WFqbgDaDuYjI5HRwwiHVavqd
jfc6PR6Qysz0KsmfXe9cIObBIQqvCMx2ry9mw/NJIVsdnfxhWmOZGCfAJzK/fBoN
qlCpI8JXQ5klDi7DCt4SSbl81kubuCpCAx2yaKv8SEFfGEWeXqZHTYWbPF5sCH7i
1m7OIEj9e8KlbdD0diWtzicP3YCV9MXBG5e6aa6f18WLkAWcoxZeSe/Q+d07nNfj
bnT3+V1UqSX9UHKsOAXB2a9zEx1YixTpoMKXpuKg8IFUsgtcMdIpX/QJDBB/Njl3
vlrLq4t2gBLcztfQlaTngUkZnFIfxEn5a9h17MELHu6W9/HJMqMzyUSZ6A9nj3c7
WxH+3FdPNtL6BsRM5w2BoKayzxB9Imw3s/42CiWl+BlTRqGHtDvezb4bonOAut4X
vFIXHKyx1ohNVrEK6NpU+ulIXSjQu5gA6wMzMOaPEBq5eDEBoBimGLpYr52Qm+1l
b7HFYBtp9PPdXviKt64kBvpGzVTH0ePTledNLi5usZJxkd5cfl9/+PsmzN0deVvZ
DKl7tmSRvo6te+41p58xvl3AKI33Wy/p1VWKmYsPW9+TdVhB5gfBL2cexypB3+bf
eX8MLjxRSvaQ+hH8s12TT7Mm4C4BSm1wdTeFp/lBaXGOosqbL4kugT09acJ9g8HW
x6ldgF0tgJ2K0CgxRT/gDmBGley6ztX++oaGnEgPxR9Zp6f1rRihHXwGYDjoelpN
6IwbULPPPQV/2Bk1mfCTGlS0M8IUw3+k0Vc2/qwuWSoJA+j3d8Teay0DRO1cPtB2
NNk0G0f2It+rk05dZ8PIZFYUq80GMewNY6i76OEw2eWbWb0uY94Pw1jn0T5ZxppJ
F0WVLcKCWIYByzZFSQcnEaaw8S6qSzvNS+wPSeNGwAdqd6D80nCH6hgEGLVnEYFK
5ia0nf+TR2Z7+5oU4vUvmrcpg0Ir01/S7/RNIdDQtyOx3EjrYYc1xkMh3z3fOKA0
x3N1imVH4T3watr8zDDbRGYVrEt9FDeIE2ozWDWggySw7GmLAenBSwfx9+ZH99f6
OBsqt3c4SvimbCHNhRgd7LqvLOBlrlUw1UeyK1iCEmGCjaKzYvY9BvGjQ7WAjJvM
HtcsETSrOyOcj8Fa38/o+WMyi43Kva+QlENp2O7ZK9vqy631hs9PHVK/waEnb40k
xaeOwTDG7X1DJSoCRSWBkdbNaMZQwhDc4MLXJ+pC8NNbUAWvunv7wnTXagJBHKit
A/Y80H2Nqrd4t9irZvZVF3FdE23gOR2nb8wNFIbhbnN8w8ZBX00i4V8fWthnyZNA
biaKZKHpuc75MVa/GJJAg4ktEL4BmCnkO4BVCbeNQWlzBae0okz3BYdr0sNBzQzV
11Cx48OuZnoy8wMAQPiYaPh7Wb5sfwUO+VP6th65wKXq/Pymxt1lFe0GI7kbWVH7
1koELlS9KnmF6uQo3j6LecREhNUzULpd5w5PFQUbL31FmOVSiPi8rmdJ08JF7euf
ItKuFCauxK9rJTjindNoaqtksDPRGERJ24sWORDC9wFG46SvwZjmOBIGi/Jl3C3S
kPoCA6wYa6iDPoGawTqJGAhDI4i2hl417VHkBJkurwq6XvkUAelkWZGB/ZENgMnj
1EfCQ2Uwawy27kXFn3p/H41wV0OQvl04veDdo4IM+5BxOVcKj0z28ke3fWkoZnv+
JYErJg4GKoYnhou4XkYKJeY5ji0nQBNJv0G7ey325t/S++IW50QzmJ7KQSINHSUJ
vtAgi4synunKv7caBUMPEn/xqTxZpOYmtqNB5sp/MB/G2ZNN7Uk5qUySmp0RgGJh
tpaHT/nVLhCcDQoAOp0d9aeQtx4lfEYZKBuYwnpy55B+NzQuUd9pMq5F86skoqiX
zwUEEQVT8t9WMxsKaLJYHFLvjRhmfviueL3Q3G7I2rsRNVcdfldPw7zCwgf0kQCY
gQghgyBPII1f/1Q5NHMYdyW2/AXRl1oFPa4hPDOlIrtRtshqGTmbWuv3zMBeBwuZ
OpMJB3hqKvYfHMouqKlqcCERWtPUBsoYNaShJdFrRDRb1WXVJu/s6ljpaBqG0JwG
AjEv5Jc7IvU+5S4aWfAxhq2igVmrTd0fMQwRddbQuoVOfcXQGpAeAowodU8Dd60b
P2kpktiwpRA9xPVazVXymx0Kr4BqbhJKCUrsmZg2awbZQLjRceyxvnEoqbqihb+x
p6hBhdp0h5Qe0zcpLQHwMPBtb9jeXZXmffZ1bU37dTb9mqUAcg8rgAq2ggPcBP2j
Gdi7hpWVxGq0zw3Ht1QHH9kPAtEWthWzh4TPFyxtk0xkTGZ8CCYdGoBhALzJR6IG
ArRY9lePA8qci+Kf64Kn9zwvrUOaVnn9HedvcaBfjG8aszdBoeh6tu0l5OVTEJGA
sccovDv8mOIx9/iXu67Hu4uEpuFbtHNq5pOXKEVi6eo2TOR3np1bI/BRud3uLDWc
HK/dkZp4tRF4gWIvtR33/0WxXWGmfLpHe9zEaX4RrzdTyBghas6pf2H1rR9QVA5/
5YAhreasVXX0XDUA22urot7wt5u6Y4osOtfrd3F0J32uGw9grNLPCTl28DLHm3of
t1vWUO3EbrF9OCN4UfET6IG0L3lcGZ3+r3RbE3Kpug7H99X/xjbPp7bAAuhAzLbf
9kQ1TnE3fMK7kHqErwtWOFjUheNGaQkDe8KnjODTBeNRt3m+SmlQNwpTMNE87Vdf
kIGNJ0NXEqR0+h2o8fzyb6IFtaUfh5iYFQ7kNyk8+VEByOeRAB7KQa7sS0GGRmh7
x6pMPk0P7SKVIDnYMgbHH7pY0jRh/wE65GlWbkvHmSt7H5c7nuq690Q70u17Rpsq
hvPOYvp6XneRR4PA7ubYOt8m4ixD/cdJs1xWQz/HbULwcAyjIuVZmTML0PhuVuyk
8KaGJUEOwngJt3jcPyEUWUj1HXrythrXVVgII9+geHsVcZ9VusliAAaAqbIQMWx7
6vat9rNU1gREqxWz7gO+tYlBXAM7dcyZHpHXYPgTvbvMlDmy90VuTh8LolOwmFW9
ESGEH+K12SElKIqys0qoHc55z1Hg6OqFrGko0ERsRGa6fPzhVUHdA4hQVI/Re/88
KQ7Q4bzK2bgqWBIHqYi0m30xL4ECu84dsTC7cqD26UgSshtzvtq/fKlvBpzjfgDf
phaU28voqg9xdHgS0OGWnYKALQTU0b8H8n2iwYe0gRmnL/SUHlfV+yEdu5+M/oZS
gRhRlBy3kLi6KkrBKQ3bf6WkfgFcJaGMapyYLxxT4LQf508fWlOkUNlWnV5vFsKE
S6lO3hzAUJGqPb50jAFcdzUVX8ukjK75f+iXI+Mqyc4gy0WUMWumFjSOlGyNTEY8
XqtADqW4WBWSoynimhyatZMefeabuMPA+3kBlMagRFK2wG2hEsbJkkec5oD9ztEf
JqGOx9INkFaqTaaymWxsPbQh0VR/0MOGV+7fQDg9tybMl1lbztW69j1r0T+7esXU
bX9qYvjHVH20dbm74rYOKSUKdkbBsUMXzjH2ApxA0VZQJohHbNo5X+d/Nglc3Hw8
T63u7MFFeht1qFFAMNMl2sEBKgA9KTMPqhDj0NzOrjEKAxR1XpEKyaS8n1wZQODt
NY2JqxKF7Q0C3dpX5JRccJRi0dq64aeiN0hBjjYnNkbT3YQNgvT7pw5H54XR+pgY
oOUe53iYJCDJNoWehwvZk8ZijhFtFFy3eowRPzp3Wp8hA0l23lSDywIkPfl3GNYv
FY0ZWrcLGkqRndclaJNE7aIl0KsOX23iem4XxcSbsxZds8Jn1rNKTFrNcZ9qFIqH
rjXgqh6ko9U7uYkBVpN9a/Vq2lxpszse2HyNfMJeLFDAEn5eOxAknf69498e7n5Z
F3dJe3Z3W/nm1J38PkM5SaSuoJTCySaIUr+am5BdwrBXD7D6NzGs/dio1vUNrNjc
c51v1IW4bIgKIyMNwagzPzgEKfYJ6g6VPXABBVqQIzq+Dz8l84taoaAIOKjpcxLQ
q8iRfmzw5HMh3/BrxqQLG7tzawApbArJMhVtky52xFVrybyVTpZe5C+STSJRX4Q9
A9L7GOsEuVCzYHfXfEY8ZCZoxj9MyXxi42Ahpxeyf7jSDsMVZVZyDYpzhHN5dLfN
iG3IH4IeZkzRnMx/ElDt8Nx4+UJzjKHsd67oFcF8UKsIHokQ2YmlrGxvvWlGLWJv
uyTVgm67hHXBHLCJsskLrTCrPnFaxq4FUiJVa8FZqc5I+O4lIeoHL1lXl1Fny0rY
aJDxbhVR3Q6KQZdP9YvG72/HV8y1cejwmm7rv+XEViI=
`pragma protect end_protected
