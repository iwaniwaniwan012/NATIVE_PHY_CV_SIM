`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
G759P1XW9vp4CQQS5M3WZbeYTqdDRTR7z9HZGPi8VDCffi2S3du5LdtIDpH31y1o
oQTCQ/pDFDd3tHvPFO0ioIMtI63gIQOkMpJ3LAaWHqTckVjiLABsxjsyhs1siWZZ
THsrdGj4mm92YoXFXoaG1R/Q8DUwfTaSDQHTst21bh0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22160)
iZ8tjAoqNDhnv2IS+mc2NKpC/XPQS9B8qYbzuu9Eg1mWZPQO3jvIbfR+XRfA8PuW
Cn63J39ShvI0KuMksf0h5X8r7u43XDwHQJW86yUj2MdtmhKBDSFOLRcD1LZQRlVY
96YuNhbzgqOX9drlq8xNy/rRzejshby8P4n5vDjIDOdhe2nS5HnHKU5UpsFzGPT4
sfEsZcrd75UraElozp9+zbgAyaPiHzmyO77690XI1pj9V0YSDOsY1u6hTaxVhc3V
uKXkTMOXNH6yzIlpM9vyE61QHexczTfv42DHyQxjtCac7JKL+eoi5CMlwTAmQmlq
SFqsoiugPsilydXrU7SRqR5ZnKW95KfYZ1RP3VGrugqXqMUnSbznJgxp/E1nsQL3
Za5OhAGcxldbl8mm6Pa37rB3UE8+lnKOenpCekNqwrFBzmIM5sYEBZalyyy/Bh7/
QksLpTzUBg08wuJ/XdnbcyykudhXc5vMg6Pw8vLAAdYh+V0aZ9jlI1PgWLp7u9ND
OdeulO/JhgUwKlH6T76Y5Gmq2BBeqCxOJpFTft4wowHRE0Sg2fCfrMOd4cbqRNq5
1Tfemk3/BNvmS+JcdDdD9hhMrX/660wOWzXlnhAab5u8/DIJSgQejvG4mvAo5IRR
rkvbr2n3Rs4QEjp27n+bD3iKlcjN+iiRvXIvS3R4XYK9Jbvwj9ZYFFLaRBO5tLph
8YXlBqbyDxroZpsn3JQdNSYOA9PPWXKop0a1Ck96eaT3QdAgwn4rwQfdjIiJbkw4
QYZ7bNQfHdjzhhUusL22QoTaCw9RtuoGZwO2VLROk9co+bFvlVYVD5DeIMf2Qrtv
9KJfmBl4CdkyvkUuoEC1NHiFr6F2cL9mpmMN1kb9oNVSxgs55pdWjI9TxcuV80xk
obPX3LNJ49K7psL2UqqUhULMjQ05X4pLKbFtwvZVf9o7GZkZAHGeuj9tbZ64jMOE
yDJM3xIN4HiifrKtEKFOg9NQoMagLy27S/pr4PbD8I7M4DCmESXFdGtrRUnGscB7
yr6RIfuemlts2sD/LVXWSP4KdlpndOpfk4tpANXqymHAInLh6OS94hAPUOfAn53u
xysWEmKV1MImPp82pq/yM54PrOGckWSr/BRCl4JKd/CVdT/aw3c6ouzQLWKm0ifF
QWXuipOXKSupWD+ad5V3Rtszup2wAQPJWMHGMdV8DF8T+q5n/f2QoF/dvKuWu3cH
z5SUZVGjJC0vzIGnIvHtDOxiR7529t5ctoSQmzhmQsEtRtAJWcII7PPwErp90VBV
FlzmHQwS+Pc30uQool1nsO63kpBRZfGx0dOgNceTigsMaTlQpADfs8EHBtDV6I4o
Mo2BLLHAwAPWIZmx9Q+vTH9cJ7ZtSYve9bmZku9FfGUbs8BcWLRI2J99fIGbNyjn
40n1+4p7WV/M+PKc89OilEklgecaR+wpWfO5OpWqRvmMlDxHI6bgyI6FBMgARDmS
7PIINwx3xGhQwHOeg7qNX1wuj0ofZvXGlqRF4z9HTkoh9gmq2T9g5zrO0Q5yRV30
10VGV7NEDEgnnFClpkKccxbRbsNuQzDvC7ozphqCTwXZJ0QBMYSz8QAAUUIS8Yon
6I7LSLCKz0+bDfLyfwUgiWoGtMjTXVuaY9PkXfCU4lBIJZJThSjCAIuB0i0ATFNT
OjWZq0JDINh7sj0XjJmmHTtKsidcE37mQ3SCtHFka3mDOPbglP3VB9pljWrKUF+q
KSHuU5xobrdZZ4VygYScE9oLms9LZPaHSl6sxyb2DXeZdcIKPqeQKicIQ9xxbbK9
5pBK9UKCbZ9rbRAGpFcqJzLl1KL6QcW11zWMQdLoOzGjzzY6+bfnPpZOCk4SRqH4
yxiNbQB9tbavxNe3YxOXRUiZgIyJltd9+KrYkxg9PPHpBHEAntBI3uCd0mANBRng
kWvNxgr6FlZ6tBLEYNgVB4zMXJGtXaThKnyiowlnDeEzeQiF8RH6A4gKxovUtDWQ
51ymTojkhT9WaNpurNYa9aHwKHGROz6gs6DqC51BCsJwRo2d0PLJjY4IQpX224zP
MgwjuAq/k5gtdRkuIVzpFV1MZ17k855h5p4NQ0j7f/hhc0Pws2rhukvwNpdoWa1U
qyCheyeaRhl+o0gYM6QAvaj+Ha6mgG49ZfLit9SO+1+MpwZccKOO0Rru2+VYzurF
AFaqHGb8uUCwM29Z2/xip2g/2ye6HwhmvLHD6OiksUYBdDyLtjYindD8r5YIakOE
aD3cYupmPjUxi/mye9QXPCk90R7oX4hINBuD93KQvhzpPRqOwoOa7/iwgjr3SzzB
I+pMZBfpv3IA9DFHgoo1+jZ2+s4RKUljOhTIfeimW9JKCu1hXFmRp1+rR1Ca0W2Q
fD9KfDs/wKslrV79Z/aFbI/HkQek1PrsxSzpRDI3sA3XocHmjHZAvvi6dxLKajwI
qU5JdxH/L6wiMyOU2BipNqDM8Y4C5h8eOAZrRARw8aRcZteSPERkMDzfPJPYg5E/
ngbME4O840dAXSU34ALnn0D9ygFruJztHl0ksuX69m5EHbiuGz2G+gdgsWF6O+Uu
IW0PxEedOmnBB6Y76JB4nrehnfL+pOt2AK3tDlINkFZqsHA1TqOftYU4yeu6Mkmm
veWQl03mBYOQOVYFzJo/ElkBy1etAabWoUMu7Mk2vI8TzJdxAlpD95N3qMJZSt5U
BOf0r9DlC5oDZxgcg4ViW6EJXpZN1RSH5NjLibBcHeTtuS1upFGY0jnwkTm1bLLV
fQ0XZo1/+7hU1Vc1hwGzaraik30M/Jlwo+ZtD18sUqz2W4hv9xcaXzPeCu5gjm2M
BZSPQYBC5PGN9+4CpFjiYqHmRBGfRClqbY5KlAsksfhyGycRh+O4GCrozmK54BiS
Z7Z3LnJ+2y4aQsLvr69H3KegqZcxrQ7XCysTSer8/ux7Xh7H1iqc9y2oxwvoaEGP
T6T6Z1VZqHlHLaBGYexJf2lwZOEe/FLzHOWFPb7YfRYAQSfJuAGpy7Xjh7qGKfoY
y2sQN5kaRqozzBIbXRNmNs5xfRRzwGYysLMgL9pcgoi5baz9e2C3J1s2TmjvUozU
tnRgRTDZvXzcibMvjGROL1zC6ThE3UI3mYGBs+OW2lSPJ1idEi+5lcmiMnc8zpxo
7uecyy6wgZN1Hdvyt2+p+2C1F5wE9Sh0q+ui9ikIAdHshPhyQ43wqPWD8tgjJ/ZF
Y8/aJPvdfEbF96gt2rkrmL1nNkXcTtQi6cXehxUHrd6QIWXTdsX1eAUTRQFbDMOq
pymUH0mNWjFnHw67eeHU9MNZu+GW5WXnGoy588llr7lbkkDEqHfA/OwNzogeE2hn
IC9c6Coir66sw1A0SR9Ea3F7uf/TehsJXdDUeBFGqYaAdS1VICDRtsbXdoZ5IhYA
9tN0xpaTeYPiyufKjpajPU0RtnKzLBIyi/BAJwcSww4HdxYxNABuAerddzH6fDWw
23k7v5tay6bfwVoB8Z3rPt4noI/J6yjQ2SGYz2O/7yoi28UG+K6sc61xyAb8LJ3S
MgVJmT5zkiTH6FfPkg7vAyrxcdiB4TP8viLWeTZC/AosmlCfbWJ3HjYnpCNVbWnY
WkbcY0KwOFVBXP9sg19G4Zj3OYZAiZIYBNieru6pZLxcko5WOjb9IfNU3TBseqbM
7d2faIjA9nxcFISeyd4rRyWviTtfptwggkRdqAwu4NDJSNKac4lCX8MfQHcjBC/g
D9hwiRNHo0JGAbN4Y4Yt1yuxIqF2DnSKYLt4q2GbXmRbga12vQkTPsvV6dNo7r+l
KI+lv39u/16Jhl6ZZPwhHdCxkjPEUWdB3Hw3Aabw9tk9nGPGoIWXygUke3jjGHWe
FFY87zcbW6+cKYCUwzjlXqEnxOqVcfcUCABg/SEuDHJRERYJEIlAmenU062YrCm4
vIp3LvjvB+YbpiBEE8r7VJy1ffoRwdAs2dnwGayXyxZe2SJhoMtXqpB0168ws3A7
9lD8Ke8IjIu3r7aeQrJ7HFqGpNzj4ENFhviMHakGlINx5S+q6MbnChtyfg71tY1T
HQqIH9P+QjhT3XGaymIOdl6IYpw51Qy3CkKgQ7A+wW1oEYHqhIPGveGk3UAig0f6
O2BHCmMAYbGBWb8XfWdwVqRgr5hrloqEztbEEgqIBckJI4eSvGTG40QCHjs6Veo8
jLEwKrOQeh3aUsmN4GLnSXWRRLY8qhBZvcGzO0UMvenxsTM8dG+xKwtzNQAVPCkD
VjKs0B+Ld2D2z85pzEeH4VEqghCsUJ/aSciMn0OMQn6LbV3hlXOM7+AsMA3G+WVR
OG3ZBjWW75De14KKT6N7ux0cBUN7EdU543xPNIpvWo5b9cIz3ez1mk3yKQfHEBxJ
76Z7fNLG0uAwmXIbVI+lgj/BXHDdSEqW+8pbMka/gjiYVVhOO6g5EVFRzV1cstEC
ydgDSkpqaZ+wK4LlCTX5e+n8YCr7fSTVDEcZtdkgzuMlIhRyTlC+K+1idq5qdu4B
pQO1u70k+D16h/psT9EExmU2zYsEiOBwC1rK5LPYP4+tnYJJVRORPPXEsXey8m1d
noQzQ6FXhzaQgwOj6taZyyfZw/Gjq1yqOK1mnrgwCKid9MVeXBZ7YvuGVF7cRXnf
x+T3YtvWl22XVohS6g1/u7z8QPbs8YeHwnPdtg6apYP3gr/exRF9b2O11eqcdYh7
mIA7t5h3fmgIqoDSA0+VyIJX1YptiVXKYo6ax1v6fHeBirvSsd++8gJNBu4ioGH3
8LXIlDksTZ52jnAusqvYpeDhl3qMNrW2KQvtuTcFLSYcgRf6LfWRYPNZb9R0pFwy
doUN/MiyRnMuNPS6DXuPR7UuF/G1V5Ktn5j3jA28l0IE5/dOyLch4Vj6FGJbX1px
ps1IsvZ8RnoRNVfbEy1Pi8ihY+cUHE6Xr/u6QKFc+Qf4B3xhrJCPk8z3TEpG+RSM
DS1+3/Rj5ZPfyECOQBbkVPQhQE9LYjuifKIMJP7z5F+eH967nxsSTGDAXMFyqP0c
8Y2dhBGIZynXLVo612qHSC5w13eeVAbxxSQfk5mejxggChRTJgQz0o8ngoA2j1Us
9TD3lbIOxyrxl5UynBSaF6/N/LKdX/w4rr7ZNshZTPhsMRz8+KJemulD36s+Duud
JU/QELHAj58MlaojxdKTbywl566a2R36+nU1OpRnfEkmnmFM9BR7Yyxe/+7bu2Ec
MvZXYNxpeF6+3K1BX+8lPSUINm4KTg1S46NI79bSEtOya5oOLtaWE0E47Y8g3C3h
+M4pFjv0ozA2UdjyXGPrp1qiFBojQsqNzOddRIZyqUKz6e7bnr0VotzNVsrERyMw
jY2xNbnunehGm896+b9IPLlwlH0Q0NJTnm953SflPjrGwnnbZxOLSlFoP/B9mhNM
+DhkGnUtB9ZtUQwYAtDr7JR4kci/WQhic6nV0ur3xAmMqDwJ9bJ4pdoqWKt4MP8I
AKff/MAVObOxP1cbpslnv5OoHR70PeAIVpY2lAbxXtGd0ZupRPVi/uYTCMr6JYl8
O77F9BOhtx1q1ZhWPMFMcGgFbV/jT53RPPpgm4XSyXaiaMibflRWETyo+1evPs8Q
BVocbjU5iowlrVmANsEGWkodQanUehAOeSlKsDfIljo7cdjbI37hk/SU/2+lfcuX
0h5/vOBFeGv3CV6fBgC0ZsnD/Et3h3OgpZefwaWTdR5L8Th8kbzqHxgluV0dYasY
ZwjNqetzL86M2qnQxiSrXrK6rg/3B2I7UxKmHaeH/NVQJ9/PCgkS5avx5EPKnEZB
UFtR0neGsECFESLFBRo24nbvEGWV5TfcZpoZEArR8z1Y6wVuTPygxEA3LSQMTHxO
xTXDwImNvKVutVrR5PQGdICA++2Rp5LpOkDYPXgeXi2ZnPeAbLGYonAfqTYQXHsA
n5mSXnJ702qq9OdiBza91fU0z2zeXfMd9n+EPo+cpBnQ3S8iq2dRCMj9EMkHn460
24Tsi+tswmsYR22uMDRoz3gvbavJSR6IN2HJRSpGSt1OWQy/PcbGr1K3rYzrRIZN
eURnRBao3fyeL7Wrvjyc9L3GXgN0ofdJdJYVk9xYt2VG3IrTNiSlj52nZhVtGP5I
aXV0VoHLDHCWt0JOsgQxqncnc7zaK3g1kjsfi79cZKe2JXNwVrBkk3bjT1D62ron
SNNLWnYCztWcJjR7Hq1FJQo37ohNseSB2PT4WPBcQrA0PSviEhOX67iZ38Gh03/U
BMmaWOj80TgZPl44Jb1mNhcSzTE7lklZraf1ewGmrtpaW5/6kpaNgPsowyzFKx/D
UUQZxl7atwYbhJi9UL4prFYHTRfB40yQkiZeo6DuPpWK+tsHvXMrAvH2DsLrCIlh
2QWiplTJYrARtlA0FsWFI5Hb5+4CnznMQJG8OH4L1KkS7djoYrDaTEvWtQjVgl2M
C6xQKxcJ0xxKYmEWtiymHcefUNY+d/0kCO8wgUNYrBui+SD8TVA+jJl7NsH4IwDM
eohvw0KMh8Ga6jBiI0CryL8231swGGpjGE1XjZgcc5V6ectKC9bQ9h5fpmHF2nMu
i+BqDsj7EsT/dsb7lHR53V4hyL/dUkjm23kDeZKmWizJstoje1iwVFbi8okCP/N0
Culm90c0fL3Jxh76Je2amttQfFZ/iwrChfaMR1LBAGCN47QoclsjCacm17mkMWV/
gFoAsmHVD0KLuVjdFRxyQkr5fQxpbUCBETPXMzhjwIwrKBHVjmXmaldztJhnCZbY
YtIINvDyk3U4H7vaixi7j6c52D/4oQ9Gf4Rmwn/G+iq3XAJxgCrg6UrrJe9oRnOj
G8fOtU6sMSmXX65LsjeOhzqcSXmK7Q/FW18oI6WH68qmGajRG4n7cqVao26JmG+b
pBA+8hF+hGvx39oc/EGzsNVTF6Usmn/kZBgJxoNXDxEjpXQAfKDiOeqMBcV7xD1+
Y8mXt5xezeIZ02PjZOF2SAjt8b6u2YY49pqyMYU8vZC+dF4vrSm1hDIMS9EV8IGi
ZJp9pSQPGq89mqr53xFD0x+EJmGZzBKhCZAjkOXFLpQyfAZ+zWAimQJVQB9R2x40
UvBild1RCrW4nhp1GueO4ZxR4y2LHau+2FGwsDFxR1bL3OexlXfF271QbNdaDhEQ
AEQ1mhX+ow8mpvfTatKW816tz/irDlnvNO/UI0uXAX4zHsXcqQSIm2Z5DaEL5zX0
iOfy7k30g6Jy+eR535TCVzFBLtYXGPkkzCAE8pbOQI/oU1roMvNqSdvmIesblbVu
iso2MWplffDDmk+U85gha3uPToAOR8nEbpNffv1YuqPU7o/f02+LBWA1tilgn7O7
taGaKa/E0PVFlKmG66XnSEEJ1yf/QYZ1CvXXKpu0CebUxoo9jP5x6yegpRMh87ng
YaKVf/8Zqc27oDpqnxg05Ju87YMwfBdofhl2WC3bYv6XhF52/SFzpA4giOXY3Aa9
iCtzLt+tGVILr855ePBz9RLRXgJvvZewPwESG5UF/xaA1p802fc1NQhmbQsmgq/R
0YJktrvVOTV/MY5+RQCAJ3U4NFjTVmH571UddlbsvKU0vms8xjF6yZuvgRVFe32Q
VwzmhRl5djl57JlZTfLGSqLjZmDxhte1qefgOjB9+LRLy60ePok78bPcZ88cJmPH
iSqskcMAszBJvwRNa92D/V4qPDEUs4IF62fArikR3WX9f/hw/BA9lpcm0v1WH220
QCkNJpVoyf5gaZgSQo3kVcJqCEXgMc3oHI0lSI7D07Q88gJEg+3qn6iLtLO8NqiX
4sCzIkK89LwitKzmS75b77JQLr7QK/UmwBQp2PgdH/5hwOF7UN6lv9AC9ECUl2mW
DPxqBJ40xQUCcTG5Kp3typtwVG+slDAr/KG8yliZnJCOExmtFNdfD6p3ohn1MBez
UO+neiUCKe1TXZiGy0YnKwzZxCkH4Ys1UMX0Mmsop30FipzR1RstMoQLlwpdcaXE
0HOAm0azKq5vg13aWkY9BNUhh/y74esK6Bb1bec63thMvjt6dnFNuHP73sa5zAx0
km15ASd03obf+XLoS3lJT7vw9fw4DaQRrNWVYhFtvl2ST0hZE9lEK/7XJv+i9xcZ
+ypPhaRjfy+m/2Pot+vAmzspkoeWEwC1YgWqvqihG/Aix1vY7GFr5O8WzriiXY7e
ewRvJt0k2TW+OADbnlaWIGgjZBY4oSV/iw7IifCjKhPm/EX1O8DWEhk4KPH221IS
gSXiL8L5UCdt/A8nNiCTUHRp8x1g3OhNXQ9g9WqN0MtyYpdfNlL7nLHUf5QYgBq0
xNjN43INGYlHQB+bJp2xC2PQtEb49W3B76rIyBhheQAbWDlsGcnUQiPZj1e9Ufeo
Iy4ZHVEPgFOZlzLCmK6u05R98CAyQpHF1SHulOHy7Fndy2KCJ8F3tOrDwZKfpFAY
XOoiiE3nu8ZKQaVmCjYn5Ojg3qv5z8pMad4nV6JReIlEEMXSHEBMOWcWtVaTotBk
vhmPz9vxADZswIYCX0YaE9+LakMOELilZKJRxP82OAN67WKoEwVjt+R97isWkqws
CUg7+nHZiM5wYls2RKqEyKtOQ2y7eyYt2OnK1f2j847dPIZdNN262lCQZ+PK/SZO
LTI5A4t34/1ZtZiI8hySwWBbcuqiDhN8I/Onq2Wlz8UVCQ0iDd/1CuoIzSLUc8bz
+hmT7ZoMhLgxT1YLMxwZcQHgglKtsfpD+fumVSf5vGHMtnPJ8To076kw9HNQkVKQ
evrlSSwc21dTfwIVdz4NrVGM+dhGGcc8ZOliOjPhZgAAiaVm3eA5q/fUBZaqE25l
qu77hHOs8vWUA9bMjKGkWp2CEamRYwGen6V1SRhKYIi7lMZQ5WzC0rptEp5eFY7j
MX6oMstS/HcK1NtWuKmxbMMUT2op/tajfunuk74CAn1oT56bmL/7UoKY+LLQ9mHr
46XKn1XAQsJA78+CdthJ4wUhcCYVCeBYy2f3m6YKQE+zzRnNIAhbgA7urPLIxekp
0txKnb00CcEPQiLm12c1CMAspO/KWCz18TQbM4jvyIAm/qB6qJmQ5hjBP9WEotWi
PlYGNGxs71x2+uF22KYrXbm84kIp7NRtkpERzrL2y1c8wU2hrMjJud5lK0OKzzUt
SrYmvKtLi3dzNF+TrPqabWBKVa+r0yBqQ/O+iZQhAayEgSsiGlRfoOCwRJVbCVMy
RmyiDXoH09/SDt7WYtmFtjV6bXmVb6nVRdQ29IHj6SelKgTg0y86iADaeSCu/a+8
9LfCkiZFXZ+GBJOOpOaM9AuGUFivtddW/i89yGsBm9kAz6mzPdqXiPS7HwjgpjxK
VfFVfh3ls8h/vj4B0oPbCQF15sEJrQlPzBG7T6tAJNzu3GAI46sG0MvmEqZQdghH
BKH0TM4ISDLJYu3LXth7xRNdpsoVIMBvy4oiCcg9ks5P7YVVEEgvPHb7jwHYBukC
Q1OLmEoxDht6ROVRiORK/1Tp98biFyklDRP3jnsIQ/xWcIfnNoR7vAj41q4PK9v6
KUMKCpklwit9CqzL3mtKWqk/XxpSyOIH/nJpAf7FIGfCRDAa9kazRzWE7Vu+RajW
I7iJ2xib+sVf2kiY4VVz6LYAiUteg3ARARfEEAmdHc5dqqmvqN+B4LZeczswfzgd
tWx4gF77aMMXGRxyJYIgrrIf7Ke+tib+ilDWOCE7/ZHf9NCbNiET79xUHfZReWjf
Xf1TBo022ikxUXb0g4EWTn/N8+VzXCofGHQMlpPHCKUqb9DZd3T01gaV0b3Y8BIM
e61gdcBkUfFTtu/Hi0yf1uuKPfHH3wG1+KdMiV5q/yP//7dSbsx4DOeqHorsW47S
LV6dMaLaHhOSc9vBRls3ZGHdxh244A4//lKCHbV3a1b97c0hAT2juWtPtZ8UCu0Q
OoiQ5fyrtkPMyPv33h6/d4sy0ExHYrR5LCP2FZ1jlpELqp3oVr6D9zig5DRS5ESk
ErkQM/mOOug+dUXC3buwH3/dkNE5hHgcZwkbbRrHFw53OC1lecOdI26Ehti43m1n
QTZ9d+5bSgQkdBLWRn8uKkcHBLX1+p80mJuSrahQhXPLuszTxfk7KWn3Hm+j2VKn
hsyN+/u+yZDNEoei7Yr2rzWpRFxR+1ldYASitVro/4ke3Mf3nlVeKkXIacFuk6+m
cKSOisme0v2WlSR3psVNE7Pukob+aWZznprC6bs5KJB6iXXf3sR7fw4ANwfNkA7h
RLlpYDdFo0y+HJT5pFLaHnVkSZtqlxR9Rp12vahhFzmdmKfsYImv+V5CtBKEHfKw
g9CI6BYdZcfpQQ1r9v2NNEWty9Lc6lMet3SKlFxZWgRbD/TQ7mGr/Wsfkq/K06u3
UaTKrt485rdGvgsIkQJySTJMn5F2PctNmuGKCc+QiGdnXttlSpkmFDNKJiB5FCZT
LG7xVJe86lA6/Erueci8P/xc2rKDWuTQEygJP/zQtm2f2Oo7E8B9xMbvp1jWy3Mp
o1J2BrSsq35YvcigLzi3cinO3uVWi2UeGwUYD0c8q5M3PEzMjj9ojLuXZWeWXvta
eVUFwYeT3YgwzCw+cllqNP3P9ju3CRGlEkRNEmJsnTCx6kCoHI8XuuFz7Q1FDWry
0lcawz8RQpjAin972naj15duwVrGZCrIF4ig6Ddw2os+/rv1R6z1Na5iKNvacBhA
ZRs/sLO9M3kEXYOJCTffN98A7Dd+82O/1OxyeYaN6JvSylx7Q+IhSfQKf2Q4lRVU
BCEeU7TgPQevwpBiYiCDFwOVwp6Z4mtj7Om8c/c7LtCypht5cAGlTCDrHa5Yzbm5
VNEsh/pCEcsg1HYprC8N22EtuKKnxADHp+p+8lEYb3S8opj56AN9QBz3t6CSOdSS
DY/9tr8Zqegci6kgALUm+m88Cg+8B4T6JCXADbQuq4CayJ8YukdJnMwTgZEDtnh0
drk4582xBd2DldnnXjEDADy3e5/HwPaV3FR6gjZ+KITiz2KMRNfLwp+c4XHNr1N6
vFjJakUvVQSRWTTqaltz/P0AG8YVXwk1AD94OF3Qfh9eyiTt4LfLqwRuco99mTmY
5TqOOGtCThxYTkrUOPItMtQ4A07FweG8M+3l1iLXRtDN6kYIa7cVDZZ9JA/xXufX
Kq9dlG4AICbOOCCkB+i0ZuejDUe8xIUZLOYyJwxboSV967MhHTi9O10W9XvRKhuY
+BFvVDIVzlZUZx6Yy6CF2/Jf8NtpVujvmWkC4bRp9GRGLzn6Lgie1S9Zawxo+V3n
/mMImWhot65Mbht4kT/xBNIujbIEWr9wBDeueGf1yFZlyPTGy25KZX152ruMdqwJ
UCA3Ghvl7GM0CAnAdGjXprK6d7Cgrh6LNQCYrs8KTwsp3SmOlTMqwJhmeRd8xHvz
EmF/IHH/oVSNCeNJIHtnZZKgZy84tZhGd5C2/YBaR9MvgcpJEdRPVKXRHeh6mag8
WEGgRwVBV+OkmfP5FNf5iculAo4OoObIIHiZ4peu7c9IaoqaJPxzRs6hF8/0RsvO
WP4VRmy/exnycrWLFnyN2JlPm7BERAQpTftcoDp+nKi0nhEs0Ie0ymokgflSQNaO
dNIgApf9hnDmERLbXlbatR5o6F99mcNrxbwc1wkvVpnEW+mT5yjRwGVRuG5HlXVU
wzTcFQUUmrGhYB5UxJmEw1O4FxuIUokjpMelCCJGFIolfH3FGGYo9+T59ohbfYhB
JPnUHOVxVHmLlw+8NYCgqiPOIGJAjj/GC7YpQN6JWTkTaIlazL2v8BPWxHSPmPoN
OCYsYuTpVHYsQSuQPdjjaMpef9+4EENLN7HY1iw6Phsdv6OTtjolyVb2V+rfwx57
FiBLms+3uX2EAua5S692oj3+tqPD0LSUU3Bf1uSbfL98kShnyHqXq7w3izS1/KUS
BkxAswgXgelM4hYVFVGbsJpW3qMCESTNsOzwMhywQkdwOCskVXF/nVl4cmCc4VR2
ai1LWijXlDk+SbI12vLsMQgFxHOB5X4TXgoeEIAQnUGuyvJuo6HsrV66pK2t2zaR
k561lr88M7jZVAqinqI5O8LWbi6kzriTofKo0Pz/Z9EYWtt7MUtXadwoldfygl5L
HWDDxUL9gBDPjSDAS5LikHqxsMM1rC02GTHpRcOzLGfVQHu+11xA5NX2+5xDdc+w
uUlp13dl7uCqWzrxjn6eelbqLs2u0Dd+cBRNLqzV1NSLw2rpieT4cPnSyde1QnPv
wA16929JXjfXP6+ii2jjPlPxZO8FCOjRF2arsfa6PdEGn99tDIMp7GWdxbSaLWMa
nnMeRkiEGpA1/p16cbKpdc6c7CWowZu7sDl5MPi2MKtvPNidTV71Aj0LgtU8gMSe
RxEBn/Z5/P6Lb6rG/L/EJ9yBsHyKflnGXW2SR5kEDTrKeDONUKFn+oajp+g9o0CE
/LbW3cHpExgAa0OrcnQF1fNCfKDiUPuQyACM83MLQkN80wL1FxOB/xuZpd8UU71y
VMOzfxdzsgR30JUwagkQ+HPMMGq4jH97Bwe/X7DHn9BW9f2xf3Tf53gnUBgPKpu8
7Zh3nUERqZxCoLfMGrZEu7uIC0tcFMK5pvlShHA5t5fyRZOKYVRyhuY+KMruUA48
Ibt6pE+vYLcDz3WKEo0Or1GVIuUZYQLKb2BfMogJfh8VJoOHFizvOX31ENngmed4
J9Ky8s+mfGTZ/rUafFkgHwOFq9bNy1GGc7ydsmzfMPpDaUULrqgNAtWziXxFwwHd
Q9QbyQxa1vtx9FfXDBb9rCozqRiuKiotz8/yCiM8tTYiLXL+1ZyJUVIV8+hnTi1V
iGDOEKfH2OI5T+mRzllc8gI1LQXA/a7df/YFk2mb7rrfZiECUbjoduyej6PjblPX
ozyU6m7tNs+gCIvcorSX/3lvOhfa6a8SlED3WPia9D0gGWcbIAWrfNOaKQBSiMcU
+iDmbA/RfO8L6z1XESkEIsYroISsvq350vnTQkwtqGYK+zeq8KqHZI/KQrhNUJ/3
O4GUE4Jxn3MiCNNdrls62sCwWIRg9m7C9MMmrQJ22e2E/WpagswGQDext+L/XAnO
UTS8J4tDdaGoXkiQ9h7mJaIfusZDBljNi7BOcqhEgYLm5HjnStKheZ6KEuxmFg5X
bpON/WyjmjwLLjvydt72/L+wuD4W2Pa8ldQeiXmPL/JXPFZjyFLzZTQeJ9zwLIoI
orlaJHV99qUEMhJyNjbx+NURKAIFM96b2YPXaFSL1X5wLjad6fNGRt/Fi0/oTrG2
RPDc1Iawq4IGUYq28dOIx/7cJ1Bj2xck2EciIANLPg4HJBHo0j/LEDSc8vMwzBKj
e8sdIPjDAGFaacT3AH6H+hE8cL4JzVZK3LQJPyh3z8ENZK+kxBlWQcifA3gmR35D
3joTFyLGojupzoy+avDo5uGFpOcQo52Cbs5hKbs4B8zKwAiHKhidbfCEaHkQjgn5
g0DfVRTxqyN+i+traZ2+oR7Nu/E2uzHMkkAyuT2QMKcGV8zGWsl8PZKD6xs4ATn9
X8kSi4j+hV4mIHHoVW2OP4AmfIZKGDX7UK3HXuOWsLX7N2Mq965OR3aV97Ss4IWQ
oYYrGVsju0lBWRJxwiPwbZJtW+lznEC9GT7MZ1jIUJ4G9Ktr9KylGPd9Cs7uxn74
s/6KWuzdeFZ8B16LJ3XhAkOXYGFcJVhGZAPh7BJaLQKVhyL4FJvHKlmY+gpuogn3
4WA488Y9S+b5eAqP2pcQkUSnFQUz2qy647++Xix9CWCxSdKPpj6oy2EYR43TkIFG
4k0MHUBRgBy8xqdNck8F3l8ClfQ1/QzqT2s3TJuea5a5aqWQ8i1C01LLVju9o5Rj
Yj8c/eFU2yCkg6q34sSm2OpH8hSKl04KJlKqQeMDXj6TaldwvTKrpyt7Q1aloRuk
FNl1tLTQ2XoP67uBljVsws02lGn4mg12MohfVGLsjvoQR8yEl2we4fnGtu5/wgm1
y2g8ngZGbyVJ3Xm8bpDMYs0bUzVS7AeN8TjySBhGmEiO6P7cBSJBInxRD9m0uAPb
aJ6IzbjFOmKYUQk7c1WBwrfAEI1YZmHw/cZyqAUaepmxSf3ACs/Fl3SxU+UZ2OgR
aFg8TfgwEPy8mzqjGp61/0MDW9o5dcyqdnJzJ5mpWE+ctSwtGLNwZlCHl5C5nscM
MaLQkD43hCQObv4cpI8UtWpoz9NYA3egCnoeadY8xbJIbk8+zs/2K7Y8ksIpSbrd
DL36d3YoSs/OgWeZd7jYuIoBWStlnioCe8d/LdOqr518eiPGJHZSkljgM1WRNwWg
eimILZ6zsAwS/qCtSH0pM9kXUwGu/7DscBhOcDYApMDR8bz4Y4BzfVwwv9rWNEGZ
Ru9uedu/YscP4BYl6nwHeXBGOcbV+17nfAOlcHngE8X9B8QEUjKLzzXFP6SCPZm0
hBoLnOG32OWijv/qrwHYSHSkGquSVTtyMkcdP7IKGLDVcxPZcDRDtXhmMowbjiwM
kdBQ9Yi4hM3D3wEkktlOROwIkVD44woNuG93TnC1K7s2qbxpZQCiA05LyGXrrdwE
V1UMfDHKA1huSMxLR/fpfXPxVAbsfUExa2wE439oRMC5iP3R/7ipgHEFjgNI12Z0
RQwDvqMzMkiD8DjvQYC2mL2IJirzH+BoJUaxn85UF6FNsg5w+IBg7H0L51vhIcYk
nj6FounKyfuAk/ZckJ3AWX9eV700HLE4/lyxf87D9RYqiVM/q1DIRy+gCuSumr1F
6XCtpmqUUsxH7YiTYVxPu1tUPK0B8utg1GHJm1wy2Wv2HYF71k+xBxENKXG1Ip8i
Y8cJZcJT/6908HA84Xu7EeYDDiV9SupFKpqmFpGDyB75hj7t513JMx0Y/tTsZ+Nk
DWWjS7HnxwGuq5qidO+JHrfYmFf4vEjIg459r0VncRvSAdSgCw7VxWhL6m1flQ+X
O5sRO83AVT0OrpBmQ4SZ9h5xqapDYC3OiTop330SWn/Dn/wJ9uVaDkAHJb0YURxs
0Jyz5wtlkELd/TKNGDMPuaop//2KxuVs532tWc/gkXCz9PvtAqqdfTUrArd46IrV
QYb8KytzAgnjZDc2xs0cAiBSFyBBNHJwvtoKudv18Fi6wd0tRxuBbnyHbfWXE30V
jlqq92NjAOwCe9oNi8ug45+6wj2aUNgl0SKoCdTU73joOo70RdXHxd8PKgJykiKM
6iQ49vEfU4vz1xLmPsRP2Xq7GGz/4qCbHacEONXjSSCS1Gy7A6fW9wX5c9W82+uS
i4D+vHb2eFGM8A6DjShPk52UUOVhI4rxDZK+XMCnvVmxzGKyPBMbxcjKAVlqlNsp
cthRg18AWh4dVZdHfO0XTbVmRiCFYOCbmMI3u/wUvObI4Qp29f+T2HpddswQoXQf
GME4eOKqTga89hzv62Y7j/G42M6sunoVscZEtSA34OFsnDyCe72D0+iYs2Y8IOn0
wVwdGwq+f6xToflJh3lpTeSQZU2llmPt9NMnYIyLBQcTjL2wayhKXuf54pMfF9PM
+1DJ/wwSg52D/r33392aP2trCiiZ2WHZPHU6c5kNc5bnTqG8E8bklMdPbI4mKKu9
H/nCRZO2FoopoxRr1HP/rhHED4hMKB4HE8+Ojpv74qIJdrI2IIpzifIowh9YDcIT
GA2IrOhtnywScTXN/gChGgRWlnywgIsHtT1+GRNXC4j8CcMAd/mp/OLYN31eYwMS
9ZzC5kAYIBndCcTCkVcJBBNX5RMdtu+2y2ZSK+jD7ILvDFaL0r2QbKeSPAL3atNs
18x6ImThDo1+/DyJ+w8pZEQzQwaq0N95Mavu7YrQx+EC5YEGADQkNCau3IE6HeOs
xSICFf02jU7Gbd+wCrJj2fSjIxru0io4vODyiy5QgCV9+YdL6/lWqe7KLh9Hk/nE
VcllJbv3dI6RvKHEc3DOPRmsSlMFagoNX7w/v/z94D2AVUK/KSW81YxuycPHQmok
h6IeNEh7T4w9ewpOV/m5+my2gFLiNW7wLUsIy8Hn/lyJpHoKAxsoXBcYRJhSDUev
4JXjb+b+WhxRDLN7RVm33zaN05+aMZe7NOFv6fgqF9V38hzaOIIWxcsaLwdwcmuc
t06/zytRZHzYphNvK4Wbp/OCMF1kh49VNY5jku3OsV3eWcXJVynOfqMuqLFa13qU
BvQ6V6mQqpnJ46MRPIs/EMdGdk+HCn+iuVQl3n/UZN5bApqZ9l5crddjPkXI+G/v
4AxKtWtRI9E50k68yfxUcB6zdPD79Aui+Y8vhnPOAkMFAwFz0YSd/NQAx0tAxsWs
bj8jOUfs7esxAkawtETggVjvehT+xyjFAnHCZ6BIkWAxjIZqCCYV4lkTVhlG+W5Y
e0qj0TYJQUXAWFBcWs7f3YNPbU7tjKX/poKf1L64irTBovYVw4t4raoMzHp+fe50
HYNVF92aYkyV2r7WLLU1hl5xdDKnuBYtiX9BU85Ku86WWFQNagO9/yPy2TQPBOF2
XLO75b3TKfQbt/ez1el51qz4lYDHn3UdMsSFC6iedyOgKapGY87nex4Vc/6ib06x
KDlLFbgkMCAjRsPNqM0sMqyv9o0jMFs1nrX6xJ4JzJTBP9HkZfDe89CnhxxBE79m
Rps/Z9q6HcDXivKLDxSVe2JxSk5Vatg8P/NKoIN5KzOUB/PqDhd4uOw/JXUzP9MQ
kwd9q3OtAiSRHEgbm+PISXzbFw6XHylzuDDUi5fLtV3Qk4HN/6DFkyKEyzILIWkA
zjxfEjVaYjAIUHQrTka6gUR6k+hLiqWwEzd5hOGiJMpZ9KvNlOZZgPDiZA4uoZIE
vifHlmixm696/bRLHjcj5QsfnIwm0I7eS5LApKKJsfUC8jul4ec9U8MKTe4YkNyn
GS/J5ZfcIACXWbKjuvdhpZFdeyU2wXuvApztdBAvRqD8UCO1EblmasPF/FrcLdhL
DUho1Fo2rtJRz0qKD8P9+f+LlXvQclUmxy8R6r/R5CR4HbwIWMpIS2ZP9H4ig4j5
/vOHib9Ui253d3EPfY0TxQGW4lnD0eTtuTk/VJrLBtgd6hh828Q4hyHJyZjYBA3q
E7dMHdkdOGn9JiRo8q5lDArMCbsz7oWB0n+gCd2xjMIsgRyC2U4cHZ+ZxcitS53K
gAn0TsggqtOZL0ZLk4J5hz60y4BoW+nSdfDffZ9rhOgRv9cALGiCG6kXjEbHlZE2
6bM9lgQXEjv85KLF+wtjkHNPbgOdLwqFibIuNXWlQkbxdx0IgC4Cl/OPcF2LgRZL
m/NKUU5z4IexCGX98upcVkCdaI/Z997kKBCGPi3OVeUZafIYhQk90WBiSYhueW1v
zFyJvk+adDMnNwfxWjNPpmOobM1hsqdcRhdeiLPTfv+0H7EmI3blop4HDu4D/VGq
ZR8S5b+vsW/I0jkbuDia2Tj77Gu8RYySs4myliD0ApBflkqiEySMXA+jOBoRnrrM
sjT0GJ4NdJqbXnt1RAWQMvKgahKOqZeH/69B/iUkjDZLwjCqX5qm6x53T53/OYMi
/9BK8GrUYqHehGHIZ52Ws/OPMg1RFekz1pPb+XYkCnvTozIZnwoBLiB6xsAR7jQR
1sRzj4YcYgv/CF4764QGYD24egFqxVhmDO56M40VNytHv+2EnZtrv6JM5tSgk09l
SosDKGcOdYMS4ybctvJayTLI37u79MFaHo1U42O48gamHdp6MDS9ds3szniqi/8k
e9BU19r8EP364sKn6nueylPryzT6w/3RcV5sSrvhP81dvXhFXYLpBAfGvPw5s1dG
akWPwKl8b2HClX2U08KawgmIDRSlxP0hBLayPBzppaLMIAROQHYE0PRQWE2XUbZm
mI8D00PMmyj7StvlAOJZUTX5yuDXojaKv4MS0C64W2KOAUdlbdOer5ecG0J8cELI
uMSTxPqWUknvgAWxxOquUlW/RiJfpwyCYj48T08U3acbMltjf/YbjceRIHxPABt5
DyDCMaN4eauUKGulD1xSvpqgURTG8Wa4iGvqIXNXOnTQhy0x6BFkthiiPvdoXXPl
q95MM8FRSymoo2C5NnNendzrYCuRkYM34ODwRe5R44HDytikAJ9Zsbw8lkey7Zku
hOmjb6nfRUJ3/I4fF3vLy+KsOqBGDxF6LcjK0FBfz2On7vhIx7N8MEDd7O9KRVrF
u0zBLggb9TuOB3QMyMWBcPBD4NpkIn007N9VTGTAEaFE3jSbup5TF4WnwvAjS1ig
OuPGdpkaH355cH1f2aQhyMPNLbKxYq3BGg8yHXgkgKumVKhCymGyyKNviHLp4Nm2
EQX22rQ/HKnCb6aT8NWKgNIO8L2M3QuepWOW5kTPs+yFC+DoznVFC0wC1M+WarXM
1CgYKc13zM1n2Cs4D/h0Rrl68kiOdEozthKq/CiKLO4bv9JYVbndGYRHP+Pf1Pe/
R7iBkiDlA/1QFsfspafbtERJRZkUsW2kqPoUc1T7WsZydS+lOjTNzkYkkhnL7aRJ
lflMNYeRhcI1JmSr6SZTmWv8ejuY5x9P9Chv8DAnqYXuUR9hCQBgUb4dJfyteLx6
Oxp2tZNbT0GTR9lSfrDvwTwIcyrLBE5zjpoADtYwuZ49KdymQtVdJEgZ/ZO1QDrs
1r0HH+k3zrXErvLm5/8pWgLoYipuajAMBIHcFhYE+2c/GaUoqWp6LOGKGL3run2W
dsNcJNowCUACsrXuIDg0Q1bGqKgfJXHg0HV6p24WXE+mN0j2GucWs8hcDxyNZQ4W
UU/ZzW6ZIxbB8hv/b0Hz0nhh448rNq6xeykRCEqoqKokO2nAbydPwHk8CWTeYNAi
xvVbhC1UygzwDWxsB+lgn4vFTo7qG1pdPTZ9yUEmum+7BL47eon71OrlwKpMk8Oo
QXIakwThRh4Kg6Jo38PrjzWsZSDJh6y+a69AF7mIXJkr+tAvuKt8QvjOdSyxZ8Ql
DNALvi/v29Mw0oMYlFtT8Fq5lAok3Hvl/0yQpuMFZBc1h6KaIek8UNurV1yUR/PL
Obq/bXxlvBNzExCcJol9iPs8KO3y9EylzQOY4zeqJrOgUmmje9X92QYW8/BIMJwb
QySwWcLiPJbTkyxYCAbRGguJ0mfqzGnDG3YnFbzPiyCwOd2P9730xCUKA+4bqRXc
t1fiD28eGLSa2EndYjOCQhHJa5c5zJb9gKNj2AJore3GnllgeJeFy5eXRab2uaqG
MgZy7Wi5lmT2C0uRQe6FplEUnh5mAFTfWc32BRo6KIfY56qXABTqzu+ktALI1kSQ
p8vEBPGXDnEVWpA2rt4Pgcm9EeLt0PdHdf0ugFMYaPXtv27ODzhhUrIuRjSySpis
1N4TPDn0eLLqcgXJ3rx35osDJuy934wT4ImCL0CLpsJEOLynwOjwQKMU/h/Xq7/Z
FlkBRPYwFWLoAbqro7iLTlyCK9BqLxnt0bx3vddgonV6+HBSOjfLD/MCoAxnZToR
KoKunT52Q/T/MOPHoflIrOVOWLqkAarJxEZQDv+W0CbsgrPZDyVvMDUobT/F39v9
L5ka3Uqp3vuy1YHOh7tMxJJDYbH72ZBMPeKdSOS5YC92cliG2E5upqB7GY2yPT1+
hpwH8Hdx1z9/8GZsYQG1eNyDEAZvHyvBGDdN1YmwrhJiOysSxOPQg8OSnA9I70nB
tyARtfAFATQD5OBcED7h+9F4jaGfC5Lf0J2XIHK2iGcTNJ4X1dEvH7/wVX7zjP98
is/NIzI5vs5PeV50U8SQ6uA+ZUbpug8TFMvqNjAyBcElJFhriMw8eVDkpx6Tyd8Y
g52jagu9Y8l7DuEZZNenWdtPlG+0sBpTVe+bZUXwZfKvTH3D4/0gGV1I0lSy/cNG
tfHzfKlYLlFiJtAToR4csdpt1/MnKvW17uf34PsPtEWr2ov67j2g21Glk09ObxnK
BJFkm5MJ+8Qaf+oWeP7vXkFaz09M1FDD8xz+lWB773adTHAkNQ6JYGx2qLxHtUFk
RYS1Q6ZkiYJyOANs11jBRd4QCWbSB2uT0rzSpLG4PljXQyWVcHvtbcFvQkzD5MeJ
rn1Cum2d39rBI6NUmVlUT2PV0m4xervBkPEBGR5usKe0jWFYQAdthfHctGvjY9z9
aI6oiXelFkBQxvUepui40ua4l4qT/tpuJZrrXpzzU3cS1+XfSCkPJKAnmMVcB6nQ
dQFFgYoc7PZnFK3pnZhdUupgBPzCov7QDwxLLUFiogvMaotm1sIIj45tqQSZHyco
C1dizdp5rHLiGf76HEcB4W5xWFhytaSvG2TC4MRW6GeADUzFDABfWZKkyUjK3Sap
wxEi0etUGdgZNCEVS7a/irl1/7mwxojicMLFHzT+H0x95Iqzo3zjZTDetemBhGNr
DOSsMAxoyjGtLHOl15bP8C6p3SF5+fPRi7dJKSpQynhjRf7UBFYUwbtuuM35CjXs
WOCxxLKAYeTn6SnZ+FuK5HTyxkq63zpgb9NF7thQ6QEU6O37K7GcsJHIwGUaaQjQ
/gVPRZXos7p4dGKXp6eMGcs4sh874d0Hb2yGiX6wYdZtiIKR+m0ebP7dzpYHsB4I
bSFSC/kgDuGP9/Lzj0RA8JzoTEd/ok0fZF/l1uHTZtaF2XkyIu8dk4kLDCo/rAvy
PJsvHue0AhN+qqWWUljqHPXfvcx3CQoZMOvGO3gEz+5nvu+Dxnf9PZRJYKIZSWpg
s0QbQWork2GtgyXhyz+VTSsrKX+FgpGS4dcDnBWhaW7okREhBsNwul9AXwZEcHF2
47+U0ep3aqz9u0YxvShPFuRI2kURVDFt8oR82aZRLKD8/ju6Fqkv3DeXPCJ20fjt
xKE0tS3f/O+OE2uO9Dm8ULEnH7eUI7MvIGMf0gv4m8oqsbqWzmfizmcdQ1+DJqCL
x8q+gVB+XKgeUvY4qIQkWYb5MlgxnJ69i3IuEDoT4NucAoudZEnt3jyjvoh40X4V
GOu8/nMyT1d1JjR8TFKrtejXIYJqiTQc84yqR8CBpfyUPt/w6V+Z+4nkazmheV/U
Qk/IvJOoKktzTnGNERWDxqEs64pLX7J14mfsFyPlWWHndLmUZMj6+dDeHc1+seSB
nmBh+xJBVm6bBHAHB0t2329bE4qTdoCQjkKAOP07Yj4R7LY3mghIT0eNnvH98J/t
mKywZwMmvV4SXmZGWMcOPWor/4Y6OR+U1wvhnK5odgIo86dXj1x5LAxuT3nYt+8A
GmEWdz5/jMe8a3qc1QF3JjlNq2aCzTPEWhufht7YR1Zd+ipI5Bu0Pm6jH99YDUlR
n8BYUEUk5If093OuVgpre4RuDJDwXLs9YE8+0TO3lakuPANEg6SlKEMi03QoCEMw
/l/3ZK4x04fZ8cOZw8smKq+HyzJ0AnCYjQS/gPRhBp5cRguWV0vTu20Bv3eFbCmv
QbPYsfvd/GDASMjXf/KI+OMUzykAbhPxB1psTaMPE3Ny9YhNlI+A7/+dFK/Lwhvw
EhvrY8JSOkKpbylYCRyLZvSIipSeIQFJQpCnbsJnR+dLi1HGoh3Qz3RKRsALEjZM
dOipEQaeoTNlT+cG7VCOCIKo+CQZwP3qmKjc7JhAZarVYQQAvy0mOIJiPsok2rwH
bdsu85qiIeG3/PWC5j4Ho2V00bbX+Vm7zZtuaoI/lk38AonKEgG2rIbgQidRz5My
rGiIqLR/khNIw/sxaIeHVZ1k1sD8mMKrDU4G/qXDZQtue5hQ3xXpSsGM2//fr3Q3
DHr04jDx/mMx5jhVggBvo8s1YXUij2DMQ3jrpB/qquYFVLhDpWLByiTr0uKNEWxD
aayXCgMKNNemBPriOUS5d8P36YpPmZyer9bBGpzdtjnx8wtDdq5sFi1+BN0kyk7Z
/h2GxtUU3ZGYXpeTm+crjswxnkP4tKLLMmhNmx9jOJwuJx5aMDEjHu39vGjpUH8S
/EY9Am8Uw2/BzGEQJOzhFpi1EYDoniSjwg0U61mTIxY47u9XRFJYVzAeIh/e1Dvy
mfqilSvjyCWzUK7+LrQNI+slroW3quS24mVppKYgOghw0XGOVvddrnSAk+pc6ISI
5DMxfCLXbDSNu8zsgQHEoDFMy5d35D28oxrchAVdDOiZMmDfDKbF1tpEdCX1MZvb
MoxbVFUH5m8g8wAI9CPvqXc80MvJtGsjhPMJ/fR2P+j25JC/lRRVvbUJHmWyJiqr
g7B/UfcLH8id8zgqCngIsT9gI1kpnnfSwdGb4SmY8GQiKllodBqKdD3SZG9voMMc
2JEfNiBumfHsw0miHTwg6raU/ZKYB35twTYumlP7v9sIqD/ago57cmr4aByTDV0m
2CHTjaB6zTDoZNWcRO+/qq/zWSoN3dY8q71TtzS0FEeqE+L45RCxwfigPzdu/pwu
bLXhE2MHg2wdl89sQ4iNY4hgYd5umbaU9djyHu7orh6IBT+35LjRqYb/di0nMhas
MaCFiHBSEdc+DgwPjh0jSkNoN8jaH7M3fBXWNQ2NnzUpK48reS0HDyM6q5Cf15v8
F0Ys4dLoOYtX7wdcOQ0ZxnuosUK5xdvdYY2sF12or143/ADAR7Pm/Ka5YE6arXj9
Q9CzUQdBLSAr5q0N2yXS5KjgMGNRp8/ntocu42PWP/isTyJ4Rz6RaNa8kYU6G7KF
4oLhc+AwjSrLZb1C3ZvsWA72eLrl44yIk1z8TFgxE/eL3b3gobcGSo4E7x5EGcuE
iU1uaJ7yNJfTNxTwdJBUq2rWYVlJn28rYTWNpWTYLo55Ijj+uAGwFVoAe1LgwVCA
J1QewZlsjTIdQN9kxDU0LE3nDeYrnlJr8rJyT3rl9Q6vX1FPNHQvIZ65qkgKfFAJ
lC2GwNfR9nUtsKLtwKn6JfF3lsUXgW4YpLWPtic9Ezzz/3Y5EckhEU55kgKNg7m0
jMMidw2vsm43e/8M9hPyibeScfweq7Ebsxc/pRf+f29+SuQZoSbrsynaygy4kxpX
H2clLksUkCV/WJebm9txdOto2vdpNwCkmBBlBahPbMUCKdny1vyyW805uDowebmW
0fDRWFg+V6PcaMgiRbeWxXk+/WILd48Z8z7jBFQ2492lCNFEvyhf1sLBdfDs8J/d
ScTq6j2Y/kl7b6gQ6OODP6wSJP7/3/yurzmBTigur4vZULS6XSt4krydnAvr3fWv
kfKzNl7KT4LroRm+lQ3dVcyoJM9kAO3eZL2bJI+fhnoKcWkWP1aOQ4A6xU+Yo4Ad
f5ZVECYYwBwgeu0wAvHJN0fMl2x9S6a4bdpxa+7IeTlUg/kBXZMVLpn3PGgYJi9+
2DoXScY5zT7fqJV8KbpnA5NJ+y4aMqceV1wZe9ByMais8SSJhEpuK/AIJpYOl48l
ZE/lsaetpZTccrM+cfH1jVLyqmWrcKfCuWy4APPEooLqs6AZk9HappOQ2Ue1EE+n
L2hlADPSXLvx6CBNtL7uwyXGvsRpfR01oHZtjs/Bk6mvaOJzBPqxwLze68Q+eFPP
5xE90Ie1bg0CyHgMU4bVJpGwF18+hpqeNiSvoBlpTHWZIu2+uNuxEgvaPmTtNk1m
PK+ygrAkdZ7pRvNtDNkC8Zl+3R4EZ6OYfffZahzGVItUtOtkLjCqIwYPdp0X/jIM
ila1fZ05gS1SwSWu5YibGJbIiXBTfGX+eGCHx0RrTfNkOl8nX6Re7kAOdBPoNlWr
8Xg0NcoeUuBLz9JWfnR1t6AEV6a89dZ8cN/FuTBP/E1OBx9wT3sU0PmItqWGfYU8
zei+QpVmtR6c1fPEy3t1i41rMK5GG95p63lefKaLQ950Gco6q+OAUyBg4DsQ6/k/
GTegk+WSlNHsa2cBsiAhme+4nxCgQjjje030OLBiytRQ/AHcSihLboWf0A2ktgXW
K4cjwSgznfZlI+ydrAzS/IiU6yo6UrOph3xfpySRdN4iUQvqIJ+LjhneH4vgI9fB
2wJkXPfKglyeHOKaYmvSy9UT4j51S7ImhNI3JN2NaFybS2O0KiUfFyC1f1D+p+qJ
j/NM3GTWd98TBT+gjo/41aopO9HWObHBaMHvdBSXe3ndVhnWnD0Fy62Br77ZBG0T
3mZUZNy2oJwKKGGMN9V97b9ZkIVM1K5nUpVjPCsylTuNzBo7GW/TFQ8J5gJ3QtOy
pujY5WEvtrcTGSs4qRwzsER68ucEfdjYoZFFAnrfE3rZafT/Ha/AsEzGAvTiOYxK
KeU8YZqQiTZQfnEBa+g+AUN8x4z0qZ+5V4pCuOZi1QS9lzKUO1nIkBZQSLAwHRL2
CPfTpDvZ0Wj4UlouSisOde/rAGdFQRLUJM+3z8upYFCIucRm+Ympka5zeSv6tOxR
h9G7dNYNnCb5cb/tF9W25Wlr+9HGHH0tkEAC6XzZi1QR+spS8spb9tH+CwcYCRMk
u8ZLZ3vuSKOx0o8iALN++/dUS8bpnUANqkdwH81sMt4YBCQaa9Y7dKFjca8SUm97
+D3mW8GW4rJtW29uUnix0I5l1pP11YtlZ3Kz+hyiukfykSWWjhol/ZV8bHCFc9wy
LRXXsrp7tXXCOp9jUBH/QnwM+ixp9XbBeXCgKbaUSba0X4J1ofKwiha9OfuG24/T
oQnMdzeeM9UluxpRH9ALGodbX8EOTCzLxNQt38umqI1jdo9Xd82ljhGo+0/9xuf8
10JhWV78UCTh7uaOM0LSLiVvO0xJjU7Wp/VWjXooEvCsnhX+dIx4NN1aPr1b5Gmf
u/FOYVuYy9/lvZ9WyGhRTuwMk9nEA1qiUsyX+Jld4hbRBybccb6rk/VPx4ibxPpc
U7xqaR3wGKIMxFOo+R2UUVy+sPInSEuRypXDQmiH8DjX89vG+4utwFy7fLXAAnAb
qcWeAsxdqABh/ky3eJaPhALKIlN5yN1UkGiuZJ0ScpwFBoquqM5rqeBlBERze9Eo
JaWvy5Qvz5jNUl/O86Pn+3/NhPGM+f9G7QjPpo2BTPYBFJ/n6mFxXgTZqhMKROpj
TVa39Wua5N1AoXNTVJ9SsMz8btIHOJg4Nidn8yXH31ulOyMQJVNTs4w+uyeJYW5J
1LQAj7fC/iiE0EdqXFh50CPfR26HT5/cHX4XQyDx11ndW68LyPW2nHjQJZYw2QwT
mFCbeW5TK/RbTuIATn8KAhYgO5mJVDIOYqTnIscbd/ZfUokYvEBy3Vlqv1TzLID3
IvBbS162icKy07izit2RKTZ8wVH/Jh0Obl15d5HP0vQe/Hlq0AO4VTjgDmfaIOHx
xu0eMJcKSGA59Ko9MwyZ75uIz/UtdK2x5r7j60Xbvelt/NaPevdmd+6qzvX7VgoP
vFLHFuVhJyk4z3BEeXc9vmdar4KvXNMyygq1PyzN4tKpEF0QDk4aIFslUIltHXKb
VAlHnm+JRX9UUfA/6IybtHZMqWdZlETOjqzDcZnARG/M6BBM9aAg+rrWbOejIBnx
CvhCQ/5ACiED2OI512lLXIsARa7KmC046OPbcYfMfrhDck3heIdAUr06S9hhWrwZ
wSywgfCV4GXa9TWSoKVUukdBqgp1IxSVMhBtNkkQ6wXL4zQevwi4izBUvt2bbl2Z
ta4F5pVjLtzxmL7Uog8n9iAO5cksxIUawSLH57uwREuNeI4kTVkvjsDS7jUJGzt5
R9+E3PIdna6rEc3KxwxiJhkX3Pz9GK0pLt4WlKsbUPFVTwM1dOpLd2pUp08mhmVD
HulKkmNSM/udrl7z9m+pOBDTKQPN/kaluTaVziah/lbyemxuzlxDfumuWG8MYQR3
ENuhkAMUkaFmXJ2k5u1sK1YKi+Y21kTg0twWDaUHfOecKuLiw2J8blCA8yIS0ZR+
Jc3d2ndFls2vtaJIixT5WEuFzZm22R4ApNWDDP+XxWY6IKPevJIImx797wzkbcP6
Cq6fuIcBwedycNPLKwLK+dQpQVBspgSajA3UaIEklyh0F6ATAQX5O4DbbLl2VX0n
Y9f4KqVW3vGzoGUyCasThJ30KLDU0bWgMJyP01v5Y+4ISPqo0L9M6ujY0CPx7kDr
sjH/FWAVpUlIDe7lng3noaUpuJYsLPsodxcq8F5LnER4/Dcr/mCHXH6Y+PjcO7EV
5BHFhOWMjTR/sTUxbrzmooZfiws3iNTlyVKSJ1+PmWS8ii1dV3xBSpY8tw3BASpt
je6X0Ii8nERgUXkF8tbOwN3wpb3w1gdvMo8iQiSk8edL+FDaEyc8pxYU42Toh10f
xGWOAyKhc+Xs/qkT5nQMtOznnAXlJrNaB1qtSKWa4SZJV8ezbSHZSyHo/usD7Abg
+82KR+5Ymc4Eq9bGgDEWyI+gqg5wUkfE5eSHDmqD9f1LWF87jQUJq6s8Gj9YJVF8
BCq9np0g8i6j43yd3Ffu/OS3V/57RqrUrNx36bdOF7WEtLuG71mJ4X90T5wv0H1z
gY5n9Bswlt2CxxJiIMHtBVTT4E7Be/pLdtg06JucI5uDMDUFPMUf5ZKWhZlTVUBu
s3MTvVTsUXsOmR+aX+BfhU1Kkdy/t1DpNv0WtPg1D0t0XkmBcjEjv0qCKV8YLzjE
BEqVIzcL4Ir+5pzU+7OVrF0xTSPdkvuW6qcGg8VaK7YTxgy/H+SpXVg29lSd+LZT
k8jxvQ7u1O9eD4b0nFoAI3BexH70sRxE8uePRX9ukn8q2lu5CPPeeALZ8KFBBGm6
4OsSUY7u3VGVjXlbH49OD8+tNcg6TG48kDCKnYZSHIKYKF2RZVGUIN4wlJeZPRu5
lzhDw3eXlw2VnZz1z4991LtniEYdK3C0L1O9u2UNut+ceXhR2urjjOHnBV73fqUo
UwzdMi/3bHkJEzeyWpevIvu1cfpXLAkglfRM4pfRdm+8O6MK9Zhqht/6RHD8kSrJ
33BuM2zeThDdNk2Jjb9I6fjRUiJRXzKZxjVwTD4OQWrGEm5KmzZKVH7HEoD9HjLO
eimspha7g5WRjhEoST5+KYzYRq2R0cDYtwbtNBfQzFzx5g/PkDEzCk4lBvBjahoL
WnX/4NwBcegbwkPPipw2ylW4kVMP3KXtl2Kb3uF1kxqwnredFLQyRUHAJzzaQhcF
PESSUTQatzrgaWLtKOkynaF/dU6WEM89h+qLbNkzuK0s0yFHXZFMrifHsMKp/nyY
GuTdUQitzJ2SyCX3e7s16IJEAMgS0XAmp5COkZzsceXZyeZcnHswMKtiq2SRvU3O
y+9HylG//t3LwzVcUnMIZGjipRekLm6T7jaEghm7BBngY5UK/5HYE9WYSIfApANP
qxdHO8k+Eb74aVsaRyCSMyVMucIa7trhdCBnoN6c4e9iT/mkr8jyap+JEQx1QRkz
ac47/uUmMofV+WKgQTn5JkCrq1objnXLM4tz/gK3T4Wdpq8t903ERgAdROvPlouV
OlAab6gyJh23xoZonlEy6/QWx8aUvhrVQWLJwdxdHNyoFAlKn4mykRsWO5PSqQSh
g1DsnfaKfB7OGqZrHfHcT3nK2GSKflp06lyU1kmBW9+9xrDQlsSfyW4B2iknOhio
LftJvAaAa4wbYvKF9MVuJxJ5jMJZ3nOGS6uWR/hMTLA0wFNe2N+b93ayvdHu+pbP
j03WnGRdGoMFdCK03GXJvrQi0NzZ5CDBKHfUlgUQlSEl2l6Gp7bBS8pICUfzUD2a
KShmDm0vW16qmk/0w3X/8Yo/FSBH10khEFDA1fQrrMiNXJdK+qvaLxCrAtm+YqnR
3XUDqallbsyO4KpqSF5j+c0H99m9jinlXucTkKXyJWPs8A8/gUeEYzteIbo9E9Nc
WtSFKGqYDpCDH/BksmWs0Rw/PG7ce5gnWpW1Ts8yPJ0Io8Sj3MEZZhNmmVbHdLOR
jBs/lcYvWvI5sNwwwtjzG69bNzwt0IQYKEYVIwCaFcPMrR4UVSHMEk+wOuM+o2Gl
ax7NFfLUv8gKO1S5OGQ38CT+CF+hq1bRLb/87ZhjWzegnytdr1GrxI4k1SkmjQXM
w2Wd2wj0OMDnWQWJQmL4ktE+XVehm7yf47055GaB4g/fKRLmbbIOzp7P1AkrLbG2
18euiSZb7hBtcNZ5N149eYUcg4wyEjXysMsQv9dKXe0WRAHtVzDjBrtdPCW4r/oQ
VDZM9338jz5zwavX+5wMqw2jPrH5ydSQZen+Kh8GPisKDhkiQkj9tjjgvrRAjkOG
pwji7UMGHRzNraG42pI57VrvBGDaRbKo3//TxGN97AR2BB4K31V4dNdUGcLzq9aO
bHYxA4lLBWaonInSHt6svSaQ65NwX/f+alv65e3pznZZY0wCz6U3QRY01qYUEhTf
BY9lWr4Mq/lDrgczEP0frbuyXhUVd/BPZgMBC+WI48W3eZK9tf8tWTn3T0NDZpTz
ogMLGY7zB8054L1eEiFJiinj4ulNlLjUD50uy0Axv8G1GOISVBcsbFUCuk8dBJJo
FGyZhod5HsW1wNBtuUJZ1e40uRm8tWZ2no5zH3rEpTRcfklf9OM3nu23xGt3TGD6
sDg3794ejg0cahO6f2xxIZYFo0Ez/IM+OIetn8COVRSRjmZPDhYDe4lCwuQGTAw9
AG58mEmGVu6zgf3/0Oq5YOEB8Zd2kyl7CDFc3/aGskM5JPajiZi6HxN5fsNkSKij
sDA2RybRZtzkMj2Cd0jTGlIIM7b6/gEPjKkiWQlNEPcbyJkuF+k5Zbgju713iTjE
ZHzaKpe8ddPj3rG8JHfFPn7XkMRbWr6uQWz1tBWsHtKLruXj70yJuyt+5ANJDbcx
pZe0EAAtRCWZqtkvGJz6IKxjgl/7LgqMwgj9qz20gPjSdEPCM4AOZiN3wmdwjvLF
jIhjQfpJYyS6Nujw3Ro8OYUkhAnynraOl8fzfd6asD24xFzivaXXBH2vIUM21lNH
1DRKm7vWIqLGO1l7qDoPBrJGNib+goQHcCx5/IBsVthpctR/rpbtV6Ubj9tYNqJn
1kB7ur0xULjeQHxZ2kHsaubpTIelKeAs1ttQht4Y/koNaK2W8GrheJ+MuqekA5rO
YuuDw3H8mJuwLwWUacs4kcQZyhpO3hYGYM7vwzvcMXnlsWkMULRwXxRkPP/CIirU
s23TVaSc1MqqOl0m4Xoo/ZbpVhErKiuadkyhGfaEtHWXkGZt1Ilme8ISn6/hm3yR
RlciD0S4XR01+HQEi7/TpUSxq6XHULTshaGVzsYiqUHKNP35kdCur/lVMQrv3Hp0
M71dO0cPJlW+OGIGwCnr5dFc/jli+M/7Lhc7Pupr53udDS92nYb7jPkcOMbfjrBQ
pu9oGswIjjtHs9WXknOU4f5riZ5u9ruvc2jHaYblZpvTXxHDZi5fxhczM+IZyrZk
PHIHYKlUeQCD4oeG8yzOko75jvtUMXquti9w1Q940iEwgsYPPQEUr6EhI3frgZs8
8HVLqUlm91usk+yq7W6mItoNukp0u7g0F1sw9uGA6gHEradYnLd/8IEoYCqKasbS
IkpCYBtkL15of/7SDwzapJlVGpHXb34/2M5t7r8MR2rc0Ye+fRyEOzWNrwv97w3h
ildBaypVAgfnHWixizFrv9REzuzp4ptzQtfXSZ2mbTp/7HBNNNgoUu5Eia/r5izn
divZroa+DAHQlZzDwmO4ItmKsQ6yrjrSQgtTDBB14U8PHeyxW3FMOZdiz3AfWsIB
Kaf4uqj0BIamm1tIDs5xHZKewsqY7Stkp886nnkJkkxEEIHkTRzlKK9K/rDGcAPm
5jyxQJKqPlfgyUQJw5n0qmGUgmeQP3GH9PVxKd3e4g+ABjtep/EvLqG8AVjxMDHM
t7+eX/1aOGWP/YJSqjeagc8MoC4ND+diFFl9/0B/PZw=
`pragma protect end_protected
