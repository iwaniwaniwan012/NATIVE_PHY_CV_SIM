`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
o1CXsL3gyAcCuZSRn7RbSwQBuvmB1kR6tMSS/oL998Whg4WPvLg8aoei6Xu5K9Br
RAcaWXl5QBDpLA8/ORJXKyIsKM4j8U7wuTXbLLFF8759WIuZAMQwvGc4ptp+A2C1
x8CmQA3BsHy1q/2M5wCDHsISKehsJ0LCO7fePEeWY4k=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2976)
5DQmUBKG4lP+1jh+Q/TKp3lQOOqLstMUzET5lMMgr+o5E0uZLLjewPa3bBbC3SDv
RC4lPkM62E38d8dq/rVWsZ9L+H/N8994u60VY+J38XocJFx0HdZ6DlOAHd7c8H8d
evXBGyhiqegoHEeLodjr3ln36q4tbxBakurkvT5IRZUZUyfkspg5prV5Wn4G0ZPf
wLe6MuNsV0esD0mK16qb0vTIwA/ygxWkun8UjIfM37fslswV8+YEADCw54Ox7Abn
Zb6PxzB7OD5R80p7h1E7Fm353MwThBciZTY1r8hMn8LbpYqdVhlr4T6gg93ByGgO
YWCsMJJASBSVM4UGERqpWJrTbiLrIaCpm4bENeSkgb0rrJh8/ydUQOtX7XE05Z+X
nktgp09yHDqe4DksonNVZgQ+77kt6Sp6+hofpTZ8pdIyOvGkZFPok+T5UrZG4nqL
Fw5jdxxNwnPpu0B13UnC9tUN7ZYTBeeJEKBiDQssLJck803OMqmbrVSwzjJ7Lk8K
yt28au/4c25AdO0eSp25aObqRAX/9gX9EGPj00vdA1FGd0EGmxWFlVfOutSf6t7m
aoic3w1ZOaSVi2yaY8nFTsIAyUXo4wBHL6HcigvbfXWUWZSwoBoE8UorGoZAVCPz
v7FKd9gj44yBzL6wJT56St6idKN7fYkS1OdKdozens7xkOM7wWq2qt+ZUepKYXEH
3uOgGSqAIlylUyzRdAQY/mowNsVmvknJ5AEFaF/mtYJi2SuoTRvHZkkrWTfNTPuh
x1Fl//9NknPMkW4qpnPen5OMDbEkK+TVzcrmpx1Ic7cmYafkbZHVuwc34sRRTGd4
wbvDn6eQqofuQyUhA/p8/P1AE/R8Jw7l2S5Tx0/QXWfCYH2ZtnM5OSUD9LRLf2sH
0I+/stbRiYViZcPtsb18gWQGYm4/y0XJSL+0kXpoAdXGmkpE6OCX0RZ/HyA5C+tX
F/t21iIKyv5q9P64g2PnmxRHWo9NvjNv8Nx/1jeDv1BACiAVUFA2RvGeOe7olK1D
g1clXA+Xj7NkqmgxG/5/7OD/gGO3amcOGBrvA2DDuR3Ho5zPhW71EJryL0wMx+FS
WtFO9dCyeqDF1ZvKgZWzoRh8Wns9oQgLuDct1RXvJpaT5+ZAOAC9T3cH59yAQWf6
YcvatczcsgojN8LJB5+iMWIvgsfvcYTuWuZlC+1sXIJ/J6TDNdLFRTLiVp3uNYoS
hrkkHnMrbhI4Wy1fIU9vCCtEEqB6fotYR5Zw9wzzSdq7yachLUUC/yVLVZgvNheu
ZBfjqu0kPujAFR9eFWEoPGyfzLlfOrhSk9OoIszAHnAldpjxXavTPurwn4GJydnO
GJdQ31j9/UpVNc3tKdNFsvPXS+7KVq96eJ3/ex5Szp4z4/0Zf1La5cwNdxIY7o2P
Ig0umCBub6673fCz5tVwliAEv7egYup4T9MjHBuOIvThpl4ookbG0CtYBnPbV+9k
TtRuwr+RjvD356rVB6QY/xVvH61QM0PTpICW8XwykrpbzdwtGZyDkBwb2SNPk2Ka
PJkGWcMcOPSg/m9g4LmcpcD0MPc7ObqUqc1mEoffu2nxV/Eg64sntlZLqGGsFHA/
wIKMgnjs/0GAmlxMCTLGssbRVHoAtSkv0hprQlp0KOJZ4V/ToU8NpwlUprwQvA4X
SkiTr3rMoQz5D7lNxORRDR9m3T4CFIljYXsnxcw2bnxW2AhsQL2sZhMQrS4tAuQz
m9VW2LmSGzUrkpCoI1LTyvOYYggmkWwU5+7dmV+FVJUZJ2TieNMWI73PVdaphmVE
GGEU5KIz2Eck2br/xr1Uzs5cuiB9HzddNum8Ncym3HCnvFO93jTT8YZUUpemHFZn
HZANMakY7GRr29q3N6h/V/9hScc2iIaZOPaKScNgBmy51kfD8W2vSaGxLJ/zu88I
sSRaDj6ENs4hosIt56v/9heMwOAbcHFnz56RSCIf0O+t+z1kv/dHH25NkLF1Imss
J8ujluPVjqQFDnBjXQ+TkwZY6vQskGPs+1gEkmwyRobWFYeZA672uTB99U+M5Fi/
fQDdIscCXXDCDpLcXoy5FoYaKjyPonO6GfSpQD7I4e7rgpkSSGNThVYzuQ3tbqHb
1A4GwDNUEE8A5Yus+gfujOvxzA8ANaVLVOkTmyfOXoYY1NFN3BjjuYLNoE3ugKpD
WnYIxMBp82i5EU7i7mDnEXoss7OwOe+Qh8mkXC1LpYlCvZLBYNqbj+vAhChCBj5O
rworlK/goMR15wPvLziZRqrk9Cxpc7TsB//rDjBbchiSQ/hwecPJ/QruFWrjH9px
Yjhn2cFQuRQPaAgE6xmdt1b4HXSJfGASMRlEJReb+UKxKlNMK/65mnV4whmwKBfk
dz4l9UZYgUeAyHrx+G8eB93UtRNa8HGC7e16L/5niYvFkFmkF9nhHfvCHr7ZdeRB
UHifT+hQgE/iSVmFanC+4YshhGgjiDjPjVecwxyv3WS6uKa3YBtEiAsK+QUL6ZOy
tpkxCSa6B7Q4rOFCUrBbvSdSFjKIcC08vaXzjfzWUiRYIhwnwn9ftxurlIxmzpdP
4qX15jhFgI0U6pRXPNrz24R9En08Rv5jx28Z9/4kQNfMs4i0Jff4XUwaUJRrJnwa
FA+29kAfjjgUkhJc0W8NRz56GYKGR1XofJ6KcoDLGdng+EoaMt4U+xwOdnWViHXM
OKf/AjMNc54prVLAoqqanVrUc1iMCdUjlBHmV5XtwO3ujceErSBkuhoTVxDhlLK2
Mol+zh/ElounRZqS1HQcVeZxP0Z63Z9yJVIfgORX77JZc8vDiCA36VFH4EZzMwry
Obhu8kjXfUYmcbOWyH91xG4Vjz1NhLTSW/Se+xmDdD8xnlQaVLx3Tem6R6pfMGhl
XT4Mn8L7n97G2gX9P8AB80A9yZCuUHdjuvtyEh4lGC0Qy5aqVJa0eSwSteD8ActF
dr/TPiPtwucFKIOFEhNxLjvXYcbYsqxu/pravUgXUyhCVz+rZ3vS7zAIbZaX8ea6
ExHv/hkqeb+mZTDHFlCcO18Dzf/0xGKa628uz+u8qLWWXfgf8FUvDzOLakxWfWz1
KJijqUYUff4JqKpW1nsLZ73QlXI+6AipKTikiYXnQcL+hdg1DDf2SegogJqKCIvl
EWomJWIHxkOQZtnmBBP+CacTcuuTnykFpRvweqRTKdXVVTg2bQZM9fBWuQxm2Hg9
Kap7yNAEs6Vok1hwHI15f19LGVJHRevY18qt3KrVHfgUV5ph7oCU7gMzH7EcVpMa
ChF+c+1Sjns/jRslU5H2NmvZdCA0EtSudOQcM+1EYVQtguU9zVxqHq6G2pHrR7Qn
YsM07NmABlXxyk0+yVFcj2rCSfWA503pwi4Hz6o9UPkNkjYXt8SXYW2oXc7oRkc1
nnIdhoY32j/PiXfjBEra9TdVxsoOqtUbixWkHM6pvgfrUaywwaHShYXEuF5ILOjJ
zaDVtJTLfPGfUDet5OnN7hu5WHBMZn74LOlVLSgQybMFVSAZbssRBtRCxmNZR/He
JeX5nAZRJkN/Vs6kXNvunTbKIqnNbj7NeGEqMvhf3HJV3mXgwG7kGHS2IlQcv2cH
1dVv8KtgzjF60aDcDP2J7/DR0bqZML+5jOJBvMwpjpnjm+nUsIZQ1p95uNTwjsHF
LGnq/2fmFKEwA2kmlCUmIphoEFftMX56XTRiWnfNAyuThV06EGYY3VyrSmHdaaL0
7dDMfiOUEc+4CmyTcEjH5WeQmhp1ggtZoQAdT1VSIvhPxo084Rh1y2yZ+Er+vofV
If8usmIYNlq22w3A7fpCxgKYvS0vBohNNGV/2pnMHAdVL9IkyEhT3U09Q0C1rAyt
u1oysB7i3dSF8q0NVdxWALpz0ZdkHMjL7XtMdkABKPDVxSCFHuQVsBRFA7Rl6ZOa
QtU2pI/B4/aY3dTVYnduYsTET5ISP0fgKCH+rgnZ3XnbAFPCOYuKoinJ2vQ0aM0Z
`pragma protect end_protected
