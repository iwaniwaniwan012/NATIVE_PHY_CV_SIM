`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MPQ34z1h4qRCUnUA9LhBEIE0SC0cFZp22HU6TVxtIbc1LK3pO7i6XWFoOm6AI23A
HGnZKFsCnrm2hDlRiVanZiLKOOA8HOFIwJhPWEyPieYjnD2AaPDp29bupDM/Wvor
CJGIz8kN8vt9bdgfo6rLnMjTE39Q9fr3OIm58N+ysrU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3200)
Ju3FSXYhiDeBveiQpu0dOuWSbNArNw02adoQi+lePLIVVDN9v//Hj/cuj4fBq5ZS
pHUD520C1W2QVbwQ/YpzJqWcS/mSpndTZpd19XHIQ7z82SNRpLQOLkZfu6mJSfPY
/EDGsfpjWtBZwX7epZXirAC8c/Ahn7/sHtveNvdT9mBREowLEi+2Tap1kY/za/HR
0pDYPnMxHitW3eMcREy1UW8RuGuttuuLMheKclyfVgYRaN6viuRzbyTKyUy+mMgl
sngUTeer82TDHz4MXPXU4Th/3ejp4yNfefFu6FDAhpT1hoHxbeIbLqSV6h1veq67
4pOv0xhgBvHcS5LV7NpTJ3l3MR7O5MfLJTwP2ZxhDQIZSOsrEY5J5a1NEWZfrRKO
4K6GU0UOKl/KT22JY/ZpR8m3gmljtErIWSJi9eDagThurT1Jf+C5P1p8z2KaGgYA
k3OazTH8gdIMeO9PR+wn7WJeKUcFdGRw5bJUVJZ8xJv15DGtZW8iDwd0pC6HB2OV
zUQ0bwBWtqdhsep4z29evapNo0qULvxRlRBX+R3LHh31gHJEjeZUtiUj/1zA2qmD
8FT4R7kQ8TzN/q33jlTlDZopCuF3hcTE48LnJynALv5aGgzrQTnkmPx/PG/mQwUL
HGkWzlolUkiRUq5S8IIMlYs0dlJ2UwjeH1j9ytghMOMBM3Edpb4yNUj1Zkh5i/IP
b44FNr0aNtrUzSHftASvnaAbup/hcUXu6tH8gGPMMvoVArfZGhsvfR03XnwO6Y3X
WgH2JRPoujsVzfQ+auz8Wc6qnKsYfaReTqoToJCZBmPewMmeEiZBp3pKnu9Expcb
MPFO56j7G5bGEvD/azY+UYFbOqJj6ZhkMC8N4SjTmtikLn1Q32WTVgefrQahPfAX
hJ2tvCFNqRcdXh8sVBKcnofj+/ZR7nzRl6Ex8lf7wTU4xeI+m9JW2rfxZ0ulpVbo
cONY/2YsDEbbkuwG9C5HzPntKx7qzISttagMExVxIYVdk54Ud7gga2MQPcAIrYgV
R2aMOjcc0eMYMYr3rRlvtayJL9D6NzEVKaWMVrv0iBr+qfEuIcCFPS022ydgdQ11
706f1nj6iy+GQPh92vByMhrnsdZk0PUVvrCDNrdQgMxaYi+pBy/GJSvepP3d2xp+
3b/svkbVdQ0AxoOoYBDPbhCf7KCGKYS1Y730wVtbG+9AUrYLqKujqfdDPa+Vq0e4
SWNQYuwdAutB7zoEopZjcmd6fi/UKl3Kym32xe2Z03WNA4rUQgDkc13XCi6RZk1y
IS4sJ0BzD7Vzh3fKht0+HVhm1Uj1ppsq0ySPv5ZYdFfKtqQ0zNGi75kPQHzZlaJd
caWQ7q4JQZ+fqBpvmTTZHt56JyQs495toS7jtyb4VxyvASXNjGQ4D3jReD0SwDVD
XJLtKgwGEZKx7JSWkZ+H3jaHdtU8Ih+EyNj17sZ+XfRM5hVF1Mcj+O6ckV5xKVVF
iWa7LACApt45Hbg6PEaGE4awrsTev6zF5JfEZZ2rUVOudxLf1rGs+BvwAb24M+Ge
5yFktDxhgMEJPREiV6VhWteUowUdZS1UbAMnr6BRGYj7EmOIjSZpSzGib9Syvf33
rBJ4nqHaxqWemLfDbMiTUFpHV8+OtZRmriMjQgyxOxsLhVpWnu3dWM+uHsLqMJGY
+MqL8losNYmw5fsTcHvJL/cXaNrKZZE3F63ogkD6ncyYEpad9xGiga7tgaY+1I2m
g+zlf2/tARK79O8mYxFA/SWzltSLwFr+jZa5Qi+YEM2SN4u4RyUhcRWVfLRcfq6i
ycPCksdmFKbwn/VoCYq3ppYTQRlyV275Pf6TEJ9N299Ds5Zqx7U1RQWC1jGDLSoT
DScBVhFuNN0aBk5iUmihMu1WDzeYQcC8iIixBY38evd8pZ/MBzBQBQmLMTjE6oXc
p+H5wr8UJNvYc7g26SbOV4IYgvcrZD/4cY4eax4urMOXWgtW29n0wGcBq8/+55+I
9/KoJMQwp9/XNzduLL9TcsrWJA7B7UgtvfnnQShVAQ9uBjZ2VlagCHtmK9npMDIe
6SJmpaJHtLOa6OFKBMWgHobUHHtjF9xriSzGwuUAQlWhkw7jcvPhiWLRb+qhFASU
nN3S8dH8a6hevdoDwXkiHKhhZW++iewQR8B+Wza6PXSQs/ZP5xMqwCQLz/hrWdE0
Pwroc7OvIpjF9iFtPlsmWflVHldpX/OMNnNgzwS0DeSDLWj+jgzrbw3Iy3lNelnV
5pSWIBrmvmUeGxAqK/cdPTl60ORlIk2QSECKdYBUxfgSk0a+mSnwNhapbrt/xMWR
QTBFGX3uIDuZN2+uBDFEMS/Xrc8WGt/dr6ToVvMMPOeMAJ1Cpwx9k50qtKuDjWpx
uINEblnjRQY8JS//C/jBngi/NdB5GyD+6usOkYgLCWUuszM664HNvh5eHgg7LRmY
ZrSMV0O/IWqAVqwXSn7bIanu7o35eLSkgz8u5I6hYVKv4jeRjiwIiJaaB+skCHN6
arfAfdi28U8gh1m4FsYB6qJdWIBjo7+06nvW9ugKQzRkDHBtOXxggIrcTRw6BvZW
xAcyQB8xG9sf+k3BQks8e5Vb9OCPscPJeOK5/rCzJI3kOgchZhXGw6aBmi/51Ja/
QySjUc9X9EnVyw1WOEJRW0YE1xYf1bQ+ineqMMqJZ7YosPn0WRb7jwaHrot8/Cve
SS+zMaey+ql7669RyOXffEJbd2UIrUXILYC9OcQrxK/ukC58Z4CRFGIiSfeI1djE
BzWBTaPodQE5ur+2IW2QibT86hn3qQDE8yvKL5WSJ7zeh6RG/94SRlxB48Z0/l4Y
G1izPz0FSkziSvNY2R55ddX/lCMLZNkd4oRV43UF3wiLGvKwGJfl0PQrMGFrz0qe
3k3Esll8Lk+W6BACMyabQgMkc8gYrEYiAShGNYQgAaYuSpA3SsPhSKjXZ4136gRc
0RtREjiCxZzXkXO7ABQqIPIcSOxZOxtCWVuHzFi77Zf9RzWXKJFWamA+9vPc3q6B
Sm/w+W2VY+m3Y7YOshE5skViD2/p4t2tPXlGPMogpdN/52/iktv8eymZVliQzqLD
JD15An51JZABKFGEu59GfBTBXG9sNfeemS9J0yJd/W1cmCKWkFmhdOmU2377g86k
6/++SoWxTpAal+DWSHlRnV9tkGpMf3uNY8SFwstTIXvkSrNDtB+7lJSwbxU/NLqQ
DgjXIc5WLrT4RFn9o7Dqm22ogGb6IcRXTHr5apwogSu9eHMwMW4dhKwy0kaA0/ml
AiABgnysKj3MWLVqjJPwKDMpAxH7jD+BcE1iXOdxVbG8hqJH7BB0PCPXzckqJolZ
EWRQawqlLwj1W5Ojak+B6/qmyQqP6cIdkGj40uO2V0ojrjbgznihDoXScp1rAhla
jjr6w5Zti9xfXBbBjEvaiZ0bZ8ljwb53SaIKm8lqbUnPyojLA5TuvIYl6R+Or3V8
rPRt+QeVD2FWH9nKM0z+Esq0rR06TSgHFtuCHb3nSW//I8bcnNH4RUPGvkLK7TVu
tiF1G65eC7vB0wu2nIhcnIi/xmJjInoPLgwacvcVU4q8CjXgjDMXyBIR04hBgtwS
Uz7GdJXSsgDwZnGna+xEPgXsQcw5eB79ziwWwOOiciYCGQPo0IHU2WUeDvWOQCpf
IRa6hJcvDy6cTsvzz8KXtKfIUelNLgrzE5qegyPC3TOIghkDDRzsGtIfE+nynDul
wXOa5R6lhbfLc0bQcHaxbNaeznxeN55E8cY0Rh68S4c2koWdmoKcwEaeDEH+v0Yh
oMPqxIYRRghIQx0Vugv245p5ImaZYgWYmBJfdZ7dcIS+8Likml3aB8cEljVsEu7l
N2zuBEb0DsY/mSd+XZ7+o2bWDzwKwiXwF/yZYhQK2FG+L2AAi0jGIumx/lJHSy2N
k0YK2mUepOAQkRM/BhyBG0vieB6qWxK94EgpjBRPI+Vq4cE/clHd3eILj/bPoqrR
Z+1EYR6f3xFlXt/7OK1TDLktC+V17Shv+++JW+qHhTf2XNnRK3BJ3hMnwIpHvLst
Pzb2Yi2UEkRorM+IF6Qw0enuhWiLfEH1wM9FajSDq+R5go+RbJSJVJSiZu8Yo4rR
lNhU1ZnbVeP/loYS9i1COUEPMZFYKOOVah6566TpP0QnSu/QegtE3aOfEAOaprEC
HFrUPWnYfLudejJy8aJH8pQEoAuXPm9ctzQ8pDoGqKdhF18dS7mIS5dLR8kBj82g
dk735bHJYBVFQFGShAlPg6dt28xnBXX0pCWi5ff80xc=
`pragma protect end_protected
