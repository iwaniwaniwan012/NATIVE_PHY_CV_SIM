`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
to/NcnX7+iTvYrBaAAs2CDil2RrSBPZYkY/pCVHAPiNv/EqyzV/rO1uVZQHQvur4
9TS00PlpEpmI3BQv2xVT3iBWctE+4/MC2/rNNXenVBSPtbTCFNRZWev2d14J3fvs
UJrWn1d6ioU6tlkxuk0KdawuqIm00ADEDXG4ANEwGhw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2976)
YpSHMzfiE7tqT4UM/R+VBqb02sFbH5LmnnhIwfMXf19amTLpTCA7ddp+DdLwQq1s
Mc8147ZD75TSss6Sb16CJjJ9k2ShvxFw/vof+iBBCSL49VXF07LXiYgMhDXt4c//
Bm49uyw7tPwycZgdB26vVUpKy8UrjXpMnSdd2Kd0IOs7KGucmPxJnXyVitv2o+Vp
fl5GxPV05NbP5+vQ3Ct6dXOshHoH6WDmbqBr9ayEBHLadC1k+s0lp0njaLKn/eIu
DS28nQIbgk8c45K8KC8WYEdOYrUV7EO68t7StcQMJZNoUzWo2EQqyqw5ht0/HVd5
o5L9wTwsCt16cFAjj4Wxhiim0emDEJuIbgIwJZEwkH+/xSaKaDT5cJB/ZGD9t+Jg
GLkxdCA3meTBSAx49HQKT8hHb76dcV7BDuYNTyZ/0wc9BbonZ1ARBRuMjli//hkp
KWbX1dl8ZNK/cNt8Ks5cDc9vK0VvHWYd5NqGz3HHzU5aqh/pNAWgVYTkZKiJku0F
SQZrGxwQDAlJMn3DiOpQJ9yQ74kKPPf4NAwOciaQUsxT2R/arw76afRgp8ca3Gis
AD1jJxmYNfPWqKl21szDC0m0bhF/bBF/e7OnodSX87e1dJI8Yn1rGeDiJGTAd6nw
QXWP4tfPfSf8vuwYsE8TAVFpd0kZRDRVDfIa84r/EiPtSQtsa+3o6odVRwwTN3ME
arqVR1S21udFJd2b+wrLtj/vuU1BO6xyBN9td12AoVc+zvDJGYhS00fpfsjMY7Q5
w2NS5iTGr6XpedNTp0UfYEAWHlF6+scYRJaZIN/bwFl4rq1ae3TYTvI5XTiH5dlf
yYiPnSLPp+kTehswexftpjKQCfKBvMY9VEcenRbzROQvKMe+yKfe1lMzuH//9wRl
tUt4OVFnAPmbdgEP28A7Y9Uxj3FXj+Ihf6YyqQymxmX6MXKiLZbQnIj/dgwyzwDm
u9Cwf5MIo/2/IFd4x93IkHVIofsfreK2wHe0N9Pj53WZ4QDDg8D4cidWKu2SRdjT
OsHw7IzE9PTxzAfGpC3jYZhyczZjq8p62mXOTrZuJlVLbkMP+hshEm5bvo+Bx4ap
U9Rz+xbtf+z5vxXF+S4JlMLyEuda6bWoGrMxfdAiEC4MfOHjubyazLFM1RUVlePb
LQTS8nK2HHrel3BOQlVAfbGqiA3PxhkDSwX5CdtUxkALpa1hxO8Q7OWT3SPcVGU7
+680eUeRLxkUQKxZpNjtKzc7TLLY23tlMTzQ9n0/mL2gkxB8OVu0UFqWdPssKrew
HMXNDHinkD40/foS9zxeZxY+/2rMp5PprDjOBk/eYXY86K5pjgTrJ89NQMx2OnMN
L67+8Oqfy9BVh1sb/1XkfGq13fgKO+IG+RqzY1H2xUG0gihkkFvq5OX4oq0gbX3o
LV50ow6z6KEkQP1IzpjrMMsApydMh00IPdAvuy3FMa8QMaM/2B8iEBNlfnPLmFyG
tfjMZKokWz3tK79JsLrDuEu3mRqidFGYBjMIMlL69eArEC9oROaasZk33QRG/lzD
eWB4miU6GTQhvCfMDFUXfzCPFyr9WiYpp/jvS4Q91n249nq5xoCKe3HQoScB3krd
UvvS2MQ62lCC4INlJGK52s15cts18o1WgREZB48aQ42y6Ex4hnr+B+UA7M/okd4g
gOpMWMXOnvK9mibsuXpVBWlhQ0OuVEnuIROWNstotCKa83B29F3klkqDDHwn9Tow
c9V3FqW+JmAoUDYwRHf0R3C18rOPlSDgY6dQWZrCdvY/04lFMhdRsahJaIP/zVJv
jd5mpMrDbupBh4OTA9Bc2i7SVPzamc9RHwDH4ai7DAui06KbwM2J5lrqMIQxQwWF
vIgR7NCbI8yidmjVe29TzvfHxOrX7i2ysfWi3cLmNfY6HVqQ3tGMwIonSqZfMeKk
6+7H6IdFeZf/yYy9gfCrkLWcPvmsBNgHilx5Ty8UU7pbQFB/rT9uBczGyvBOMVV1
ZAfyWWq57HPxqIiV5eGzPeN7UWXR6LzytkHtNNx27+DItpFRaMcInh167m5bCqvx
nPGKXNzTX8dcUZbzstSAvSyZmtKMFV1k+F/2JISIWXF/BsUCuQLQ6mDoBb17NQ2l
Ofu700zfxI4LAdUzx87GXQRY2Ze58J71BXykRm3c3fh++D2uYrLm0EDW0GWV3ro+
TqnxkB3KDLa0BJXPj0U5gDtkUXs4C9z9rsYh1nND76lSgNp4iZoJrKHiwPaB0E/1
7d6Dva5kh65FGrqzfDvIa1CjjhB7o3Tntu+4IANpgP1FTiOZCEIXXHfuoWLPjM+V
GDcyqttsXTa4aGOLwXYtuumCnOwr77DwRkp+ViVXQUCj05b0IoBgj5/j19P4wD7M
zicur9pgwadWWUK867uesYAAijdQapVHAtowzA56VeMoGDQgn2674qgwYPEe9Dxr
iJCtoGEj5C7BgqbDRi4w4pS36GIbK6O4WYoxxipp2LjPldT1XJO04J0d/yyjO0CC
5e6Fkyvu3UMAJ1rJK4V/XaRe4FERCNhJ+GWrO7s6GnudpwkbddogP3g3hxLlf0Vq
SoOY5MPh4fH1+TeUoUNmkXdjxsdjeAZWgCMHdPgWs4/rTO2FlVvcaqWD4OGZbK6L
lKOi8oOSc8RWUdiExkfK1hSHkIJhlLTkrt6ZF8OzPnZBi1zSuNz6NAmiIAYpdmoJ
ugXakQUYGC4zdpOWgni37WIa6gayLX14DK8pFP8McTUvtXvY3hfGNLfAEWsW3wQf
ajLv0uh/pEFrWjgiFehKYn7yIXX8f9hBpWxFlSEaoAoagjiVLVAe6CGRt2UY0p97
DDOKaAt0JMeUwaK6IylFyR1OMOXfz7dBaeAGPzUllJtr05n5gEJ2dbzgk0pU/1ow
5Wai81JTDgc3BejRFHYVk4mdZ/w0BaH4dJgW5M/Gq+oYL+FFigouossBHskXKxsU
S7NhO6gTIdLcb+E2saY8cLebG+mztx89XxF9rdeEirYBeTCBuMBPWcupQM4dzANS
NEuxQA+fwPB4bKVYxdQ48mC/83Ww3eVeMKQsqA3OyE9Z+dCilk+H5wmg7nno146u
rR656wH1vGy7OQMFkInrzvzsdHy+H5NfMgoAG89iiE5ZV6YgC52/cqoMJK2AhkRu
Rd4jK/4eM09FGD2WMftdmXyYeGHooC+rAIlU+vJYoxK62QqgudKfPojiRUg0Wrz6
q9SO2BWJD6o4dxNXFRTGWR0gjG4OKShaPJ7OSZSIQvLc9oNRNX0AOQisvw8kydRB
bVp6HBDGDXnFrc8Jf9PW9XzFXxn5/t1TWGFH45uahUFCkQdAkNhVLKLqra77vXU4
53MA4EWtmS29n7YfnXL+26JZLedIsGIv8LcKelynyxXFUf251YnwmK+lfR6C2RlL
UVK5+Nx/8HZbcn/w+uwQPtqbiMKZMvhS362IbjY1Xc2v7d/e5rwUfejd/EaJ6YcB
ySt/ZLixg4r0VG9dwGwwmhuVCO4NwHqZH92M+LS59Zu6pWU7/jGvoVmrWuOIr2zD
bwG+bh1RZmfEKHrBHWoW0jmrnr/JbnnGDHBHrsL7opmevOYtMq67VjL92SbuJs/l
Yhp6rtpFQH2ml4HUc0YoJXOZme1mT1cRQme2onlqR25p4YLaovVTO8dgm5XlJneg
vgmjTqMVu5tHxGe2chF3MfDNj7Ie/FnTFUWk7Nj87Yucp/YyIQr999YD/avg1Om6
vd3ZWx61m8A88nKD1arh1L4E7oGvFuJdJIHrC3HpB/2GtWHuq7zQtE/VDvzLCI5L
98ccaPdBxNgM+uRBlR9HnzIrfalMMeG72Af8G+bzr8CcAO4a12fbYvB0la1obDmS
w06jPsSYXXPqj+Cd0OocRkHGRnoMihb017Ws1y16jxGZXOFVHGvkhg9ht72s4LXq
dhC8wub8B1nhYNB+12l6PBNh43J2ZeWtQgSzkysrtXhlAepbNSdXlb0Vck+oRZQd
`pragma protect end_protected
