`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NmRROAF7imhi7G0B0NXBT4Q1qpm5PfIUhiBvKzdvMzQZ8f85NcqSN8khUFHsOOpw
n+lxFYD8ZHCpFwXXEXyS1JKw7v2DPiL9iqZ8Y1e8hBJVLWOT3W4VCtDih+wOD8MX
H8QE30Xpm501GwyFinWqik3Lpr1bI/erwkZry0omytw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3696)
B913qpawAsleIUij5tRrFN5Oc9i7L91/vOLGgu7nVUYA2XtxhWruOfpjzI52v+a0
qXMvtEDn1Pspqu1liTR6V8SUmR7YS//jufDqY3VDxHoVSXtXVtWEhHsYBi1Tn8pV
sKz+bQbeE5mRF+VXj/+vUOAdj9VUvhQ26eewj/SFzYgVYW3N4+3rht/DAy0//uac
8DC4mMlIdmH5tDcb4k1Ju2dDR0Ipux6+eTAYXyoVXlp6A2TLbqNmSKPy8aaJC4Sr
vo14KPCqVUNCqWJVMhIYvU6xouCBDUFAC4plGI/EvsTjU0r7HamvLVowBnYqngq2
T8lSzCZcR4dE5Lsb4T6Bcet/Oa4B0xlrv0zZSuWf41+N3UYvwA9EkDGCVyWROksP
gUOrBdBwUPq1+eXAjE2Zj7JCErlBvQweECaVrSRZydq3YysuPvFI+XpwiB4K1kxz
2C5M09HtHQKRKuKpQUWAYs6MdfxWURAe6beYNk+guP+QvRZDkSNkbspo7x+IAdLi
4QiLkENwgaOkYWMm17Q6PWE6rrKqlsp1D1nU1fdRkXseih8y0SX8FBEfRx5MOTnC
3sXuwF7hIPuEbVYj9w7IxlRxKWE59BakbS1IIZi5KtnA3w6dzW6z6ozhronxj6Ff
zd6f5PtyZ8QOa8+1Agxwzxsx9w7jivZCQq8XnPMDsUFW//3ORZ5/HkpM6cl0PTLD
Ky1aY42CNfoxwLtqSedxWC8ln3RfMYg7mD0N8fJTVtslPMDG0uwuVDQ2gGuM0IJ0
zfy9uHgl0y4IlNjsEKwjFAzdYLlSVWT97ZAM0K7Z2xVR9uB0zh0l0MSXTM/7+Wvm
vqHdDUq4dkAXu0665DrtQ6uT2L/Vuo1jVrMzPyljRJbYFeGlDNYgpArXnZB8Tnbr
l1WufBxXEj8qqqCRfInnGKopdnmYG+UOm8EOnRfKKTcn4nds0n9RfBBeatF3UO1S
LYUU+GPNVn1dKywei3nrt4dLwJoT706jQrA730uhiEdxaGnLKRsNq7spXloOr3k9
vErtcPmtQUq1thXFimjcoFEb1n47PY6Gxra8rUVMEwXpjjEi2fxT8tM4sCdQXCkV
Oo6lXlR5RktSLtXGYCLGy9RAu5gQJcF1xUcndJpNgkp7zsr1mGWZwp8FMha1t/Il
0DK5MQP/zl1LPMhA/mmnZK/l7N2hrsaHBNMf2xy7mXQL0vNEZhhoka9E/mQtXk4p
tjiW1sT49XRWZ9R7C+XcQEIKSCN8cqUyo30VJ9kxG/IgYqDyxBKNnRBSMj1n7mKv
B9/L6OpnxsMciB56CjDnMmXqgjyFs7Tii+aHlmo1LmrK06YFs3b2jUdQQe7JJRPd
bqfS8HykwnWnEXzou7a9WIhY5thGQJAczdZ9WlUXpmNAXynnaAq2mhH+nr7aHraX
PV1S77LD/dTHi0YYheuFd3nz1LZhKHsTLYP1FzlwK5szWaVDE+bTLcKKpHvvfhDJ
aFHl62j3tfZs5WTYGN0+OMvCY6pgmNkZL3OFzPUubnPxp9ghpbfhzEqxsnAKr+s8
xcWQXNKxJvx4NVWJ82AqvY4hIaxf7eYkAymbfvUV8gq6a657Icqh3SXwmdmEpxHk
9m+Nehuf2q4one9y8iJeNjQSmNAAAGuZNkUPEPskN8W3mLHdzD1ksM6RNdAmUeHs
oqoq7iuTXvzzzk6m7JANrfmgXajdoVz0t5ZwnrhLLDzxWEQsb/ozHniYYROkmcU7
rH9u0dZo9YHXbfbVkcFugOC4ggbR4xrPo7HNqpwhcCF76KSbXexG3WC2dsOdpqm+
EvVLVGAdVtg3OvOEwysq7UuuB+eglp7DDDF0pbGnqsKUXr3mlZHWthc+5cNG50ct
9gnr/AUpTIrqTfyL5DFxFljtISHIINeQ8gxwFgxQ4HDH1VFsQ3maFbnrqmRKNeUR
y1FMerg+BYglxhrLBq9gJNzFS98jdHSk7CrJTNZT8+uSMlwgqFykvpIIPvo3j6Uz
g5Snl/XoDnTr6peqYHPy4g4UUGWFn92L5K8UcO0BqOu6Wn4nxS4dwDK/5FcMd+nE
mAXUwUTzDw9YaIF7QYdljVC68eOEgCGtHZ+4ls9M7xyrMJq58tFWrbdNRVdQ+uC6
/WKge+Zzg7u/OY8LvDi9xRhFnUbXHdgWJ9JKdTxCydaIoSX9Dj4pFhz2rIMZkMSo
oncM4WOa/h4zQhIE+YQouq9YQGJ1ywLP2QggGzreDjgP4d3pIymume+l960/g+Xk
MDOKxwYd49o2h4D6l0moNYCIZ7OhalnedgivRzrnbx3GuXGu4sVWx+QQF168Rkko
RH91wVIHmny6eQN3HdBq1c7lyvFeRu4c0SHNmOtmLaVxYB4UeUOOhIhLqKtKvSW2
4rhY4sv8AitsFkVtifQUIy3DaufHIIe92h5EdE/wBHmacdRklSSydtiRhQBO5APp
5dGCEuXhZFuveR5dKqkYBQ7sJ8AaoohY4pg9NGJEtgjWUDzdefERuWIq4ZbC9ukC
D8P5/uwXWCBys9bWRv4dlFiRu48+KivPfsaIdOxLKK7Q7AwW94iTiqk0psWwZ9W+
qK2CddOLgXTls761EMt9wXbOET1r/6Pl9I9NLtNXRNZga+Zn1iC9vMKHdIxNiCq1
/1ryMmcw1dpAvkylQxyjSrp30rohJlDZsexWPFsFpYRrncHsO1CVt7bEM9eU2ZvE
Vj0bxDsdsr1KGwj+2Yz6wGSUmkDQmOXELX5F4L9YLW029RP9gq4o72/CQ8+eh+Lu
x7CnPZHHN7iE0FFs6kqMrDfbdkbKKbsOZgxTAi5wrJ2xUh7EV6OUi5rIxwtDbj0y
IyTQpeak6cUcjE//+spNYoMI7G6glY6nbd2X2BlDZSfmuakUOplEJjaUfYeldskD
hpnISJWoNgy1By7R8Ov01B8qUxK58gL5pWd2EbiwXnLO5mbC/E/oqMkwAzhocdVm
UJKXj1HgFn5dHz3ap2v9XgHMI4Go3GSREkjE+IuLOlcUAHeh7L/UGnGi1OOl0LNR
znd/IqHgHA6nlniWgckh6maAVniZWKUhnfUd112X/D0o/EuZWfWRV4KIGsH8QYCJ
kJ2BQYbIwGDivixSjA4o0MqLkM9IPLko/fQeIX9aGmWPPPNFHyDxw0Q53d2OANhF
X8Q7/buYRcPQT3jZaLp5v9yjFIiOF8mOGTonVmWd3m2Wrgc6Ch1nnAyH3RLjjb2F
MDbQHPxEpGTmImrCxhTGZSAk7l5q9cqX7EzMyhjTkjGgO9cC0Gb5y6akn+eu5PQW
GhK14P87vHRlNeXxrXVp5TgQX8/mlTM3CT1epHl4D6trvK+icuUzCnkQ9C5OUXwz
kS/VxnZRIcu+XOl/srL0ZGdE/05TCpC+b8EBjDfeXUqWcSAXhMrdsvcy0oXehPuv
0a6N1fqCRsIACIOWQjepVqGXdD8oMw0NYJynfyoAcgrFMZ6bES85gjEutZKIbU24
+WMTlXUFaeGAFZeYNQH9LPP1s1o9dbYqoaEE4JPEiljmdMwro3wq0N30DFUgh6cy
7NacHaX0khFe6Tfpob/lAuDrh+czlGd0uchwNSJDUbpZnGkueZd/uKRe+wDIrpZ/
fsvJRCFGofjSZhPIrB8rw5uvcHX9RDGuZggc/hTzRzf7QmlZHQ0RaP7Ps7sMVlCh
vrlX4Jb3s0ri2DwZmG3bxOU/LQE7D1OwTnhvnlF0uLMNSaZoeaZxaCkRLM8bVdK/
8Fs5hmrF1RtZPLoF2Yc0P+Kv185wGegHggC8uHxYSFg9kP2CVQqQu3rIqTH8yaEJ
Rg6uGakFs32Xw37hkxC2w3cS8hri802Si1KkmQ/1cX9eNuk1Bercmap0r6AesLtf
m1KSskKHns1XNvue53IdJfz6f9fYpF4LtQCYFqa2m64hX2WTt6+gQ9SPe0GsSbU2
CDMU2IsRDA3cY7XLcUX8I1H4nhq3G2M9H8i5PUzJBatZishL6dMJg4I4RqMkbL8D
0YRSuCADXDJpr0LrUIKwT2pE/F3EEZIDRPgOwI9QKO/PxmskxwzIBNKHTVAmU3E7
nRKSS7vcF4qTctn/myEx4qr+yAbk3eInHaOEnx0bGuRGwSVzL/cwgsmobLdihE3K
I3jTj6DCw7y01w7oN57UT2j1V3uNJo06pYyykBnk9XBBgVXkAvFJlxrNxNlb31LS
LMGyMoF9L/MX/b+1CG6gGxUaM/qLxAA/haUMA5xX2nWhXnDsPNMPYihzyZbJ7vO2
CSUVqHUXql0RZz/YY0Dc80VQReYykmVZdDj7LOe1FRi/egX/dyUuR3rfUfcnrPQ+
T8hTccL2xrPyLIwaHaBV8TzUrQ1dSIoyUG6daYyZjqIuYskudGf0EO7nrF9bOvZd
LdyXetMawd1ckrpvk6nGqqqRPmZVY4X4Nc3w3rl83wSdRUWC8o4iF8IRldS9MQlY
BDv4yD7/Etsr4r6vC18Blc43GNqLnnaeh+1lmj7nQ03QvacqB63JR87tk4mHQLaZ
xsvz7veaKw7Vd1rfVx8TXv7wzYbj7sHGFPTJHL6ePGKRw9rDYMBCxlYDf4tA8KwW
d3y34QuaMm6WLrhi6amt0D7eLqxI34X52CSU4jsD4C6OdyJCE64bEVQl4zrm9DlZ
9TlQT6N5nMF9Iyr1MLwtyOCZbNhUbpML5Q3OYQpZo9iBQmVETQSq7IBxFOibo5i3
QZ2vZmyzwQ2oR4JlJ/Sy7k4ITQzXIea/J9BkZ1e8dubYm421UdX7ti589QMGozZv
1w9IzPBLriPLkq4XiwiDJNZ0PEu8BE44hQRiMzdE0QIzZkWMrtkys+1cK/FWsQuH
4brG+7OVyijCTqxPQUZvJF+7+UzKZpk397H34tsTowuKhDWBNXEC5VTwzq/ZEAgc
iL7qoM9fwksH3mK/lXULYOkgPC/OJk1NW0W4tacXm33RkpTR3eUqHSnlh/Gevp70
`pragma protect end_protected
