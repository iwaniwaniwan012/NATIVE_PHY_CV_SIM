`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mHgEJNEsE0Xtu8PKhgB9SyePpK6NwGdU1i6Gmni0p8RQ4nJc+GMftGWWKrPLyTHw
J0W6hc9EMcON/6pl4tMqZzn/m5sCF4L0iMkHuWv8Z9jzU8VBOEZ0dh6ffX0ZTrX7
ta0+uWROOJSprgJ1nEobX2Q549Mnay6lVC5cM+qoeSk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 103456)
MUjYdRYBHvXch8fIQEiHHYHIP6CJHh+zTd4SBdiFtM5buIFmKY0vLDgjONFiuOZW
jXL1x6CrYIv1RNVpBqbKrGcRxcD+Ib27/yzHx7dfjvgsLsc6ZfPCDR2qTvy9V7ds
K7ADWNQUXB2sLbIxCagfHPVbcLXhBeT7VQ+ORrcm0sQlmuuv3AWyJT/woy0nI9KJ
efU9zv9tCMO8Stk78JzJIDzlD/5cmSCXCK/rB5iGBtlZj5nhgtGA3DGk+Wx/2p0g
E+oZ5+Sl0Pbqbv6IjSqWnQQHMTIy0w4PDvg5+dcOdpi0AnHuMqhRuW8cleao397m
0GZ9J4iVE3Pngk4IU+WLkWHbc6cjrTt08yODrgTeXVwlKZgbZXiOL98/pz3Z1kVe
Jys5wNBmL3GDErUlN2YkGusLCp+J2R+WSzrlSoN/u8ZUQDc8OL+k3qCQhTZVJ0ra
v9ITVxa2RJGhDsUuIxtOKbuMk3StX6zbacSRGWCFKVGKRmQb4hUTNwBd7tAKyXA0
ZMgZfTTTJwjrjDHlqYbPBLR15be+sChilEztCKBsw+64Xx5lUs1qBf8aD+tqnq6h
Ajo46fLClHKbLfh8NdhRz9HuUDk4E6r88j9bLkQUqiHyI4p2W4yYzeSxCDARfxnJ
0Yq0strIsugkDRSK6PHBeVa3CtcBej9nNvrClHD3PcJRwte10/Qw0bMZvlxdYVCv
hkMyK/2okyY2lXj3y1siZOCeEXuuzfFzI1ZbTDXEpRj1aAikWofhVNypXeN0Q5tB
uQqj0rBIogzkowStB0GgrTweKiL5REU+PrUB2CJdWduCGczp2TkiHNIWL4v3BX6l
jAqJLFPP7YAv/B26IgGVpyIK90kBLj/obxN1bQQj0pMZkRK6ryMLPRtyUdD09tOq
Dily9ViuucLjSXZjTo5HbCbBQmfrws92qluQ+Hzz3Sf1HnOMHDEnPZb08SFLTf70
KnCTeT8jxiS8blJy71yoQe/5579oGMcBFAtWqp7s7KdzXUoqjPZB4wY8g6G61iUs
IuN2QxLqCCjaOLqMYYHQB2WJLeqoTI9wYcVMxjbLYuyBxajppmr1MbJacNSXD/TT
htMcc+QgS+pXt0OozMDOGConKZtfnXu1FzYcTdRtSMwj/1WW9RFigMFZyD+hRRxc
MqKw5DSS28GUNP76V+4v1SKwkF2eSLoXuPBoImPC5OAV4Mnk0blIsSrRsYaR9T1w
rUs9AsjoN3T0w6TiFTU7/Y4ep/KTAb4OUE0kIn+YMB8T1uzm/AYpk+TJTtZTrYd7
OCM3zLnth2HnNkaVxzqvDLPVqYO6r+qZ1OX61tJi3BSFzHdqH/E/jFnqj8bjyEhe
/NaxteltR4gSM/On9Gjq9lu2B0KhtIabJUus2IRLfV1bJpymP/Gw91ZKj/r3QGlK
nkwghvNxT5D19+1M1LgBUWf0wlHH2JnERYjT7CfXFoWirhS2cqnvlOHNsqfszHjr
jcX5lDM4FVqUhiEf66iaV24v+CfJ1FCI0AaxJUAppl65c9Aq1mgOPTQP8DnxWq1Z
iNJRQilMnCakHk3Hmex+xpeNBABfgLc0Ts23EMHIXQtr2WIMVbGZx9jweb50F4cS
EE17/GBthZzw9k5jANL1HPvNQKd6hcUrY76/UB8G5qU0Edb33BJvLT4tLpwFaDtR
4VvArIsBYQKoSKLUcawdAs3sKZqxTnb/0ASnTxOxv8MnGp03CxrO7UW1b6YhOarN
Up94eIpuVhnHOVITYxGi1OgEG9t6SX9m9x1u4OilVOOYirFAntcpJPRKMoexoIU3
46b+xCnF8cmHybxw/y/CXIgYGMmxJP3Xjl8GnYmlvjy/1ar/5gfSli+6ZQsTE/4A
z3WYtKkckOhB17r8UwiD4Jf1CbLXURgT6hStToIzDwSwfGWrbQ+ibwGveZMp0sa6
mPh1NFldBbzRIx2u2L9xL5Dh37CYegiUq5eins9q14mseDn8PJTNQ70L4pbonk2e
1eUFr99XSKP72EMEmc55MD4vxNOyC7CGi2Wg2HDdQEts3S/BGeQvDHVaPuBQ/HSz
mf79Mj/cE27Zf3l8Yl07AQ/ZSI/dZQ5GkbrkcRaI3oCXsthyQQmDrKUDV7pWDcZm
MJMIyEY0+qxYkbSEbRHDr4w9lPzKVHPSSyEhUbVG3nYcuPQIxPa9P21ng/GcTFBI
GFgdYxhFIbDeBk0urwK/IjTFiCxVQCl2V5S65/qxg5tnjysCOT1nhK6LVnqQJ+o3
++kfxTmJWomFfcwCuaM9cL6/ukuhBeufRzz/pe+fjNbC/X9Kzptwhzo/cjKD07ny
hCnmlvSVd8StE2ixabXZ1v7C3BSD1iUZWuZUe9Fi2FzGgI3YO0EmzjEayGAI61JO
aAhH2kthUgE/acQL0yEJWjvZvL7B0lMLrB/MggOuJc2PZuikHIgOtio2dXHxLjqG
qRFoC8K2WVIiKfU8/y3N2DpqldF/04YpgNixxLOQIFAkep0NnIJkV6aiSa6WNYnq
opBBHhawIEoB73kmEXZT4O6Irzf/9RE4pO11LYV8ROhxo6sW7puaXxN6SGrgUCyq
8Wf5KVT6wJI6DMxuFhcc3gBZ4hS6i5dlfnw5seIltEH1mQe6Y3bWgOTKPn6R9sqP
5Di/J0L/B51L07XnQLayNdd4jxqExwlbBYimYld42v42IaoJ1lwI+GtqrY0rcGLh
98xNyeCUYUU1SqXoJ2MaFIT/GDq5ZZ1HAiRMeXYqfHyKRgZKw05CZ7Hg+aBYi4KD
c9390dFOCUXnBSmzVmO3Y3uc1mbJH+DP8nITIX9k0MGNi2JfezsAiF6JiGGnE3Pq
dF4xs1sETBkx6Mbyv+T7TKA1pEkyWRaCVI37+ma+aMGmW5RDJ4Y4rsjw9lFusQ1m
nJBug4aSUR8fzDQm/pNDIIDk00bP3sI0Z0nFerhGr6mp6X/A34/3xPRCvgOTMq4z
lv9wfeySMBvBHGhzmgtwNKCyzMcLEcmxoGp2HFC1kSk1A6C7511jAsFe1/DBqKit
O+WmWARTBqxGdxHlnsw0ChhdGHhdhaLbIZb4SZ72rwygafoHyTGEYNeK+oTW3m/0
4Lpxo4AtUpO8fbfWzQquDjQYWlrw7Vbl5BYkn/mCp5ieW4eicn8rSni5sNNXmm2W
Hcq4Y9XeO5gj+JG6f8XxJgjRKMxZFguAtV4i1PPv8cGCoeF0mvjJ4E6B/fdOK5Om
xqXIDLUXpEsmvdnyO7ghWXsdQ+ZyiR8mnPThFOjty6FSs6LZzT3BfZ4S6fJoRCq6
JZdB78jEzZUro9K5LIK2tO1kzmTxC9P/yfSAY5LFsMLvLuXs9xPGmyT17vphTlWm
1nOOSvP0fxsnypqJFrO0DCKtRSLRmXWd2kx9I76Jbh7pShftP1aMOSwGG6ls1RVH
5y7zYANYApBvR2IrP8VDmEfJ5UkEB9lOHysyR8TB0XQ0sKIf3aCOh3Iuzk43v6so
vBuy+m3z0vFAiVsIyjoBUwUrkEmjgCSunMm1kfaL+EZOoUVFoBYVpa3E6Tr1wiA8
8DwQVc/UMTQpEpwB/Ff/vAvLrHH+WGkYpDsUFb2o7gHlEBqB1848LkUW69t/IqmM
RJj3YTHLyvcOmAXfLC4Jwe2OvRVbawi6Dg3udtxKosF6ge6fN9faleASRbBuwZfl
aYUvNL75UBHUxeFoNu1kHU86OiAN8jStkpdM3Mvw305ZTY8e5PiFZAGQzzNFK9u3
GLNb01dY/m0kiVX1jZBfYlCuLbrTxzhvtfvZHQGiqUjvKLozZ5GlniMC6J2SjErO
FFZO2qQR4vh5/gflVJ751JHBR/6IQ0qh/PNM30OOK3HmyHXVaWQkMtKjoVTbPpZu
Df26kfcDo+scKgE4IBeL+Wi5OZpcJg+gYuwDSCAET+JGz6ddYnEzrV1Vh2MyQ6Du
m7CN++K5W2FSxyHe347JfHahHUhCGex/526cRcsf9cISlaZt0maOyq6lGH0W34pH
uDQ6Sl/jWHiqs49eWKJ0eCbj1V/QHe2HoKwmWF+LMN9OeFj1+BkWOXZuhJopI0bf
YlwA9EOt6lHBGfumYafeudAa/FpKOkpzQj9oO9J93f1Yaz+IUfJ+9cZSLOnsoR8H
pGqrmuVMchrn0lMb+elcRgsAFUdLSvtUw0vQYqDV6tyXpwSmtgCMpvQRF4wWed6U
vhbhdOczGLOOEfFApYlupnoy3phpY476b/cVmE0IwnTjPFevZdZ246nWBggxbztB
x0GxCUlvODWfr+c/OLw5CtN1j98zJRlDHzitnsqD3ct/4LN//mKeqIXHUGVxRQx3
RElCUxDPDRmfz1dGryJBSuU+NJM1bokajvfYd2SHghd69NvFnRQQmeUEDkod5wnH
0ebvvXLhi2WjnylSpdv4nVkT/aGLoB8M19VazH6mESB9Y1Ru77/gsZWFwaoY6ulF
HMcBsus6QklZhpyR84CEC0Oy9BLezSGFZ1PsFFn/FdUfYTDO9nTbQ8X0+VV48puG
c7lLIhVJdEbqrcQyAljPz+S1AKLNMBydhiEoqf+meVYudWb4eY9je8kCWDM9emTp
jB3uXPvB4Ot3E7pnwvQ7DkgVjNws7L9n1WYPqE33HO3Wz8MGXgpPCr1Ly7anqPre
uTgMH3YxCQuTcICs5v48J2HoTpjniOGjmIgqkXPgfD6rDIldYpVdua3zQHPo7meJ
1jnh4fy7o52e+k9NCK3cmTXBbsHIZrW2p2+VvZ11r/awk3K5QEjpq1XsVxlEyy0J
TTRqRvD4E0U3CQ7gq3NADKmEtTNRBAR2SnVFWCYK1cK/SyxaJ/qpBzrR6R8JL+nE
fraSQ6513Q6szu20lb2PNpXm4xK4vZL6ekA4vEqc7P0wq3fMWWVuwzlITLCXWLGT
t95d6Z1N4VHr2vyP5hTUdwj6Kb9OxO4Uwyi13IrBiR4ml8HWwNFY7AHaMqzXSmsL
hQfF8Pnv/GQ7dLtke7vHo0sARjUowqGwSwzVKUJ8TqcMpP889avp+FBwCyIHTfui
3XZW3FTKJ9WX4OZ16H0MNdGV+AsQ+qKUNL5hAKJA9tKJtaImdsK56sP7rhWSaEC+
BM/FH03ZOYj3lLNfaXtMNuMDxmB94Ru2KYC9coPqQPqRHdxvNqGuVVmjo8mvlq1x
bdlXVucjVZz57EI/G3MPBnR5M6jDs2mEAwX1ydinITZ1tfQPOMsJjUaGWCcQsnpD
XUMOt7z/SqyzcUlwdRSe28JyOIomv+f/0PVoa0kM1AqV3eBmP049w3YYSdkW2a7r
RznJonVWqXZ5SkSqwaAL8HCPI+nClBtQ4Hf/SEqlCvPboFeZkeclbICXjHET//NJ
3mmb3hODRuPdXHBJEKd+I4RUKiPW0aOQSIoz9rZ5JyOCc1k2cSpQHawHPwyBhbK7
EKfU124cZfJjfbNt2rc78w6prWHsp0oKPEB61vs0P/bzlGPWcvHLxKqVfsvafw1i
LIxzyYiPPMLO+7wVQjp9x2/pcox8v5swa+Z7JNpzdRtKf9gE8uBkBewo5k6rTxpr
lSOsuwxreu/ra5bKIAqi/VkX89mUSywgfPvbdaO2BjFBQl72q7hQFdMqvNdR4qTK
yu3ZHWAtKbtG39WKcPz2rwtCHAHGdTXMImcCVsWAiiVEWEEt2tEC80ewrKXVWNxi
4nmzwNtYA6eHqcSmUshXHm1YpxgHaQekYEXF4/UNV4jA3hdwflmlgS+1FqMYSptx
ZoSqK8PUEBKg4UeHQTzJ+4Iv56UYacyTeeq6AUAIUAAj28+82UNHuuvLSvZVlp8+
j5PN65y+Sg9tTW6l9B+kaBai3i1VRJsKOX5eka/qCW3DQNb9NB2kI8fr5Uu8u+j4
98TtvmVI9mkPAN8RsEh6M1S7cXLAU6/G/2pdyvlSiNKsvfpdZ58l0KwRlM3CYTuP
BKp30jVoUG9wYvQSPS3LXkkwG6oz8Gh9K06f/3dAUkeldrUTmf07fOePpMExJ51y
gRXd1LK+qRImY7AycxJJQWwpU1uNZEQfocaZXNO/0DVY44TY/AKN2OUKrDCdHmrr
6hipadW6w7Mva8lMk0Gi1Pl9L30PZANnmRlHqsVh0KtCI92/cwZtB2K9gZXOa3Da
X3BUl7hmzLoDLxtDy0ZkX+TI5gmVAzIefVJ0YWq5X9aelOPHlNz7+uyOcZM44a6N
SKekbDnBTIMSjOpvjRbI6pNAjkqK8GWFys07Ojz4udWtpK82iNIEqCEtorBB0OeM
kXgegoVvVOjC+fznkID50oqTKeQkHZOK85N7djIsbb8Nsvu29GRyQn0+f51/r5xY
9MBmXCPWj2mjAIECRBj2ZPUdvEY0/mFW83Gy+6T4P3Ak8y+9xYbB7Pp/rWjRKv5v
NmXt+qaYeT8NaPRkzjNT6gYOCFGns5coxZ3CpQQ0YmKkin7GujrJFAYjWAjn3h2J
eoQHFDO25UyyY0wlFtNc5RwwY0IClWYnqav2xTV8Nq9el9S26nSfOkIGlerzsCxK
upCaqvX8MoFUfiX2jPx3SqH6l8Tk7OuA2nWgPgSOPYdazTlqGUyerKouksnIPjUq
QkrARHz7K9YT/HKNfW4Wjhu/jGw+c4IuT3QFskWX4vfZy/7xxFcNl262VcaYjfxa
ZPr6BtEdjriVd+hldWFQN7s3NO7g0Vg9rzn3lAyQv+y0irMYmpJVyLf7XCdjceh/
3CShIwT0OsAwbuPid18F24yhWinrl0NNYgqnrUN+H7CbsYYGD8ltPbGh029N2zoc
R2lIgw6NuVCQjDhG/aoR8WuZ6Dp2DUjeV4EQxSumz/CYQZh41a7aodGY8QsESRpH
doFtwvZU8NJ/kryUFMeGHg914vjNDLLpxQK6/rKHUc7eaaIe/8MZImyVCFT0rHJ8
6TCqrbTblp6AhjkYG4+lJpOFqle4e5EnbJJbZaMSnUkfPQ0j+MtG2gPrtt19J3EI
WwCwmu6plGUvz7dsW+cDfCv+mauo5lmIirlrXQ+n3LN9D8cmlpXAKHoDIcrxwIB8
WRRo9u7mNYaBiMJScT+Kai+OEbH3leh2E+GMg13OUT5NTl2K+TP42VUBR2LFqHVK
GUs7WFM/oXrylBUPXWRs/xRth3OEOLRIegjoLZnQgmyKVnp7MBkc7dJ6eUk9MMP/
bOUNHu/bEIETI8Fau30syj9pcqyEfIY0GwewtaPBsJ+yQXpbs0j+SrzmskVmhfVT
YYNWP+A/w0vIqu+ZDZwRhBwLceE2BF9XoaZGZ021V0shf82gmwwuTNYBHicmJPIS
22zLDgQnidFUR4+wVsS8md8yhlwvHGQf3WZ7Q5TWk3BHS8e1odqFf9a+DyvbW3Zk
ex3XhKAucSKPP32yoAZk8W0IZ8NxA9YiGcLEhvVRWdjw93azXAs7GApKVn0svWDz
K8RYlPnw0ckYTJVOJ8g4frlOMH1hLXoUx0/O1DHSixxV4CgpTFddiSNTcWucZSE6
bYYkhSLBy+ceKktNRxEKKfBD3LYeL6ycK2K/Dz0DVxyRs4YM6RJR1wwMqJ+OR1sH
Q2ubVlFrTO6NnlnxeAXMVjGyz9/PQApvL/lyfeWfobZgtFywiipqZdEZPozsP2W2
gdCf1TX3I6Z/sHXuqubKdIr7NybyPoYI9lEgS4Wk9TZLpb+rlkTlkBBKMQlppvjm
v2iIFVvDC6QoSsVW/5zV7WWsC9pzZTuhO4Je+VkSCzaMwZmiRHS7cCe/P6jukAXh
YeU1uEfmh2kzhg/JgblaUydaqDcu64AO88VDA3ooLbP9LEJa+WPj4no7+eSpJ6k3
5dasZYZhQiQ2b6W5NAzLL5XfIBR1yEUeDG4P60i7j9g4Vx4RFne2QkM2aACR+SYu
6Ozy55SPrtRTAj0F0FolvLlYnugdVnotoydSQy6pnGgyKWS5bkLMH7DzmNNV1Ev+
vHlhNI9x3X3blatsskMyf6VsNQbNtmNZDSYu9tqvUjqkMac5BEvZwUHLtNlqtDj4
ErQbNEGx6BottbBMyot+j6MxbFzOizwZgNfRh/kaHoGIADSfrPU6+LVxBHFRjR77
H4/BHtlHKMffCKe8dZIa/enXeAvbMB8/w8YZZptdYHd2dsl1zHvbAUpt/DaesIeQ
Hg7lFbh5Hv1Jx7hETmT0Nh7VRqE87QP3E8437JjXdr7bLVcxUZfVs835nnR3gjHk
HaHy6yrIc59SGwnqXaSCzZAg1kEcewwkGuEGiHkMdl2EI34fDdiXqdfdUfMYQHmb
qzQ2ALGuGz5RQjV1m4osjGTGuk/w9tfKflsjlxe5rXcPwZKBpKrFxB5+G2w5zDao
uPb49wbL34xFEL0SoWA9OhBgNh0DvUUw4fIxFWxiUBC5I/2tCQbOA27o3aLqXW7a
zRqnEbN+389rwyiEfjwGKD+0qxg0xCOgoHGaGv4/LKzyUe72vJrjvhbnnnfEOg+P
Qsd6rR81D0jc3W8JQzYA7t1QfRtADuu82QpwTKtGH3n0ikkB5cpsYauux6WOtMKI
A1102RE3uFtatHGiUGbBdyqOCwpcLk+nZAvPdaH02yx43SPGthORwgYjC6fBhULc
M5jnKci4wXi7vE897Gn/187ribNiXkDW2WyiB92a5qt+VMsgvn51Rh1d8Omx35RG
P6/s9bfl8G+OBHeV6dGbfJ3bY9KoEWjS88OIckYmeAQHeyWd5U/NZ77FTk4f/B+x
9/4fpjTN2wcD7CnGthd2MHhQoX72uOH2fZdM5tVj3BeyF/+QPKWAuzSemwTZehUI
8VVLn/SYrCFfzYZsGnb+E/5uYzpTlboIn0Wkkf4WtES5266TYTRs6PHLWucSIhTA
Eo+RMlIah302+PzxQ2d56FZmfBnj8i0Jw0kyeyh2qltna/RRVZbiGzLNaN1tWDAq
+gykcRQTwQ/QxJo3hBt54HH7Imk1LMJvjJGb7rMqTEOwyylalkLNi9WhSsluZXHr
V6q5OxkCtRyUPHU5cS/U9ufnwqPKEmHGhw2tSML3pp0i/eMsttu6SuXfwapQA0dU
MMz96MUmeC/gkt47Ojka5qDDieHQlcbaDVSitcnDNlEFApZ0e15pmR/Yp3M3xOkz
woP5TLpjqXCytQuWM1IzxwTeXWHG0T2DcMPrXzIotjiO6/lOdxBmvkh89XPvYyrm
X4Nx3TKwFsDJp/Z/6UvxqbYO9VZfXGMbUifRiEzCottBsiWgQnPHzeJi/xMI47la
vG+nIvKYKspSsdzkIIXf4txNaQa6gpnt+T8r210aDYTHmnvEuMbGHnR7y2lgiNiE
cwckR0XxswfII2rlzbgDLpz8jTbRgqYtiOM3r7iiyCTcuLMXC9Aa7Oa8l0bEqX1x
OMfI8FYzlLULYYFYXlJ3F857EPfiy0Os4Kf5c8FJuoYex7CkUlz0hZMzrmNpbiD3
Mxaudg8TnCG332V5iCRL8CtMPwEU+URdeSXNWiAwzX1GfeLicRxyV8J2VPWtjIqH
bienXX1/Elqe27rNAvqqaQb4D6M/ttRl9KzVx4IJSsqKtxS9rjdMw0CCjKzRKfyA
Q4IigTRLdk4LcFGsBv+0RCnwRBvm1z8fSbh9GmSZ9P87fQ/eVcVokug7ZfLJI38X
gLQ/cASVlarugS/hQTxi1GUGukRiemroJRTsEzsE6t6CjHcSOpsoVsO8wPJOhMQ+
Uma2fVGCsU+kRNJK2Ut1EgEoYks9YCQ+hyEAFZLazMw3kmWRzs5F4TFsQC4iLbcf
3ogcVHajRwdWJPNU72IpW7BBqUp1UNleuO1hVZyNkRuX9KMMk2gBPlcqLzCnxehp
TzrDu2sAQvRRtfsJvwNyZiXZbilkGK783VZCvXmmWDrhKCM9QtSEQRy1WmCZuz8r
yKGbQwqKf5zn+oPBxPBDvSn3HGu6j5ReiYjcU4RgcjcQ+1Tv/BA3rPEi9CCyfnAS
/vjdfAOWLwbCyAjcyGsHQyOq1OvoxgYldvDa0vZtnz8FjROd/xW6IKvOBXR2qOYi
D+DKsqBkSmXOnLZ6HFYzz2wgthX+1ekZS1U8DeGMWRVndCX33XDW+bEuoNf8hUhY
JyWx9L6J2uCl5cGzR6uMA/ixArcbupxKSl5YRKjvHkxkm+Nq2mh6eIr5Ewcs3fow
TQ2v1I6LAUk+0KaHzx6VR7VrLk+/7bU8Ot1U9f249qI6Gko5fk2F1ULQHMcn+UQS
FdsitrUrbknO8cyNl4PLQOD5kPpLX45mgPKhVzntcDU8jmYtG7WNWsbQCjviXEz7
cvMrsnmCPsw5HJttv7z41YhY3krNMfNNPQHaSIUJUWVTkfTo8nh7f/NBMkL442UN
gsIg8cd23Fo/7uFe389pHvyrU3Gqu9LOKqwEchkj+PaeFSADOjihbwQ8EeDH5I2z
r1xvr9Dbow5A0q1eHHizXjFin099C4Zcp4DLjHmE4XFl350ZyT8gT9ACjMPqm5w3
hABcT/1ld5Mmgjh4Pe/yyC7Va44fLwWxkjC6L2jheV5bdUyDEtts6JYltxutJZzi
CwqoIhMX5/Yqs1ELVLNj7hprLnD5/q5ajT0vpVLmo+GJ47ZL/gzqy2Osl/snfomE
dXpusqjH5lV2l8OaTjucszZS1ZeNx0Ub8447DMNIQOqTu1J/MS+33N4HxIpi+CCj
bFrSY/k354G4UoMux+BOuK8Xp1Oo4mXccX6Nze1q+1w2hsaxAjVzm9mbCXpB1CbO
PtabJSj5W+G61n0BxYGca+p9MKLtMFk8r6pBr/7wk9cVUNhl6Emmjvc1HKfLXuLW
UbwKKJTlw1/3jhgrW4ZpP6ePV9XfBWp5xak4rbA00Dme2AAO4b6ej6kaLBsFwy+y
QtFMumv3yHjLMscWMR28HwYIcB6uRjZ28nT4/4+YdMh9GYzu66cCpNwlUW6MU09p
+bb9joIdlZD8eipFdVjpruE0N3NHQ7Xp2/rlPk6NaTqCABIgkatmoHtaDD45ytiT
f1Rc9hv6lS1u55Ug6PVLcyhuwv3tyb6y/TKK7aazLBEY53R4BouOYM87yDDv0HbQ
maiHKLKi7hHzlRsVqOnUAgV1Ui3JTj2fvcik/BX4vulnSrTuFgmV2PDqHWGT6EWe
RGfBkeUzgusE2q2I1So5LxHt9JyJxUYFs2FBiyhPYyB6rJEDqaOHx9EMeEeYAnxf
bytT1QoBkKJU7RGGflOWchjM1Tou0sEwWdNYgaoNM7qa0Vu0RsSB0bpf4hfgzBWJ
5z7z6wtBVyAUqku6kzHAa9qOEJ01uCUaIyEUkmNfNybLy9fu4VdaRxfVg/VXu5+I
ZjPSKaO2x3XAaaX+Be3rHXMQ535aCWeqvWQeQEzuiidpdwYZGVkgjfdzlYT1drBN
vqRaCvUGPAtfI+uBpseM2UquEjaJiMTsHXkysewTmNLz/7W/nNyseACxxwzIQ1Og
Ka7rTiul9Qs6eqKS/cjGwVd1dBxWTTVhhKuz7anPccjwVjIPRt+wC2A2mtSaKPlh
JyKJMadEc3bixBC5Tc8qYO6pYhCAxPyGwbT7/PIBUo5DS+mk6ZsT2XOEvCLLg9kK
TZvNnXEfdWOqUOHWVHaXgaKomh+UPxg+SX/Qbqo+8x/UxARUVG50y2epDVoihLLX
7Q0CYt4+NRLLKfG3kEZGaesEJWaLmN0R+5xM0wfSXlz96m31aklFFzCKfPip0jnL
kGYNpoPHWI7ljs+RalnIMpGtSLpgiOpxIup3zn1Q1nw20jbo6kjTB8phTHlDs5ep
F1afqwkGdvvct2Loe8l2ucMbXKWaIi6GsX5CYs4TmFn0Qi9jnNATVLuZ8QVKqPDC
B38vPyfvaqzBLK67ZokiN0HPPapZlZ3cRh4NORYtwNcL92QR7syCjh6foitIR9l9
eaNzNfqzWN8nxhed7ObaCW6Y0cuoj1xm+b9jwKsA0bbQeSUHr7g8kvtK0CXmHj8E
TBaxno96iX2AQ9H25SlrsXXlx7/HPDnIEakW5Lbt449UncmD/yP9lCV0e3s+i1CF
eyzNiWlOEmkR1crCG+AmxsQScuhqSQq1kqLDPmd8iFfkEf22v1eMBwhuQ5sYQgvL
QgXxxwE3f5hSjIEUijAZU5nvaM84s9IC+nJDiKXimV9c/mxTMXdaER2JUhgBIwCq
7vFwsTYEpOV+z1+B7mpKlcjIZGgDXccrGlNzYDNNm5GZBvPiHtbMcmTknSzzEeCh
T6yJdEKTG5Pkc/akx+7IBViiDtFVeK9aLzFS59cvyrQEYcheqNBbi3ZS8rmDpYrL
TxpckIcDXfDN9Bd0XOixRYZqcBhtUmgA0FditWLArtcVO5nmTfXmT7ZlFMUzPPww
02PrvkHzMSTzPKyAItt3Grh3BOPS9RqKqJ9hCW6QAJSjB++R7hAUdb584Nm91U4e
gWrv6R04QllozAz8q+55mxlLea59aX+J8g+cGFZn8JkVCF7mqopV1LBlkPGJPX3K
zUHmpahqb3kBAEvhY4Q7edlM2owQn+uvYZ5YJK4BkaGMhYrT6ipYjKC7lS+KktwU
Vu4aN4/MQUw/pigMAFCHvG9TrCyTFzISVJFK+k242mdm/7n7kB75/055zQN0cV+J
ep5qJzpf1T81GL9PPoX6JZ0SbjwJeDbRji41d9wCMYrBRpRCxxSnbak3nmcBjK14
QxpyrMUAHwysZzKiPtCOL21u/i0Nh1gbHBzxdj+duojGqif7Xew+Mr6E/cV4JjJ/
dN35JktwPcax7mYpkftGdlo7pKk7D6iTVMxiVy1J1vEKal+AjrTBwjFxtgNYlQpz
Zc0iWtZBCfhBaRf5CLfazmYsuFVLzaWOZDzPhGYfykLeJwGEmG30x5dNZ4TP2GTD
kA9/prwKtfR/gNPDf2LsA/dJddkQ6EouaAzrgH5yNODVNh9uhGILgS5ihaNLTBbD
tIQQqBbthuZ9TB9V8Q8jNSed7ppdSsB/jMz32X2ta7jJWynkDUthF3vTcgVx/Iwg
cQUB7PlHVB9hXTg/9p3fV97VzJNRQYRD0TDVAUKMDGhiEBd8bmIxVcNafoOLJQuu
2YAtRsaqvrKVuIDlQeFlTm+UE7i2lnP003qdj/EtbhVvSB4oUi4qFlPYK6Zp6LzB
S+2loX2ky4IgSt5Yf21D7ExDLznQnLGc1ykbW/3q6RFZsNNNc+LllsXsPpsn8fPI
h/4OCXJUu2d/onvb4NlDPfDRUWYgnr15dQXqHsZqYRbx8Uw7h6wf0PLyr9lJZjDj
N0IzI8jTTra1x/y+J9A08cSrvJt6IlppoTATQn4/u2HAFu2WNezzbP9V0riNP70a
y73k11NzUaZLLTIMlGmIVE3n3V4hvfRsKa7YpvToI28qA6SgRneBSEBcIlJoAI0P
ud8WCp9lA8RBVu6DGa5tk61p9dfv5YoOV+D7QZiYdmCJ7HiuaV76Y+c+DoxptRjt
t3TkHGtpeSqluZgZ8lSPKYYefcAz4vqo5EAC95th7lnjbI7izuH3EXqSlYucn/tN
2lTVwnzL0zT7fqobxn6+FLZvZcLxkNQbmgSGYnBrAZS1+24synS4hmazmT+wS43Q
WwiaFVLG/p1oIOlb7DJCni7z6I3CAvXXVT8iNqEm5OxXHMg3+CBKvOh4hJPBzkpm
LLRsp44jo3GBt721iEQk0k4Wa3ahfloNWcIKJMP3BbyRwvqtm3JeeyrBLXdGJgNb
EcCkQIu44hNfJK2n4Ek79/VZe0HIG9eyUYgI80r5KUmu5DSp5fYOqWmcmMGRE4Mv
jUvmg7JFk5gB2rS2qwxwEa3k8o/PpmnIUJT8X/YObR/o3RaGnag6Qh23snc/BWDK
8hfJ7+shquG/GIc7QaOyJeHHUh5Wqf3I5moy7VlHf/AIFqox5brpUvFS3BzLpo5z
eist7dZ//chT0oe5jKihZ1eAoghqQMLHX0tNpAPb4AmF+aqc+dHjriCbGwuNhnlL
hQfbvtIRt4Bb4U+M1ufag1vvVXiM+4NjgfR94GrugKkbfZlrWM9k1ngeW5Shqoj/
x1AxxmnpiPGw1I2D2Te3SASkCQosSSs2qH+tiSrM1bv4FnuJSKgDSTmqldXmhtxZ
L0vKY4JDrh+/5QY9rk2sBE5VdXEwB8elk9F6txb04twYgYnqnWTH2R/ySKB7XX4j
S/GsWF+qeVVPzmlovWxV3xIwjNCKsM7K5Qiz75Kdgb8+SG8mjC5SUJ77GH11bixt
4fiWvBxdFH1evKeDP5lxGlR1F/lDJxt/5GbZQ0oNZKbeu6YGlEXNORo/8ihtr+DN
no+DKfQTI/SgGTiNzNva69FKK7j+qLw6N5UIKk6KSrZ8uwCgc7yLXc4UfxLD5yXT
38jcIm5YZ4HaVhYOp0+hPe7NVGsPSz46p0e5Hd2yUC9afrywlwvrhLAzR8N1xOWT
+gGz1UWLf2f23RlV/Arf4vi7GxYQ0L7JYTuHNGPRgLCz4XxcUNcGK6YTHRqc32iE
htU3xW3eA703f5LLc90aMuh/MN9cSkGrNptY6u7FuJ/nwonGX8wzy3HSKyssepOX
Wj76DVeLUnD/+0UyAcLV7Bh3C3asnLKIE1scUR1//PKNmSlR+QVpO/BVWBy2cl+6
ptzLwQtjWApOawxdtXdyQy++rz58estzVFCcjD4l8RgJdukC8c8fajY97rjiweCB
eac15E5Vbg0ExTKVv+ZJvmvW4pCihOpjhqn6BHZe53ZnYOYtwhP+rRYjFkqxl4cc
izkRwcsmqny4jPjhvEIoPJzSyAsaSgqotB39jnZBltZIm9DsR8n3PpoHdChnIypg
1UzywultGb8igGPX5aq/iYNTsgpzTakqBi1NclrHbXPb4DSuGXYVZAQe1ONz+ayA
WPo1t0jspYK1SOSUyl6Kr+X23XXMM53ZAjH2GueeZobgrLu77KGiCt7DBh71bROK
t1oaNUtaeEfjuzD+0nMB3X3NoWjtXVtTt24IIWedkeB2zZ1pYVqHrpUWOz33TdmU
lv2SbjDG8s1qSWNwTt7NuWN3b0DyVX9zeN9XtuOb87g/wFG+2/V6okkzKaP2OeTq
Gk3sEoHCvRqBpN/q7MVK44M47q9rvFHz+wDVz52GWmokO0EdgFcwrPOoMYW/l0O6
b7hhnMbosa9FjsCUjK8Ni5JEsEIAwHzziiQTgTaarOrzdG6dA6vYVVnT2aTFhziR
/az+MHgNdGE7Z9p2YnJTZNZqmBFof9iV88gyKjYRveAoxl5ZFnd2qOHubtDTOjd+
OmCs4RNBcAPscLYQZTIwyVqtd+lVvhGZezjvWT2+tYvD2UgW9cKQ8rUg9zHuTHsw
T8LfntK8LQudemdK+Bv0DK7BlB6VlFVlASxHS4RSWBdNtN5Kh2ZVZBz72W4OM4Gm
IlEvgO5hHnA73j3+XzCmBBXbtu9rRBUZJq/wMniVf48Affz2Y7uh5CxkWgemsCFy
SYEbtU/ihj3wwmJvGuLDpU06QBa5wFAaFyorIcXuOEp+8BcSXgbzwFD5X22DVdb/
v8x81n6XPhf8Go06YBZV/kS8JX9uzgAG/fvn0lTP9+79MaNqdVzugOdus62MwUA8
MC9Efo2FgagHCAjyZHBog5Kf+8sI+V0LITu994HaxtVYHgX4rk7Dis+X4reFI2qz
U2z4/Shs4Nq+n6orVi11F80EoquJXHsKvSZesElXMMM0RBQl6p9UUK06aomI03qi
AdgJ84Iw5/0GfnHui6t9bJm8mvoV5Zf8rWBDRXEzTvvjjEVE7hhzlSSg2OW5t3al
GQ4MnR7WHpux7AsPXjR7AWsdYfJWRmR/ve54RLS4p/wJb/C5LLzYGaarxs8EZ638
V9OIbRYn7hdQuIOnK1iPhA5gZdAUiKyNzaKiFbIzxdGXDEiCS+IMpNpUu9zFkQbz
P+gW32so2KfL6KlNP0SyZFAfN6pdVw+dy8Xme83x/uhZ1hghzwInM+0RHFMYrADC
LVmVejwxIgF4/UXLtAW717XoqJw5A2xxya/FO2Ro/sYMDHljTM35Kp3834VUsehC
y6iWshuMLf7rM9Gty9ZNGFfTuCLtPn8Hxmi9tnbJjHpTAX9WkGYGObHRnZ1ub+qh
BDgi0HtAC+m0CEIbhx4aFSez4LOUyp5IDQiYCbfs3FdhKdJRZijwuVve1ctya9qo
lgeARoYsQmvTy1s0XK+ZUHMxByEQr0eudhWvm1l9xflblTu8zAHal5YAtt8r1Ao2
YUy5S+Trw6mtMaY5e9M7JUtIDY13rMbf1o0z+zuLiP7Ouy7ZllcEUVxSmWCfQd7I
swWRwPG7xyJ/0Ty/gwSVoLOUZBiMe6OPa2aoBB4EKECww51QQONi+lxTHovf4C0W
jYBUp316MlDiArKHctlr/0aKKOM9gFROgZzMH5IyLE6QrPjhSOQz8QeF+QzVMHgl
EncxrN584gyFDZ5ZCTmKlyLouGvpwvJZTRDtXzx9kxTwsVMY69HvIbeneJDZ2Av7
bZM8xPurGBI4BEs8Iv2I9u3ks/UJEIU8fQwrqDAPCTFBuNLVD7rdpC8mbDWiGEpL
Mi4akzAlKl4s3KMXx08NWUH4tK8RLlqqOxPwAOLFqhqekjwuz0Yd9YQSxWuWsa23
GCcrdkVw8jJCBJY9eWXgeJYvkR9I2qgYkKFdIm9k8G8oYbIjjVzJ865NWYOF71pN
vl+g5I1O0E0yFY/c/rR7LeSjfFYNuWfmWDWwC/LGseI6IUgkanWa1jC2ffckdvFx
/PVbukvJOJtcE5Sp5TWa52PiU/92caAniti3fBm85YCj6roDf+kd2UNuIQ9pYW1L
Az2D1WCmzzPO6rKA2ecCS9ofhXCfGd1jBUb83Lx0uFgmOM2ikZiur93M54LWISp/
6n8FO8lKYbhLNVlYZn2HdiRbJSfTpkBa8MF9xNdV3OwIdCyN/brgVShA9Z27dbYy
c95W9QVR/LXxj2JGRnqKW7WVapCMgGwuhhl03CFMG8hhpLKb06B/eejtKr7Tz1qt
MWEFppPEbWdBXM/4QaGFMQNbVxDD2FJ/3Q8b43HOsOxqA3/JY8DuxmrADmidciCQ
7zqCHmC+ssPD7HKv3KeMH/+WJoKGCgue9NRal3q6yUGnyGCfPI18/vHaejetBHlQ
oqWr1gEJX0O3/tt2nrGTDw9ONyRXzHG7VzwQBzY01VNb1F3+7UeHVqi9I3w0THxy
dDxW+THi5VQ9QxYwvqlJADKMlCe0DBU2xsn1SgcyYz7NThEnEWH2VtAtLqFkk5CL
0Efoo4AHuJwuDzoSmUAgDd1fFdrkA9WeL9To4+ahaR7mH7lOYQWdLIWbasZJXHTe
CMmkXS5AD2brXCpmfIa2iHlh9xXtgwR1e1LpdOf3ZA2USZuolNVJMHcvFSU6EUKD
diVtVQNzqJTdme1uP/PwHgznoWBYiCublsnrd2NkIlQQ97/S+hg1SpG+oBoP5Dgk
Cd75LnjGsei5Cqymtph8grkgeNf4Fdwr6lY7Z1UvijsuRW0g/b953FJgtAGSFXlr
5OeTueTVhn7Y4OI+hroxdJzlmunB0SmjL/uNEiefoyxJdvR37LLMjFDCx5aSTNWI
reL4v3tRmhj/Zv1j1GfBZf9UEW8ILfRA8I7QxR9hbuOgYNGhXPDBKSShFIrjIPir
VMKtRMAb6O7Ru1pUnZRl/IRnNWcKwU1Asq1b58NkKOEWtE6PHPJ5Z5NSYJ0IQOuz
S/PplDAO2WYxTgv/J2FbEPsiuoC8RL8daiVhjBSJWZVqRBMVlJC6kJziRXNZbb+L
g/d8pyOTDcV/Yg1bu0TvZOyMddZQW/sI+4DT+eWi09cve6nfAteST9nJ97jj5/aU
E19kb/Gc40mUGmTl54WmqoCttlB0HVJENr/xVlWR7tOaRY1INmXVKMCQpPd54Y5h
v85aFW9OqTQbs5Ogkr9G0BmvKdKFS/Ev8szMDAS6xvzkGPB8Lep9/34eink/WQ/E
v4Ehaf1lrbv1yLiYq+vOzV1ahjyxC4SsuqXsmXaBuBTf2GVo3Vm3DtXkPm/NnGtx
iyD2BGa6BkmqkQW89SfI/+Gijh+BHmf8Txl6FDbg+AfLl7EFtPUyVX/vQ4wW+Yt/
/pmBlC+g1bYHybyy6NCuHvPosFF9DMTZ55krMNsE9mSeCxjAxwgarDDXzxDHZ/TJ
6r2CtfM613Uu5Os03EtXbkXJ4QXuNhenpIqPmNp4jkfcgXcdmVNwEQLGGqV/jkB9
wutjnkPaUsvQALbu+B7jm9oFQmdQJIqq3PBzk+nzlcDr7xmIlUST+bpkVpRr80BD
f6wwtvU2bUgG9ZTww3RklUFXBlpbE3+fSZfbHBA8Mf3b/qYXB5DT0X/ggCQOytUf
+/wsUzr/e3265YUm9G+WS6p1Xb2j6TmY7BbyYndSV9dp15Ph8JVvTpPC7UPZP0bf
ayyad0k/fRJQAV1Zz4iJaoHI5qq7XhQ+O1uqWEpXstahQ35rYHUplGPi6ZM7pN/7
3QZOj1I4q4kYqOXOZX3nyPp2gS0vwqVv56CIkH7LuyM61QKkGkSdGGe+4kEfT5+P
JydWy/DUUtu2E1+w9PZxG9bc267OhLTQEDlpadVpSk92WxPWl+bfdQz9cFBZaahb
vdcvZT5xFS0nHfB9aOAtGNoFyTfuJFFL+V91dhuuH+2LXLPlAHX7iWN3Ci5Sx9g6
4/zdiVBF8e1PHwKomQHoHr8TDFVchkX/yBIDVrEQG+qvw63ol4TONMyt6TlNBL1r
FMXslqbWbHHsm1ka5YEqoMgfnc+W8diRIDGfhWxfx2JXLfqWfor2oycIqx4mDSAm
qMIOB/vlffSuJyjhcXF4aMOh7RCCeWceZMe1MvfDa/TCW4tbpZxQ1J7Ozo3mZGHL
dIr7y7QzQFfzeuZAjWrORu7Y5irtWvkN2XOPJRELJSsLO8QwFE48oHl0heqsmEO9
zhHwKA5N4IOyI4vzuQcrudn7XJEv4+K13gZPpM8qQ1hbtTcZVMJwYT6qdLs/ksiF
MeohFPKm7Yl9tKdbATWoZt1fpWG0NhyNuQ3xB2tZm7MbKZax2zqtYA+u+Z0LGv8n
/IlrYDKCE3BfiWXbEeiaTikNCwh/XVOTvpR3EZNRqNVOqySja6RxmPIoQCJNdfg+
e1J/G4OMQHC0LgkFgFhb9NMFZmWo/Mgp7KQsFQxa+mQdbfuAUL/2mdg94WVqz+zP
PF0Nzcw/SoG8Xj8q2/X1AkRugcxrmd7jC3iky+kjoGBaURX3RuLNcsJr7hbdEqHS
zA2dTaUtkw1ondc2/QFALYG73LISKkMHeWwUgnnxpNGQrvsPrclDo0MQ2m7vlwdu
dyVe7GCXADkqOJqFqUCsGMOTkQODufTIOt4orMpsSJE6KL7cg947EsAr1x4kPx48
W6DQLDRGyHubWAnjnrZcixBycct22Iwn19VfABOpfA1fF9X3ZnwARpJE9Rd304Js
qHCicZzcGvZvdJ0b6MnFVuQqxbKDnB+VATeER1naZ2lcKotK1m5b6r3A1WCeE7DD
ygcV/rVuNsoc08e3WEXB9H+Dx23vb7/1EJe0WCybZt9lHtkQFoVNI0UGC1OhIEIa
sDoFJtCZujWQv8r5Ns3C7JEx0vxBsU94AhTxwzWMAeIfMObF5khYiS+ufvij2EgT
zQjuJZnccj1Lt4VvvZG8yGQ3SMfkPEaSfzVjaKTZLMsk7Scj0o1E4hyRt1l3rpJW
ZegCxhfq6Lay9fR3/icpPTQYIE/UyEvA3VgA95JQSc/be4NdTJ5Zm22DSg+2P/2j
DXngFBWeR/eum/wxsR/z6Ok1+ebcoe+ewMbzoiVjstSTmwVzIZct/yfqAOvtKO9u
MNT6eoUUbuQvOVa9MIF8q8apI1jEYpg7gHWIBHbctEYEgbp2TxRUlDEMDYRxTpqp
0vaIg0bpWRjXIC6YXEr9AGDX9OzYFNfPj7jKnhaIh1z1U9yJVUu9qG8ANjEgT3rA
WWDW1nkMJrVcm13ypFPN5GigmG6ZDT1mqP9TKVOhcpw0HLo4WHo6P+tvo6Hkz5V8
KAZ4vyqXM3nChLLg+0FiYZ2nriNCyCUF7UVl6SgAUWWght7TWi2DYEQi4JHjW8tW
Wr94/7pQATAY12QRhJDiNI7Ih3Y6DfHmdYsss0DmXPAZ2qgPKfP67CY638VUPJ6M
8s0hd839SKpfJiad+91Oxf+Ty9UpmKbZw/Gwd796e2tVsVC8mliE0GyeXmlNkCci
22WXcN8c8IB0+texkrY4PGa3GGN68X6fjMAiPW7EH1qezFxy/mgg9HQp1lgHFdDY
npmCoUSCje7VntDRBVVCC90yznmnn+Gu/d8fruRFbjyGjZfW17N1IHXf89kehCs9
+Lbq90TZZs00zrwWTRhRGs87d6kF122LOY3NChafFsX4zfis69hR/SdWx4WtA5rA
wgZKWLB9DK1LAHrgrsNrrpv32SsapIItZj6Mu4gxZvVhFH2kSB+76Ugo7gGsbhWJ
WHIck20jCiBPtqAF9imAE31jFUpT/1GIwyNLrHw/Sx4JXP4LcrEfOASYMq2UNVIG
H8a2T5W6NsAXfIuvI0/cvZyaHjJTn+MffTM0Yj4i8/dn3W+VYPSqoswLil3LdDep
1h5Gf3m2HWLiveZrYb601enW5c4BiFsuKwFeDzdBi79TTqWS40xTxQbCWyfjwdh5
zyRYK9JxUdoizSPuZaL/nT5UjQSNrqGyf80ABSQ9Q54SQ5MveQyMXLFhCGfy6mHz
mDI8NJMA4RfEZLy6IMKNS9SwBFI1IBG+NEt6LtI6aMdVK00lom/Xx87fH/28qqy7
p7G+iitBATQyVA1RavvAWZZulRtta0eMAUelHOhbqVipRR7EyngFgXWKBlmTJxnx
dlvV2feWEreh6y35an+yIX3nRHZ6A6gPAQaunJyLWgixxV3eDDe5zePUOuVU+mKe
HgLVchFg4CxsSNFSxAPbUSfNFc6vWEsLyQ6X5QlDg/T0aWEw46cENaA//j3JEzFj
/BqfeO2u+oJFija8kFGC7k2TVt321dnELgGAaHlo4sTWOuKSkfGjuoNb4ic7zNqM
ZA040e+hlzgNGcJhMDNjqdpAMkGg+/ccsM3hi+a5SaaHTXVDKQRgP4I9Yx6gDPFg
6X4TYrFj79fXjzRBVxwVZO4IZ/8LSmXwVqx9aKCYqPL9KdCYgQ4BeVt9mYUa1b64
b+Pzvt3FKqWjmjoj1G4iDBkNGxbNOn9OI3P+XOa9520P343TjeM3D/v1tgvqmI/h
YyTzepEFp7bRgpbXKw7zYvQGh6/RMqZZG/gmaXqSszT/7rF1Dmspeb6nbcYiiNJa
V4cTC8vAR6+AG6bqD7NtPHTiKwfAYWYt6RpM5EXZzeP3ps2pB7wH5r01nChJTMGj
rMZJ8p+Ip3Y7bLW+UL2m0uERnlMw9FkrVp1HS0H6tsbhQpeT3+XqHv5lSsFgG9F4
FcyCF5FD6fwdSIgYXwQNb6e1XxfeNxSl1OEgWy/7eb3u6WIiY/Y318832dCyzHzQ
/elIRXn/YJYTat6YKMUiQO97rNthx/NMVguHI/lo9/x47bRYIuKFk126Cc65Mv/f
yN/i6JnQ+5oy2KOLGVUXqQGUC5IOjl35ujh0Gzve4SkBOJviOR+Yso+dJSxDp5le
VjtHZgdBM4U6et1AZwwZBmWhqd705tzs3ZVv+oOr97KNLXIdTeg3Tl+UY5uBiuUI
6YcLMbN66pgwEP9J2VFQsE45W8l2Y/XXcbjiLeqQJZEEwMCio7e2H9Gb+HkG0Wdp
D/AjYOev3cxGSYWjcqfwYLq600ifkUzba1teugljlUFknY5aZAoW0ufzgmgBSU+c
FvsJRQ5lJ9DTFyjryeHKXybboCGK0IgQLbkN2trZqi+MLYNbBNnGbDVkmUoCQ8v0
v/nl4l+vzlETBPhoQj0F5e8f8MszgigkqxhijanHnQWwzClFzzWKcgGVFYXnDbJ2
k2f3tG/ArRdNd/mlrloc03ZZvnEkrwn8eVrK2teizbsMYhNeh+gaglZVkDpnGDaq
jGSWOUTm6vuXUzXVuB8rdCqup88Dq16aXsWfCEU7a9OoSVr+NBInVyhrBX6KPxCH
eO1pcTzh0IbSPdb0NFugGo9YH55e/K2i3Rjvb0mCObnLkEchTcfMGAmYO83NCXdM
0VqkDQkCRBQ9w3uyWr74d7kSbqQFqNG17zWzUKt8F7XAasSXnzpH8VzqI62XsPmL
r8Vte0TltFOrA57stQ1oTLb/nkAAWPjMALEi8/CRghmU2Xd//aIkTBS72Qm12gwZ
oeHnQIBIvGcNVKfY9vAGwByy7lz3rPy5w1H+Il7GS0G3cu0dpX/nbU0whGZio/2W
LafownjLdEQA890OGwO5HYUttmxYqdD10PYzQsn9CRqMifhT+GbHruotWd7zSkD2
5tZWy0o03JPQebAOf6Af89bLxAlolCb7dNpxueoy35jRWKVdKKqbh4V8Y9nWNQcw
3yHRWbed47MUq/Cpf3ksl7yYJrSK9GJ2yjIEjviBNGo+mpLsC3jChcPYPRSsee3c
RvPsochLGbaRgR93DZEgy/kHtWrtHa9E+jFzOLk2WJ+WfrU/YpHBkfzhoMuqKfUL
fR2dSI5uO/EQt/W9UeLOrnWCNFNClCLgtlmIWGrDxd3DKv5isiYyGk37MS2f1bEZ
J5PVV6Pp35BkDZOlA2KcDqosI+wVBg3pFGb0VrhMWGDSXsGCOd/cntrb3j2PDjDd
84T8Fsu061eP5+YJXfvad/FUC/rLvus+Al9WzRxmWPN/SYAsugV7xvskY3661oPD
6GO88cu2qo9a5kGwbmKXGsnJ4CevUw9rAH41Jd8XGd88dr18OqV7BGjOP/JUjfVU
hi6qJ6QK2HJpyPTCexXmfAXbjd0pEzmbCciuP04qtcNOoH2bU7zKnAIZGWufjiG5
YAj0mHOrrSMsWmVY4z8zDaNZxD7Qbh2p/M/kXHQ42SQePqODNy8PAnHhLNp0CemI
io5HrGQoTkfFisBXqwhzAKSy4uq0U/WiHxFYzRYv5qd3RgkBu4bONLP+LrmctKSB
gj6iuHW51qazh08aDOJejbpmHhMfYBlHhegqfgMNieYgGPrjFhcBsOeCNQD7qYbh
TTk+4wyPCwP2YbvtyHtWgD4awtmHyiOoUvsvHfR15DQY0S+MUJ0xruX6Ixtyp1zm
vIc1njo4HLjiJoXbz5s8FDCWwaNH8BVoLwwGCW0YfVC9t6yQ/ryKsV5NAlxvUS8R
jvqgYJU8/vonjin3qkbhLTdlAFmb1TRqTPlzrWQBRWSDMpSB7q12Hv8oe3MfWmjU
0+n0oI51Q0JtyX6IvSCpzKXZfopI2jOUlMtnbUJR3AEP75dRfuvfi1r51uoRKw6H
gt66YtbN8jM481OL3eqEB65WU9h9PU6PTGGkvxE+1dQN5adwEP1KPb5n7saod690
7402j7Yj83RBA05qDd+d+medN62orL/8oDDFTh6RxHHDlsr7iezmU06mbJKAbAbV
k9oSM8jsPmL+cKwkZf8BnT2f4jWD8f9Hj1fL/Q0QMQ2o5UyNyxYcBsHr42sNLBXm
pWzO47+E77JtZq4Tg+/f5FfYro44nlf6xXqLH2UKNrtAu1oIDWt0/QXQMPMrlwTw
uI/n6Cawipx1UOxHLe0d5TfSZPb7N+VnQPTiLJbDGKhbFCrtWVpblRwUm9tP59G7
cdSqo3uP1+Cn9Ha2I2MbwsndCOAVzoCOK/jBlfpzG993d9w5HhAbG4/Aa55XMNbz
YNUSI2pe4C34X3s3O3NAVFRZdNjCFU880xXj+JUWgMr9pvCyZLeSHabAT2XXuR3G
mNUzIJSsCbojevzXNR2iGSVnp0YMgwMEO7SQbkHJDHnQFPXMxvG2fhrScLV29WCc
mdDigIpvCiGZfQZyx9JB/BJJGQwILcyYk2lomjDAGmIvdkI0Rje+ihFmeEs4SVcZ
WIYKjdpgAGXA2B2f3zLo1I4quLnUgcNPFunykfrdv8KlkPyY2Ut18zAp1iN24nMW
mlpAetiH2IlnfTM6+s7BwjWzlTq7DgUZ6IK3j6McfMxUzkWdMBIuSxF7uZkDu9Yd
7WkCyYvQ2c9bmbzm6Fcela7zAV25zMlBNjKRGVcnnBWHuo8y+l1IqzYYwl6j6FC9
TzH/xqN+0olGyj6ktcr1mWP3Y5VJnS/ZKjhJQJ7Z+vjEeNTrF6wn/MHVy3FOvBir
uL02t1LmJ6/p7CBqXkPzzyySsQHRxxvfryAr9MaYZPyABIPqq+gAG29E7LSpgs0U
6oYObh5XgNON8vsA2o9gwZjBOgoVIuMkg2q/JgDaBAORtKNslBLT4HtTPk2PWdZ3
2eY8VXuQwuStnrH4CmA2bYOcR5KwOd6yeTDW4ksOFolybQxA8f9v0af6qXRq17zW
iD7TspgskGnn9/MnJlEN8apKBXPu4x4DTkS/fluN33id5Ts9+GpzzfpM9ouslypp
Yev70WjVjn/4s1RYXUD8be4q+yN7zXFOsz28xBGf3EoDMYCa975GGlU35JYzl13h
qMyVWWDhA+SjKlGKZ7Js9Aa023jLYOGjH8JvtWLvHl7tcn9vYEHQZAgqJrJzzHAA
50+10NT3l7f0Lbor7APTCsZCkcN8jx1F91bt4YncvKmGVY1T7KKTSwT07BOS7DfS
ZAwKAs02CtADnbsMjaPCt8SmHnMu8cfcFbbHp8ggFpb/wjrY1HnqB59BepeMx7Rm
wY70vJOh9cVuu5mOHXZcHdQOekpFrbdRzuDfQKjXbr32ZfbnkgHVb/ie6NpbEx/i
gkUduunemDDxDy7ZCtwamNEEpB9enyuB6Zosia546elrJciZkVLSiyGp8aVUTcuO
SBdTzfIpARGFeDVJnXs5JiXrMDJoSo0OJGsLEUcBEHGMtvWgF2WxSGgNWJQ/GTTM
V/pE2Y4pvqpjydMwq8306I4fdYncYp+oV0qvYCwLgyWltpd/VmS6RGNgyGTMKoB7
JSpTpc/rocuKWUaf+wzJwHUR6te9+AEA/OrMK3JU6tSnZRo2OUmcSvh87h/WEgeD
kD9jF288CEJwNW5RczZhf/HOyVg79s2vn4b61LAg273gVjc7GwJe9lMkNbAEHWMj
l/sP+c8zerWxW1I0lhsoU/aZEX/jH/WcDjmDpNY4aGgV25raqKDn+Ony6QBdn/52
ED1cFToayPVujXwPW8OW1TjHrmpPKElme4xQclEG/Uf92SHhyxGVBwQWBVj10ce4
DIBm2HGqzU7n0EInX7P5dmTJCucSlv+HmJK7sLgpIKDqOAPcnjA+/tZboMNeMMU+
6kONQ7jimguecSAvkG2FQGlj18c3q7Va2OnTzBXsIGVCFZK1KpnWONMorqIZXA1a
1MLPAc5hb4qs8Hp0mL9nKAYHJ8OIJFV00rJuaZQlN853w/kwyNun8vrKpZ6UjfO8
+hwMuf9wpFgHy1CCkAaDuTl2mmau0oqYIt/q6yp2pouFGXKqfxmW6Kx4IproHuz1
ISNbiDSCoEnIUA2Nh0ep10GfpC7mBaI0YogwJ6NC+thkofEVTRafmTgOOs529EF1
Eb4TJardru6L0CLatjjF7KFs3jGPWQUGRERBo1J4MaFIBscP5LsJp2vXjpPwDJRg
ZgXe7665Uh79vrxbjTr4KF+dEO7DHK2qdiehRvq/Anp2V9Gx1S6CX0lF2FuDTYxm
z9uhbPxa06bL01uWC0402bYYwqSz6QhBjfp4keagKkpKfJxxpEebjDZ1Pp7PYP5K
seoTkqZHdbuXJLr2jFLpTUNaaXV+cC/iL4xKjcoPgWtlAZQgkxbdCItsR10VN3Q+
NJa/sPH+L7JFtM+Qj2eE+NdAk+Y6e7E0u8PrPGOvgl6i8UohnW0pvIVFqp7j7ZQy
0rHojc+9EHvGmmSapy6yysrRdEdLLFHVSPr9A5BkzjDgpmhYDkUv/APBHfQuYI1u
X4pAzWLPfGLs/X85kpLakhcrpslDiP3Im4WuSwnB4lCX8h7V9dw3S2uxxSvnoJ6r
k3rBLCA0FwwlZC3TOthjTMFKxuOa/wn+ZylIQnskdjCEe0rB3yhyBogspxqxZFPB
UiZ1deYtTjIDDXTWBPU4ZFC17DItiHixQXuTOL2vYZVfQ7U6dF9fvz5gIyDeLtzg
djfmSBfcIweXod18hwsPFlpzI0vj/byjNvlHu8Criu7+IedBbPpAUz+3QWpYhCyG
VSiqx14qV4mfENAJrq1s6OEUCmXDOXgUcRfD4yRXSkcwsaeD2Cp6eodpW1bVWGq/
TzvQ6dlGlF24yNKEtgQTaYG1PHipgc6eh/ncK4eJ8kk09IvipxE5dBlDNzwnI0Wm
Y92U9Mo7gnzz+TgxUmyzJRZzCRLld/6d13S+u27m/lo0pwLGH1mDCu/MsuXYCkMW
MTSbwaQy+Xke0xhKo5zgm+vo9+9Q/sUII364vHXNpgON/Uph0q9Ad56uq0E5S7lX
zVJNiO+vloDq48Q+ST3oq44b4H2j8ydp6Zu/Tb8ogiDOd/4WCUDXelRlVqMs4v+X
zh1FKLFcHZo5+tUmRG8cCpvJqWz8WXtYSS+omp+UF9TiB3oZ+Rfbw0F5EqfGoiiV
Vj4anQLHmKw3zkWFrTZ533CMfTqvN6OzPVCi6pU3RJJ+UZ31DT+YfP/qUQqs9r0l
vlm0D0FzB2zdZ6bPX9kalwIS1RGYXqZp3rYV7w9PGF8fRwwPOpFGcLnkdoJjYF2s
vRJdu8+cLBOCqe+GntD93mVfYr5sR/eOV2AK+LPSoat1vbjwsRbZin4fTZu1IYqb
GSXPAvxGZVReFwzWSUpsdL4biZcxGKztPEeVXjqM3plZ8O9RdvG6js8CdY0bMPmz
dhZ3ekFaHbh6aZVVcWbfHSCHkEPUIE9G17gEAiGOdiwDblP+KvfIYUgdc5Bz3hSa
QFRIReOP+X4mwVyrsgn5TqJNCLzfoRC8C+w4ZaMVILZWMbOqye3ssxjx+U9uT80c
g82Y6wNZMM+uyHihK+lUKISj6PcLuDsmTow8iJq8wBrR2VUx/5ynyz1tAkJaDoRU
yeGbVlftzR9YCI6MRqsvBoUzpusjunCCVjS4KSwd35ZEP8u1AH1lmsnrnOZFMuL8
NuRNikRhqmr07OCt/N7wOVgUVsIQNT5hy4L/cjo9PTHgDRphjX2SJ5+JiJb3LHwp
UZYpdGz7xEU3ngs4RvEXK4981YnlOUK3lKN+zmHZjCoEL7ZCokqvYgSQD2HnEDDK
Dpj29lo2C2KHK/XeFHow4DCD8HNPq9+G44yk6dWGgFlTi320RclnbcLP/nqPS6ef
jOJj7xWJ1kCpJviWCWsdYoWmNnLaPj8R0BHJJB6LlTjf3D98ZCAdjWejxJ4oBVRC
S6v6NsMeuTUToCIZHFgIhGjXoz8ujgRZo2rA6ZizZxm1nLQNQ/JZ8oACL92A+NQ6
UIcbvDunx5SaKtl6UfxwqWganO2OPtzj/7XtU4tp+aptlT0LPKHNEBu7k1FTbTWb
NUhY5F3ATdmCnl4/MR5EsPKhxpj85yR2ijzuw6yQZl0jPH+1YXJWqCrkn+MVE/4l
VkZQLsNWVH2VZaVEwM3cwtGuS2hlO9eVF9SJa97lpzLV1nqY3+NHm8sifUM5KB9u
DIacsUOjSLJXN/cR5FjKYKXPb25SF+rG5NWwfJUzbR76LQXXzjC1hi14DhmB/clo
0UnQO1DHMx90aZG8FqKsfjTyo4l0ck7aNon64UBWHdNfkFkWsU/XB0tOiXyj7jTD
UsvJglE8IT48xWcfmTSX16XT4Di8FJGzakyuLkpHRciPepnGRJ3lV48ymgFgNEIS
BT1YWTKiKZzQm/zF/nR2xdesOt3398oxAkYrXDwg8xPInH4aC2WO4yZXgYbbD5GJ
rrPaDT11H+pgbMOz6sxYQgEWuldrQcvwbZPEZfcFD/0ElZBR9675wXV5oukEa3u3
4jCVCDDVVPcg0QKIaU/Nkunx7QpNFh3R9QnOij15K3QrHRiyya1mrPPXaO3hzqn6
hkrqYAKAFQuffxRajPcpbYGF5jk+oK+8feoy50qJXkRhdev/6lKrWkD/7o3WVzSM
vtJ5S69DEtd4xvoZ7SA4VnbYTLuLJ01ht+EXCzYHpq+BIW2hTFvi5dy8i2McG25S
QXmyWCzK/JVd/oApbQh3V5x57GYdvRRg7nMIluDdF0gUPE3PmAuFYelFS7rD6hv0
+nkZrl65vUJM48cm+ZKnV8wrOmULVqMSrfuRYAvqfcA2iU1Y7nxSYBRGRnryyGOE
FSzRYDhoMwUQxD33cZBkm19WUOFHwObGPMWd2HEnuUEP5uix/g1IbRuqM7zv1F8V
q3+tKFh5d5e1I0SlVHXJCZmLbV18iLWjr4uIpBHvhBa6UrxCjDmw0MIWLJStKj6b
MeYzEcdzefqfMfOG6Fjm1nUncklBHLP2WHBGhum9Pth1c44HF/2ep6f4nh80Ia40
U3bIj/sTPYVSV6m1A18xf+9M+4x8BrAnp0KG3W7f4VQn+U2etDoCIlFT/qpXmPo0
Gp6jZK0ZLiB40oGI9i/KM3fMThLB4xzSt3XWkwFYCEKydIBQ09TuSXadHCtyW7DG
h+lYIqLcVvJMvashTFW2WwqDJrXa3zANErP6mmwKVLfdLcE8gzXVahjHZOSLSWNw
ZjJ0VXceBv4RKGWpppUzQml+uWya04YTNqhpx0XB4X5rTdmh2oBCA3q4TQ7MAmJX
CPCjY+bLyOMx354Qftbnk3TbitSUVf8xfAa+0rUxZd0ypfLogqAWROl8AtkDNVut
dldX4BX2Xs3vq4WvdTUAgpH9JqjMKZw5WMr/NwzoEPHMPBzWTvlmBaSIy1ybrYwv
9icbt3qZBeKTcN7fvkOI9hl+df+lS2QPGmuNPkCCan0OgR70D/qV1/LDToflZyUV
w3Q21d8+vscCXF7Ok5UI4RSF7enFk3E19L2g+VSkSX45V5HTF94cvvd8p8p0v7Kw
jUzWOumOyBQ6KG3GnU14ZItP5OCQ1buiAD8Zb3lQVXI/YDHNdg+NKuHCbXbB2ag9
3xDw1m1ZUv3ctD5aIeqiUcwQt8iLNgIZqQ9wb+99qZwtGIMuKUuHqYwTAJx4kPOA
KZNGuEBJHy2PyjzoxVFmJD6OgCi6qGNIy8YWt/Zevme9lYCTK4i7QqsqmE6yBZBa
aBAg6q9EPf+niKGgDYn7dQ+VENkW2TTaOX8ofw57dq/zRm1EUqIMnri/Y3y5XgiG
0JEV3dm/R4lLtPS3L8MP0VJVPGlXfb+U7RhelOddEYSM+CgyFesWhZ9gBbPM/r9k
aQ01YlSEr2NvY2dUMeJ4oz8wygksOv+H2ptVDhTonUdRSSmuwGLao0Om2obll0D+
zITeZtazpIHfm+B+gmcDUccYgHJ1SNr9ZXyulaKCuvOFXyoja1NUbiGsgJv+buaP
7lKjgnQT0jpUJB5PKvwU24W7ukbJ5+G4OJm8l4+c9Rha2PZIQW7wS0k5qaBqnYvc
1ZZDI2NpPOj3TP3UmWy7oB1sz1+xSgjt7uDxA45zQfGg3G3npDzZaYxDOPbnWlSQ
QSoZOY57ggpYtO1VlcChhHdy/fNhoF8MSG0r2W8stOi453DQ4sk+dp6TSr2O2FIi
Jd4kL/h2mHh01aXt8p33HJxaHDmjV8QaZE6jgLmrTpN8i4fiJn4qRVQ8hVzUdYmM
zOQVbMPN37EP7PrOXJTb5IFTsQ3JrQ9QlvUi2vvIbTu/iSeMez9e2f5bBzskdQER
TEvdnlaI8S3G1TS7L1nrsnnB4DFjeqyN/Ronx0xi/y/rakyOiI6KtL3/oyrpf066
7h06lbXFe7LNw2qwhocnI0PNlu06pGFuZwnbYRvcOjGZ1lg7XOfH2Z8p428H+lP1
IRgZOZhlwoi/OS1YLNNa3pkexMx3HiOsyhCrkc3EMjXGWDJ91gXv3/JBMDJeb5Je
i33eJcn5dVZD95xpgm2/CWB3i2rxkG6AF+y4GiAzsUoTCSYRtrrsOBaXUJsjMOmM
FQaFt1X8X0gZWv59L/Bm4f+mnyJ5NS9mkEc/m70maJjPj3/qz+dPAh7umA9J5fdp
1UY9qnwjMnYnedgSobSWbW0GBqfW/tb2sgaB6d56jwde9uSbUFkMW2ncznM7MaOi
mRa2JdSOLM2ycu3OvpRIBSwa309jxiz2+IbGxAeQ2ybCWoqqLXgRDQ7VlYJyiaiS
3+w/oolfptEJkk4wHXSDKZTKA06T9AWHNt/iN0nkJTtHSakNsPI4x1RkRZpRjgp8
ynPiVAExTAzdIA+vdvOsON5n75BqhW/DHD+zuP1SIcZ8HBWn34P9r1cBgKrH8Dfx
YH1JVmD08/u/x/KIbQBSBEdCRj3GhlTMWP+ZdzlXTy98fZsp+cnljMTtDU/So/9x
PmkNo0VHNMJw7n8ekf1M9nvLb5lHxLeTTu7gCEtvFp9Nk0v64o5yPQrnhm5jgrv5
WWdepxETv2i59tKfAMyLLp4WyVHkD0hqrWpGlCiTzWgC5sx184pLPMHw0xVSmN4V
jOJ+k9N4JZjL6jWAKoLS9XqpFvhTVoSp/MYH+7gSB3PBK7AakcPNgyje/pW5lolZ
v7j4Hj4muVvkMX0oP+mKnLtjMso/EispY1yylLsPICqPSlR+yy42afVAigCslTmm
K/Mt2V6LTJWQfrxRrYX/GJk3VMtNj+RA0MvilAZ3OzGCi6wgd4i7W/rOVN4qnvOE
1H1C8X7FX/gxCos+IskxbCHo7UxjMQxQOnu4ggzYYRjTHViYcWXgSS4XjE562hj9
Kie066DXBic1ZYM+HK3EPY4as+dHUiM9/fFLpciKywdj/IF2Q9joW+0fWc4CW8gr
j6FyA38HYxpEeIPeuTv4qoK4oyPaJOT3ZlcGB6jPS3gyS0Prz1wnJ/JCZXezzOCp
vUXUJEssTcXaix5pAPb+44A6bn8o/C1NW28oJauLCMD1I3ViPD/+dFuJxZEkLhaE
aOarK+H7vIW+3dj+3jqHQlsp09BDD8ffm0D2NZVg6bHiOpq4EXDKD+mNDb4DzkK9
fFs3cCcpdBpSge3aGQ3f5uUgJCxxpupcwJLGtHL9aZwXbvWh/MBjIYZe3O9WhXnM
M7A6vRj8p/P+duIwUJUy8oAKY83tc3LaAz2ZatQaVQG2hcGZCkz3+yOioG9Ll5Lv
RpsrO1y8aqIFx9maxPaUeqSUJxrKUKkL71F/rlqYWcprjxpL4zvSsGDFMe2jPv5t
XzqiviDt4rc/zPTZgBShfk3vsHDTuhRmGuf/wgJtz+VN5elF3ywXnhlQPYkYk5tw
ZpWp9HPMxGLJP3SLEPRtKeliLlgGitnCHNve3kOkGRzJl9stqHhoRpOkYvwZC6yf
pDTlG6ccwsdRouQyxzsbneS+QU+sG0wKKdqesqnOpVhfGpFhWZGLvU+kwgOspbbj
L+RpgEsaPPoLi8GajNj2psIbF4F4KuFbHWmK0LhQZIBUlfx7VWtx5i2lS6SGIBLS
h3Xa+OdYXaQbI7GwCdlmaTXf6ceckPzfP0tqlzyB1VNmqBpByIgiKRS6aPOmfFDw
rgCmKcu2QgV6Tb02krUoEur8x411sR2m7jScSC/ruqgxJ/Sxr3IM/U0UW3+dfEaN
UnURKmVd3vwkdU6ckK+1XYIZYLuoQOSvAzTffhKm0itrPomZ8gAizj2kAkn0l1LI
CKYPRtthsZte471RG47YAUlrxxiuaswPA4wdfS4cUBB5y5t6W4PkMd51wO6ReSkh
/yEMuLLgJL8NoSvxdOybhFl3fK2AZkCXsRwiFgbiKJ6yjKZmhrinIN+GCNdF9zZs
pLN/cDFjJ5YvKz9G20wr0XH+aHd2W3zt1/SxmBJGmkEimA4YcJlgd/lO4lAZ6Y3/
gC4sQpwRxn+bXdwcAEf/1dNgoz2ggC41vD30gFjmwRNGOhRgrp+Af9M/V9fTLC69
jamFSo2Ok3ajpHsSlJD59aD626DpVcvv2YmTTlX9s7G03JtRQldhOTXm3eAtC/bU
HSJU5dvveZBta5lE+x5/A9jEW0JTM6RnIv69TPpHrz/3z3Vm5rEcFjud5rJpy/Re
eKKyOhOsfspfYmbwR5r7UlEHfe5rJ8t2w5O/skNGYiXYPiDVu2jHRfEhv/ZZ8chr
QNsX7g5DAc6NQgGbqm6rRYWAHcV4jM/CDJIkGVcqI8VnjOZkKExv1+1XPGdIailP
qf2dMtJQQ5hNzIHL9/JgGzkybYKjkPC5gjZYJxuB9VlkOVqZdps83dPrgYZS5K5K
ymh5/pPVK98Ppt3SOIAncEn2pDQaWKH8B/ToXkM8/XGzy+n2u683p5QAh0mPdZJc
F/8glOb8EhXNJ2cHChL/XKly0YRRFwnLj1z2Gh8x6EnF2LfRTaaZEihBS5dZi8or
H3gHJZLGItoZ2dG0QF4itE3aSjE/ar28wVS33/d41pjnQt1Ch5jwYUEZqAKjimgA
xogavgcQalrpoElRPE/bBzf4cwu7C9jQYi44vYx5RIiy4dPSErgm8Jg8BVFucYfT
2Ei9QU/dZLceeBwdd9LzWS/QUkkrx6QscXUI5MWZ2SssKDomLUdWpSL/Gmj6QZoz
5yJxAo7coTlZU35MqtfoJV/fOTbelfZqYw4pdzFLyFveYz5ffFoK2wgWMMRCpOjz
zBI59koP1i77ok6/weUgge2lG201L1wsOhmp+1rqfehwhr7xV7c6kXisdSu0Et8V
d7SeIfXLKUNnyvFgqUrJIoQIyKKyeZLdFEDnbqjqKgtO3hGuR3s5RLj/+6S3POYH
PSPqbKnxHEJm3FUNsYPpXjdE/BhIqVKJOzHWltvrBDmU/1mQ5lCOt0T4DmlK8ehA
1ls8eAhvO11jPk+FHHbBKKpCmevkYXut7mYvtB48HsEAHEx4CErTYiOtnoU/R+md
Oi7eLALwG5OGqx0f/li0di05KR2n0DkyZRrbto0oh9BPPjaSH9N2xHBatwnO1m2v
o0koaTHGQF6khnCV+jYZAsRRt+0NmmOfLzRALOtmyBqlWmKA+qlQgQRkh+5HL0y8
Ebw9Qo9GL/QYsjmKhdwOaLG9zT4zzHXPePk3jJSFoLfJRzSvjsAx3DXh0ApkbnoQ
Z9oxEW/IbfexwDYhuL0rmSBV7dKqglrGVjp4l8fdMhNutHMqcwiIxiK19SRiD443
UJsbaOYZepOhmA0QhuHqYCsGUfek+v3kkY9OGb2p8O5Gz2zco/RvsStw3aWvj8fw
cXqlMmBFJ++nBUoaWAfvPqDyXiNN2jh1D869j5yP1kLZytrNBRIKFSXkLEMcZ2Ac
G2sLnb2jGB5JcYSmkCmT9wewLVdbIfSV6TnSq8qtRDMgTOtLIsQD+9hOvSYMgbdB
2TVDtPl+MCnsMoXzgz8Y0gPuMyxTGV7Z2FHDHKr7pJXyHHxZNoXlGU/u/Zf2e2SC
MGMrxB+ME7OqFN0Wbbkzp/BZoFMZT9SCQNMDHlJHcx5kvg+J2u6P4XaZySEcQBO/
t/P9rMY1Qjt3bfyBQ72g9StwgDx2QyqJ2DRGrrIGZM3gHsSYIzcKqCmBxJqohpu0
9qhxzXoPS2J979ND5ZCCU0Tj1kYXwBjVF5MvW+IdbZrDi/NDervVd5YIL6o6uYV9
DGhFGK2aVIys+1WsHifZmLaI4mE4YUQcxSA5MQcHm1bkQANnA7E5yR0Pw7HtYpr0
Cp0Vr5HgkvZvEARaUobdABKaNWswl4l+QZDPmck9u8B96Wo8J7CuY1O4nFNep8Ag
EgRFMR0uTAhQh2CFeasqqppGAZibsgVc2qSTkL/6nael+De81knp4z1gZCB51kvb
rxKA0zzM0Bh/dmWKmmYZfEORyWtkAJPHp00jCIXqxIZRNpA3WwTA+rkhHDRyLzVy
OkLywcfk3VwyOJ1UfgEif5Qb7/HDY336w0Hbho/lzn/VZJGHlrXqGBGhAiuyzGF+
8MVPisl9JHPloWUViORtAsOHlJ/jMY8CgBQBI+cEhFx7eZy8qQv8f1ea53dpWMiq
Mpu8yoqbOtLsd+H03XinWLKkxYBo0VaK4sg0HLrO7/Dxc4Xq+Jb1WZiV27BWDqHN
usxCs7v/FOCUoXQggQCEyOcruK194kIJ5e+cL+Ok1D5lPgL+UPQ5uUx5mIVWTCBm
GgIKSE4Fn3D+kYDri0D24wSnL81YwwTut5MWQSyio11T01lbd/dq9GUmjb2Pcjy2
Secyv2B+gQjLoy9t2b7+qH3+VI6+jQOhWkNIynTncdK+xzzT1418ctz2W1Ptaz7z
QGTZSTZhYPF5ebRtGI8It1/33VPk7cTs4GhkpdGWANqmvVer6NsLH9UldEV1/3sS
PpWZ2gv2ezYabSxtkTIY/YyWNp58yRe4ppgSIL9iYhLmJ/pRx3Lx4+F59Hfcswk7
G72gwQ9IltBG6uav/v+95a4Uhw0PJoq5u6Mwc4sODL2rhvU5F+UNET9v60E6bZiA
4s1Yp6gAfb1W5hc9IuTMXgG39fy5d93eSUh1D59OTG93+AaCi2DivRZ+WtqaEwxJ
sIvxiQtTeJa+yksUudT5XKq+iiXQYjJJdmktoX9FqKRWXeqCaP9H4qdPicyijYcF
skjIj4af+fDBeHK6YZbOegI/jgemAIrzw2l8ko4hVLXO3NfVsHf/duMsPaTPjMDh
ADt0ErkmjxuhY01E5VDeC+trbt6Wb2U8SSbv7lB0QVnH6t6pyLDmX/2za6TWSAva
6WPpLrli5xQfxxp/u9Nq5k7HDh2NE9s/FfqLsvVHbKHaI5Fs6oFXN2pIVOTsnKkr
PW+fZhuCWLZS8Lcsfb5U/NixUabnp0DrnF1+v4HjBlVFWVM6i6E72PlcE711uaqO
xBVgqJ3xojT35VbJa3xaJfW9WhKkOb2ck0pUb9te/ROKoFG/TsOYwOVNInZ2iwrh
ZCFowQIEijdYm7yl+f5sv9NlqMxeFqDbDkj5/okKH3roQUlFtvqIGJjwuFlS0nhH
IAHh2v+zizNFlLex/NKHbKgwddqI7synDIUYBBWl48cGHnlwZAoo/D9uIwk/uLnY
6vMsz66izraLTYxZENtln08Xntq33kPthPbDyZjeD4rT2VJ80S1xkHKf+R0YgorC
aEJbOcnjUh0QwhfePEHkGz5OsMiYFb77fGNdA844tJCP935jWgwuCb7zTzW48yeX
ERTn/3c3ixsorjNUyVb/pt9kUDTzhvWhHw14u3XqoPY6GddtuUtyux/lDg+8lTIi
vKfbGaAndDVMhJuX4LiXu8q5vv7OTQ6uDg2vGCuK3Oe4hQ82PK0hAxt986DfbnjF
8oQDKO7IlYgxyrk6NtpgeO/VH8UFY2XQaJQjAf623xMBoWB53THIYKUthxlT8NIY
pV1oqKLglZNKCI2HV6QflMKIN7dLicQ5IF/GSFGYgy5v0cP40x9NplKROsCowl/s
B4aXAqI+UdnudEPycu4HsiZKBE9p6ftj3Np2c/yj3832xaM0kyWaMhr76AULgaK+
wPGLLhjnDT2daHtfbTXqC/zwJv5nAWL5wQ6z0Sb7HZQtKkFb2f4bFJop+zlehtDG
4EYep6BqUA0TxNnAeAHJJaFpopuSO+z+cJiXYorMmk8tE9FpejSJ71CCyssejcuP
s578Ea+94XYbunMxccuDgNKJrXjSPpckHCztevElbDCvhXtl+hPu59PuEefgW9VG
kNt7shEKvKme8VcaPpun589LFsY+zKsgVQNNE0GYtw9hfBsstcDJ1sGJc+5WQ9yG
diVt08bZ+nrfbi+kZ68kZmp+e2CLag8KW/bTV7Fxu071qxkJLqlEsnZNUnzoJRRh
lv6tL94JgcIQRKvh7IgSx242yoCj4l8SHL9zUHqke/YHWsXmsWv3lDViVX4EOw/m
RJdC2cTD+QAOMH4g7lv3cPDUH+E/x9jmVh3w1sFAgfTjecZEAJ4rJObUgwXPeFdE
ZOut1HSou8JT3E21OADmlBG1GNyDTAuTe0o/GlY0FBCC8JPi3+B/4xVwUOlrYPsZ
HQIx2N2JtzAprqGya1LhpkHTZggVOkZNh//674F5nu0SfWsuGIUazR/hYEuTC+Lb
TW4HjuDVn293Hd1eVbPMexG8H4tm5tNV9ShqSCgr1rVHYcgEfu6GElDweqR9tWg0
5gBn2jJgQWGHqNmk60LKmCO206bJ/TYd5emqySN7HReCNmslB641E02n+zLnk8SP
lnXxJD8DSFuu13o8BKEtyHmRPkl/+KUrkcZhLJsWBGeFhxAgnCS64omBg1Ch0Lb2
0+eROBMUKil4JIIi1VIxPuuufKrfottTMvXxrIeP0Z8gsTNidHfjlI2nisON4Mi7
LohKVSutyctZRYPInZJSG1VkwO665JgJocSbouc63ajunNWgNyYoS4WfDNFUrs3L
qBnqtNgvHWyxrKzrF5W9G+bu/I18o8lVybdvfteMX/taV9JjizkwRN7N7X8a0Hgo
c2LYM7/nvXbdNz2aMgmfmUh370Y/dWWaI77B3buhxaav9NVzCSLM/upRN3K/R3UP
aOYzmVIZcqVvUHxZcBVTxiF3DDtzTcyz3iVPmc/hgMrnkEki+pDS6NhnaEZRMoO2
RBA0zH47vsQ3Y8YWAmrudqZltbdL5nSc+dCa6N0ophU1NYD1RPO8el00NNBoLwgM
9WMcR68NCKGU679PiOlSC5WjAgdEtDTlpLAMPyUfQ4RAK7N4QHwYnftKHu4YbLPb
1bL+tE5WEBTNjeRXc2eKp6YHsVekL6u/Z/L0zJePToCdZgg8aXKjkg7HD4zlq3Fz
3FmnMLkn/yE5BC0mDDxck9/IT25XcanhvflfgESdyYbr0/dA8SzFWhDrv/41/Sd3
oIG+rmRlZQ+DGNx0XzL+XKYhBrd8PP9klGnEerJJO0pMrewPtHbEi6EwP9DQYMAO
2IGEOAczGuVa45blTLSSBeH12ikMEgd8uiz+YAlomCrnWCJNCpgaeZMWEv8ntxZk
lsUrd3zdpJo+VCb9tTPzMtzsKavKb0VkGFJJIALyeX273TC3xvaV3H6K5/OU8+Qn
mgLcqPtdw0oOg92WCuiUy/jksp4dZVcrf1Gwmc3kDJDKj9W+kAfMKU62e7w7dFrZ
SRjJ1fjUl4ONDUx+PTJi9BSWTFxS6zY13Tptv8rlZ49eUkvtvFtmZQD5qAgv68M9
mlUa0Y50tuP5sTZNeX/vRu2ZcxeRWOkkTxAtuxTETQChKKQBEcvaQxMHvwd1Kwuv
SVldXYNf9+yx10wLZ8rM5NF44ifNUc5lzyPPNlPlQvqyKvECsIy3CBXtYsRPdLJg
RgFD3t40SdDYoSsaJMkmyJ927+G+F2t/p+7dFTkR1YOt1NRRKBKxC3MRJ99WNUIV
xznWWIuwYHjdasG7zR2NMy1dSzhYYP3w+50m1URcnsJPUSE+SZFYTlZbyBa62kgk
hTF5yxewzNGRaXUMaYrSHNxqWX9H2lUC1mAWEGjcY8dh694l3WTXCbY5BWEls+It
8ou0cOm3aanQHYl1ZOVomggr4B/HD0bkeaS6sJpUnpprnDFvYLEiS6K/TkM3K9VS
Zy95YQw52UyVULfpHOaaNp2MP14OeKsTmK9nJZVWxWGbtwGM035mxMRvZpTqr+I/
c9PRTP/BAm2ST+qDoRRkt3JsXtfLbbj6HxPm2t/Njel9dgb2qyX+XBQWFs2NFMgJ
zSoGRwGxtv77+E85qzap85+SsRw6YPhrJMsti9bUYGPb/m0ATA683UrSp2LFq/Gr
mx1l5deHB7cu92M+k08Q7/qPkdtPAJQHy+eY2nRlVv8WHInixGoJZx9HCkYxCw2Z
vMQ83lWRogTy9EXxdtY4vifWIfH0tvIuznUY0G/hw/pQtkF1wwO4yeXOSy4eWqZb
HTFPC76LbC2OdfS0pvfand2NJHXaJBVrCHR01L0m01wPtLtWftplSZFwXXVgU2qE
Xr4aL4iiMC9pyFWNz98Id52kxtQF8HZlYKkqT/j0CEM99SLpkicZ5M0iL1k6OSnE
ZgCfS+pH8OM+y61btNRDpFmfnQMkP5gzQ1U9556Tdv3P3AoyMqnQNbiSsTqZAiLA
xzNpLE1i04IUn1AlZi0YoZ/oP3eKb3dL8H/Ew9HDCUJI6V0BUlHrXM0N9sJdJ9nF
3CrB5sS36PFwpjZpd/zNbNL9URgC5r8hSj+o9hWBwT6tr4jaQuxS9PVtilfs3IDI
zedmSWINmzWUfR9Dg0R5mFsCWidIypvlUOone9AmFAJhIUGyxFGNDPwCeEqdPq/w
sO/7/yWQX1SNIZg+M3kmTykDQr89PHXNmJDDHZ7rj57yBcBGJCvmqgWoz7LmmWHo
2A5sy18ceU8K1Mu+LxhjdF0axe6FES/gfwKiDEuc0S2cutSKBZ8DxGARS04T9ro+
4SSEYUcsCVD4nu28xlaGPMiMM71ucyfUysByY+6p4N3DZJzmRWEbqsNgOi49fj1n
6XHgMn7Pr7V1kNdrZCdS16+xe81PtIDK9GkxQaLDsk2GC9f20wk6/2Ao0yDYGKQD
zibEemuJg1KY9JcC66YCTBX6S7qQO15KzteoEH0jDNR6l6DW6KK+42RjN/OX5MUz
3VdYu3NqpKUcr1JUxFPk662X41hj8juILPmfw+MAXzgQ45XN7Y/b4OBWxHxdNYnB
AJeRcnH6cpQy2IlUYvttt9YBqU6oPTLCTUOIRGrXa0VdHEdvbsB+RuRuz+EfZBUr
aU+OV8evRTjADD5i3OTT/CpNdU+TPCkIeOIgFi6H/yrq5pHBtPozqC8eFpjm7Iic
9EXUgLKRyufb47Gy8wqv2FxxPD5OwsJFfjMWc9/B6soAh/dquplZMSiTw49i22Q/
YJc4FWeeBNZJX5h+8u/A6pH2Bve1pq6wzhUXAk+hMI4Lvwfi46yLOapgdj5NaYIc
LEHh7az/xQaLYskOarfGZ1IgSYCVTo7mJAIr9Gh8DAcC6iCa54g5k1FjjKTiSD13
V78Cf00xR13MPG/RhRakVMcewM+dezfIM6S++fflagZNoSSRHNYf9ULVSpypc2X+
oq89rDzh29c8xOXDcvBleBUDKikgd8t0/26jdO2R2APVyxbxM9KEMQDEzzvcs1df
c6LpeuDAuckfW9Txvl2dYoSojRJwx3Wq0zTZFml1KasPJ3IMDt4q+OEBkuhbVFVe
kmiRuqjo20qzfg+Rwms9g4CBNgFDppINY7N2WrJ8C8R4IIC+/+uviyjr3BzhRpox
T3ZEGEDoSOFINhAsbqr2ZkRE1YDPg+gEtAmlkFk2whLCjvMJD/RDv4i7QldDCMcI
hfcyocootnlKqzK+C4JLjiJdjvEwFZHLSN2PMn4WpMwfhz/Hz4DFRAZU6zmGHnZW
W2/Pv753e3pcfL5Saj0pEkXUZPYdkozUWwcPR9ZDLaKAlPazH2mmu5iiW4spPuCm
aRvbbsaQXgqQojL7rPL6mVJweCvAjda8yn1Bn6JQeccd9BU1cb/fnpYhZIxLkVDa
0WFYcolPdzKbe8rOuN9qB21Cpr9HOgHBD5YgYd1Zgzpj/hneSlpAB/EgkF5MzMnk
rM5pgNxlbLpA5RwxiFc29fWDXVdMop/UV353S+hlHwgc8IXCEspsHQgkRlkNRVMu
VXZ49Y52YfT4Z/opVOK60duD8zlPe+vPjop8nZyaUIB3kSFwnrBArxE1XoNC9Llw
HwoV07p/WCvr0l2pw67hW7T7K0PGv9fjvKYgiuziBG2/9jmEFMgTys7En6uGb1t2
3NDvgRm0WGqVFlfdTqqjssK229IKDAWYNY9RabLDN+Uk5AS5YSrcxDD1NH+z+UTD
BB3dv5u84LHNURzi6zEc5YPcMfHzqn5kMnE3bvGgN4vnz4jo04KELpVqIUe5zf4p
G02aLPrPqN+qNpRLJ8iDfHPijCXjfSObWmZeHRJaumbL2PbPwFkKelQpJLrGV9AW
9FtG4z48e8ZO4WiGJeA9IblGQ5eAOvfhZesvh0m1bgk2ZNTYTisY3sHAZzS7NSea
ROXoX9KrQS6ECoyfRD9RTVmzv6j/1Xi6eN2W7ApWR/K8dnXIW2BYsBwcHl781CT2
D4emspg/esQSHQRcejyonsx8egY6SziWRWxl+v87f1SLk0UnNgNDb7ygxcchYwNW
QfrkTPCbPJ8dHT/zFkAcg3N7n2+B0ZvxCERkEoljUbN1Wg1XGbXLrDisc8AOlUpl
/l7qxkR5blOQP+1ciw9qJ+YPV5xCb/1/CYPnz/JT7Ho8WCL+Z3TK21pW1wqNNR+o
DqWSJ4PFUNVB+ldcvU+5tUdE5PQyly6lDYh4MlmSLvJCH5BzLpZYV8gl7+I96LhY
bz4dU+Xb+ltl8kdcEiPLMK8Qh5Lag54qQrLjv9P5tysuigF/CNQnc9EjKDYHuSmA
wXZo/fLSkXS62ArpYE+km88iM/WnBR7WqFQnYVAaGJ7AqeI+VALh02vLX3AbluM2
Rs9ZI6CJlfqQpJeSPEh0nnP0vfSz+Ctr6l9nZimBZruoxBeMezhqQeBXMOHND/PX
2CujuHvv8GNuZe3a3ZPcDcu/Fb6tC5iKUhk3nsibHVsoGetbPB5G4xE3Zf6W2Sox
OPBrAWYmbJVmub24II7Ow7p4JwNBpr8L6CYL+sUX3LiCMt1HBExA9loc6rYwT/ed
Z6lOzlLwcdsBIbhwcBxyPWYswD8lPyJP4HvRUr5ywisy8rtz+51rRNErw4/MW0KR
s/3GVZ5htLaX9NsmEIrJib/AFmLYVcQdk5rdqq2dn7BdDcbrgYBFNeE/kT88AaFW
C5aOaHOC+ZmiO8Xb3ficAaM4d57KG1T5rcsMIEa5hgMo1GwWwMpMnYCAAEP7/wTf
FHjQeteVFj+rJV7JZ5rRqQSblsN9ArVbmPEmG4uUol+LQgC5XrbbNNdjKZ/eDFM9
W8HWlrMi6k6feYuS/nEiUIgvTJqRTdWm9g61hY9I7SVEXGt1+FBRlMvLdCZJibc9
ww8J5S2a++9DglDJH2u4k+Woimynm3FVToZMaN/ZOfuJgwiPhJyo1Ir7iQ1KPqCP
CG2bx1sz6rESuPKRg+EDHkR2X8C2Uk7Xr/8yMW9XSZh1gqxns/jKYoDDYkAH5C61
konzlYNbI/Cwar43vo1NG8mtVaqLj9Bui4gMtE/Z/gw1cHOL4R8luy3xV3jeQQU6
x+3w3O11kXJRXnIarJVxYn7mpjR6OaubH+SMH5cJXs41jrkan8GzO9S0GdC8FkL5
nnJhXEMrZ4LRjJFd/9sxFSGylWJxK+o+x6ln2BYBaAWGMAHki8rT5urLeB6aHsyG
OeLcf9utdOi0v4oQVimGEpFpux+YdC5ZNsRzBYIZw1owAA1cyr0MAAXjxLdZBvF9
3SDzE7N3zvThfHiPdCcJOn/FyJnIVYiyoY00HJAd5/3e+Uc/lbAFLuOzQciQSgbx
a3lzYj6IaHPLqGCQE+HA7afT/1dyM6O9E68noKgTjnGkt6KoTiLkWz9kLdqVHhex
pzNdT6SVeiahiclDBLHvpWlP7M3wYeTm5Z3zHs246UH/1tEEu85FkSn3FGquZFxG
uqT1JuaCN0GETMCqX57K2fm2nUFrxZYD1GwwwCTOLc0yRzPsDFgrnuN+UgLmO1IP
gsHqAoqOslH64St5hZ8eLciOU/LxfpB9C9V8MJq6V3/lY7BAP1OW8bpdtVN4TaGX
Dd11YKgbvg4CrYatcNHPk/mkbh3zagQxRr1XwAMgQsUUFNfLg08l8xpq2hD04Vtl
XIf1YDdR7AHQNjmNoI/BdCifKtjMrY6D5fhDIxA956nWlbCyLrc+3ur/IYWxG6kI
KtLcjKt3XqwopzcC2Wwl0uARoD9JH0Tbzk1cJA8pColu3rrFO4oDnjwNfUx1V9gx
1O3J9IN+o/CSUBHgmnYwJvM75Jq9bfASjt8uffzyCwhTlUmpmYfTRItsUBm8lmsv
IKEgmR4ncFeYOvI2rHDRa0p6utJDxMdSZG9/GYIbsRYI8rQ0eYprlMDGrQtCN20A
yJZwXA7+YUvxAPUMun2aklCj0uDIYUcrWWbXJ/ZOpLaxp4kBrx5rKS+cduLEbOdy
JFQrJbTGDqymUYb4WP/kSVRCw3SkiBDbqMO1nEYrhe2PO8e/hPVbQ3zHcEU57CEk
UXflA+UCZIsODyltLX8ueklhOz8LEeqPiysW15IcGjlOId3iT02gXtvtSIyzilsj
ZSB3cC8RaVUa/XKHYK6rN2UfZeU0RXca0MsWd23IgoikKWkEzsIkowUMhmChlFqV
mniCb6DjQ6VJP28DT7Ae2+nsaCe66lhmWPZV+k0eBtCBL9GBOgZ6nw5ymelTyTxJ
9XCfNbgW5WSxfFwS71056V6873GI9v1UesOglPmkAAn4SMMr2k1DF6bq0IW8aiju
szT1N4FlAXj3UmWazrrHQ/Bx1CHBT4MLZ4RTpXS/WrAuJPQ77grsVSkT0Em9kQId
lLhD2L3rCXztMDnho5msz4GyinmPY2DT0aQVWQvzI9JwjOTlevvOv7DyM4pIJpPU
byuKsnG2asLSyZ8Jrnmti1cemVwkc4Mu8d8gihr6U3c1obAjGYA25f8HGNDLINpe
9vWNSAnlRHqL8PNa6zsSnrocBgA1iz9y12ZDw7MNPd6AkV1YVFRUv6LXfqsRXYZv
a14sy5Fo6Po/3DdzoCGBlOqz6kNMQllRDrrNsNMa3u2v9aGanxckCqOY/Hb8hPrK
+BP6z3sLk9O6VbIBvpU5UDlQ+uSfh8jx0HINrEj47W+yfdaqRlCymUmBTa46KLB9
kfbYq4JFHHlxdOkQnnlysynyvYlmAomd0dVMyGQp4XR0eovM9QwzGRMdRxd2zn91
MB8ibvX8C3wUG2J141TnEGAVReG4u24rYXia9BxXtHKLJJvBB+WURs54SB8oPNRh
gEc2apHD2ueBd32uKvnVIEFvatFYElp3+T1JgMSdxAkHxvzCpCDn4/OMbCJ4Gajh
eLbwEyyNTJUAtiB7TUBooSjgi9Marx8K7D6xJx1SGXIdsygiWa6YTVeq0rSoSt0Q
NC60ujAom2+SKY8BUsMP2ly+g7pGsOpJyi77rDQ5kXSDI4Ti0FQJBP6eZ3xog+xb
EUyOggcZeD6GmvvmcQA0U+TSceZWz3bNw+Ci+biShV9kY9NIDbXqTfpBU/kHji7m
LYjduUGIVALJflthirEYAhgsPt1tzZ1qEjX8Xyzq7cuKOQ8MZPfiuK9whO8cQlhZ
tAgwTM8H0k3CWiuXwk5IES0imronaQImojGkLIRn3n+yrRLuJMHBMlnyDxNzSFTJ
eBVLWBo/AUGnBYrpNHWSHE+xY1+Cjh6zItPwcCuCSFp9xIhqDtM8JVBtwPdrf3AE
FrAFsPlMKKojaln0vFYDBKkR7BwzGA58oMgtxRbBKkjepZQPUNyLSuVN3rfB9OFG
qRBHoM1GtWmKVEhFvg2ArSRgI+cAXD3vzBq8oI4D+7WrVNMA47cuOO8kq7WqlpPJ
uRoKHna+xg3HFxt6dWoSAdHeRD+4VKnwC4EywO0/y6xT7lz6Zk8uTnhNVDSf4hMi
EkOoLCALytnfTl45a6n+KoIkmHKRfG3kiXIDryZtQRXhJp5VzQ7gJUo5kk3RYsW6
k0TGVFNYX3Au2N+Fz8l5JazkFpcNW89VUCxhIkGz64ADT8EfLqwYYMdlCY+MvaEb
bXgAfQl280h0+zQxFEyhdbYtpgVVSTxocxnB/rNdfbGAavWLx0ea8OnQOCkcF7Ly
Wnel9WmRe2+xFMwVyOCrcbyxId+SXW7zmaus0ycymO73ozAiSwP47cGZLzdb8ty5
L/plan/np9p/XZ5Ois9HcWgvnwa+gFKawNWrASfmTXWSTpoNiUDMZCzmjUxokmRr
CU63Jpaa0p8MV6hxlUXjCs7xhK4OLCMfBxdn/IWi+6mUmQcwsVA6dinFv2QvKDV0
RpvczqLap64UuIsUEL9BIkRwUkIpqN/edITBiUALVMU5deXzieZF/m02Yq49FuQ9
nF22L40BgXLLSINC05IqDmSSamBjY+InaxU3RsuF0U8ZNguGgtx0A59UbHAFT4ph
haklev4QWzeKbgrhYR2q/6jzjgRu+5bfZE3HtFlvF+pe2Z7X/CV8cB0Hgxb/hBuA
s5r4hOkMZ7/xFSroCfjqKCNpd5ngwz92rsynXcnAz4Oc8k+hgO9Tr4m8+ikP35a4
6bg9J6eT/LdkVmB4gyfxFybA3mM9gG7/nvR9XDgKnvcHxYC/+qCPU6/m8hMl2sHP
sdWsWrOOvjBl0gAdChgU3WUpS8KBv+OeVrkbOdpEA6t6eDzP//Da1zbKz7P2mayK
kpuXbUuH6WW2bx2zgshMrtvKmH65rUgLyt5EygMchnjxH0mCXQeRQRSUpcGiSYRz
nNN9LNo+xQfySzjY2cWrN1IBEZSfL6DUIFlogaCKcdZ2qOSxQEBVjDEE9GnpIbtV
nVc+qzHTE4Z+iwpNTNHSPYFgHk6ko7V/2oxCwh8EIz0AfO2WwkBE2ppQa78Qh/bc
PBVenaKRmB7jQomwUtkDINTYdKPi+5KtDL0ss6jAFg67G1+asG8dCdZqAU4oZ5s1
RWg4z0vunAkc6ebBFAwS61UJAZnWVKs29SVaDGvE5joiL9VUNcJcylDECkWThxnQ
7ITEKt9GvHu3ewLdvKs8BUOMQDHWUGzOJLFXYGGKW3i9i9gC9myvueaSShzD7Ord
CO6/MIDyAeQlW2WlIf20bmck3Op+6gkRHtD53kSoSfwTqvkP/7JCJ1qU2EfpsNmX
47EFC4vLiNgAKSd5Qzuvb/5aeShdAGcXWfkmCpEV1ny5NJcFo4M4ygu7Kkkt8laj
xpsyDR+HSd48ylsBWaPZeL7f+7eI9GVPq+AGgufNSrvMGxa/Z4icNE17yep7U9aI
hf6VQIfHeYgEt1Xx3EsRUZFIVqNTlmngTijMCdvbjGinudgG2/nqmXYPoeFbiKgo
p7cmC+HIdd2qvU6hUeYk/7BsaodIYXmGqx8KLy7I0NEriEKgmNVuSVxrA2HObOlw
yd1QcfQCnqsRifTIr3vs5jDgeAMvBGe4VD1bIJT4HaD8aPenr0ykCwuM0GA9AnwU
S2EWK0IClDks+52tSth6O7JBkl/X+jsU1zfMKW9Q5u4Xjeia6YWOy9lKt7mNfZte
3a9b1EO/vlbOCL9LexnEifewx00tCe9dDd6PJmzAOYa+jdYtrkXuRa61vS/2e8ZJ
OtEpZomxGbgaZh3s7k5H9vwdwGH3fDzoxgQTQaXqcdYNouGExnhmcKtwfA83uyjk
gQRjHN2KzW59VE21Upgtn7yDUDqz0BKtpOYOYPT107gbGAXeo2El2yoK2tVaFm94
NlazEPjNk9mKOOYKwKs6xYpCrc4RUCHqQrLHMG3ufoNaVQbbg8RXzFjXn0PARcMs
15UgYWzu9OsRZFSdToW8tRTv0MchetjnFaN+TCdpKtiez+YqtJ/pf2LBxFOi+WZp
w9v+kizmbLYF2bXVfNwiTDCEDyTxeNtd129gBZqgcecAwoUhOAJCSgr6nbDQJ82O
Wkkqj2ThlWPW4AVr6hPEEdHniDJOFGC6FThplS5aeW8ewazm9s0rm2LU23osOHh7
b1etk3lBRPgYxo84G02my4yDkO1tQaa5JnX8hJ0WqycqP3Z+g7nZmDhXXcT7/JnE
SU1z/JGDQUJxmmOZPC56Dun9HbdcbRjsAM2DdpfxxZnSlixc8NxemWFCXEAX8rVW
ZnO4mrZSyTcx80A7FjbUPm/PAzhmKHL/VPfEFZ32kIeUfochallKf6Jzm+25mCyF
pu1WF9twJMSyTSi5zpJiqBybpiTNaKNe48uZ7Z1nQ/OWdJrLa8O7FRHX6SWHDd9c
og/bcGlxKyFgylZdJud0HNEiKOX5Oy94GrZaAU9gMp83CYcgbcXe+nyjRZQOlI1l
RvqHrFQchz1q4shGbAi1a0RTdRaZGIZfon3OCvTDr9GIzZ8vzqYvkTBvOm8C/Fxf
fXHdqxlWum9r5ywo87+FCB2tnlAxJAmHjm2n3WNU2IqH7pNNEwGqxRHF2g9RVAR/
ZJPUdROWHG2TRd75xvbxgwQgrs63LRTsuNuh24UEYhoDuOSn7kaVZ843Ru8OY3FR
68rNw0GcBuDUqPH76VmDsxCZ7dhprovEHTNmcFPPnrC0TWOZTli6CTivO9Ix2FZL
l/Etj9pZm0tRDskhS/kqZUMIfrzWAqdDXpFFUJ3ErsjxR2bfnKgPCQ++FnNodAMn
imiNKsKrjaN1t4sZmnaPEWSjO6fELgLA5h8c+dnqZ3zfozT676xXOc45rOjJXoOB
7nA86pOOk5EwfFsphuZlqJbeFxQic/9SP7unm8VcUmFzocmDNBkGXkG94OHLp7cl
5mFFMEGOYj80Eu5Zedd6AMTnzBRSlNvSRg+od2mQs4MU8oGtvnSvYM/14EUe2AMh
rrUr0yT7qweAVMQofdSsrpHCdW/sd59DcmdcKS2dIidqz/V1oHioufFE5DvtCyau
6sDNaV2n6arx7wC/crf4zWjlw39wYAeiWun4DdhYliojSS8vl779DL6UVGPqf21W
hUzkiyqfmNWTxz1Wc/px4ghsdKILQRK1YP9wApNrxnqb7D2Dqj1CPrlzWhYu8ILk
Fjq98SrcRN/hGjLijYG5KLTUc0k06Zf8QmPAcAB2DH6g+x0BokewKlkdYsPL3GZ8
1CZE/BPsDaHb7Sj5uRNWTa3ZDozLIO2S2zSUjGNMr6u83WAPtxU0+vTtRXSP/lzY
MP6VQFerX/ULDnesyRD+NX+YGKzim4wZQqjmBNjEIgpIwNxm+Pyuk5J8JzEgDB0K
fVZSb++3QMFCUu8o6ogOoOGyZQDpe/3iyHfjJyC491i0s/ycIOimDv5VGaj6821v
tQ9N5B9nVFT3GCVYzzvKVvZnET/nMz2OvnWJrA5sApVjsLwqtHse9DWu6pzZFgr4
1Xq9xJSLYPbT8bNPBLLp6HxxSePUjMgjtLcopkOmqVWRKDvRo5sk55saY5AY1RzA
HhIAJuN/mWqDYc0jdHGk2VdT5vfDnatE3HCwJMWoNAJ+l9OZTsL8ZTycMRVgy4l1
KIDi2o0UqMuFHtigJZxLcpHmIqTo0pg6GK8aYbpSBC9t4lwp8eQXu0sniSkBUETL
5ej9UCcTU5e+DXNoX9DmkCkXXG5IgKEBtlN0vZWSQr+r3nXMA/p7UWdf9aD0S6tv
8VbVGbA4WxQeS8SHMYFugkeaaraETEOH25AQEIJ54EN4jdYPR68xjIojqH9XS7TC
Z0r38ckVrWmDVX7LRSA7gJVwmzPI1gpf6qIWv6zo+ZNPQd4HuutDBuwR7CYDa+lA
pB/izxX6kvdtP1orXQKvNYsXC8a4QPn9Yz5Qza7G7CeG1da/0HxZKcj6QEi1/PYS
VkMjIKZrYXNPO7weeykv4OxMeG98m2PG8Hi3bxayHBF+ImpFAXclpgGca8tT7opl
7nXDIWaP3TdcpLjlK7ETmwxsgjGB3tc9YVDA5iuO1Um3sPLm24cq2e/nSuWmXkCH
ZNaG35R93CLSpmJaD30Z4vl/tqkxQPvSmF63JTKLl+oQKlO4/3gQO9Ovv9DHJWVn
hyXQWFHJQDb9BRVQdvGDcAmW/mKQFacgtnvy7pfJ+rwSnfHPoWDh+zQSUz7tufiJ
PFOiBu7IdFf+qwJKy2VSC4WrwbTQb4fm7ODt4ZKLP+dGumKxhNH7KPQnkM70gVuC
n51Iyh2uCCgKL8bG1POAVVHlkjoXE/4RM2Ms/ofaH+WnT+DR+P3gyUM0kuMKnMBL
qqylr7B8/JaIkj7Ia6Z45BKPgTMoyX5zmHYSVKJvtDPDCPtvQuwDyBGw0xJTNU95
jS5REOZ3gzt+J8RTtHAZOKv+hpoM7e1e3Eabf3qgu7geKzWnMrigHT5B5myiH0BL
ZRa/WUYnPqi2XqnZZILjyADMYxEY3DEy1EXHqOZZOi5AWBZOhatNs5GCwBa+08zo
y3vv0Nr/Jc2yaTDvmqq3xRWBXhNenDrYpbX3pv3FvUQejviKc/cZEC1xFtADjk+v
EcmWsXxiW2dLCXfwY/mWS1dDInXbIhHWOn6k1qRQCPWdJU8A84+U9A/t1Ax4B6kS
UTD5Osxo1aew2Bph/OuGuDimoHAuoxEVMtaIqeWscOmcMQAF4wm+QMPIVqnoH9BL
AytBKk3idUzXWpxTdCxvtclysRl1a8RVy6nWizOM9h6p3UjX+HdqS8cI/sw2CxhX
rhjmQXTKp+40k/50F+ciafWjSLyNbq1yJ3NTQRo2BSc5GOVHUY/SX3uXhzE53Ndk
Zoe2ilbiHXnNfRo4xBwguwiMZjnn1IcY199NKjZcT9rafYNrgC0uGV3flnFA8/+y
yR+r9oL+bB985yX9aWZZjhhmj/XYz1TR5T+ptlTxQHXx8DWPycGgtwtsaqGX7c2W
ge8V+pGyDcCOm6dv6Ff9XRjgifmrsrnMOhHWD0FD2wsh9s4kRxW4pVDRkWQ2d6we
ClvfOjsMOp2gxzWCWcV5QKkaXuT8EP6BZsZdGuM0cTzyj09p+K8G4Vukl3VgUXDY
1tBl71IGZ8lX5ik8vTasLR64mnYDuWKQ3AlpUWO8YWj4Py66TIT0cD7KR0Aj5RXz
JBqi6ZdQQcuzEKMOLQt/5KsswhaMHCZAeslfKy2KUqfm0zn19iWpfFMpsc1U4BMd
GEK3d+EWz8NmHQWBFfr59DxbnQKcwNJySHYkMwk62PfRBxs8ZCwkEwuEwNJ+BlWA
wYEQZLw+XIIYps5CDSxUGXriaih3on9YNOBMSskjsMs5TiKGraUcQhegS3PBj1Sz
y3Uy8VbTUBGCmwsWUyHuJ3uP7eygB+SFDTaDIFB9+XgxZHyJJuRrqX6oms4erPww
nAvp5jiI42Bmx9/m51C21WXXAF9zfmiS1x3UeGRHnOEVIwhuX05Kkhh6nyr6y2Gp
1uWESxN9DwJ6kyTtd7cGWooBLVldwWIiyLZUZgcUbmJajHn6EFSmptiljH/Hm9+0
eZKur0hcxBYauHgpwYwlwtCp5qDjHNFIgH59HC7FyucKR3fv9SwWMr20nhl7TJ4q
kFnGBLvht81jMUVKWXA+pAxSm/Pq8vTSH0mi41Oi9MRc18NMPond2ryUXIx9D6k0
FVixASgY8aXeOBuGkzLBVpPhxTrcSFf4yzVrTaS9iNxQweNgoBcCgO5Uled4bvE4
lYPvzbUwXjIzHSuBrFlkHMkfBe+8cv0TtmMLL4jj8lkmGMsQKKmO6jNhaFt1xEfs
2hGglp1ekUjZeQQVbMml70Sj7WHz+ZNvXj4ffdwLBblteXMNfwQXFvh+XLwWn8ku
G8JB6PkiPYszDx7RzA28fbvDZDQEZhLq+5CWnLQPglo0NbdEbe+Kaw/uRYLl3lAm
wAd6u8iKvlw3Vk8Jas+fufJa05tMkqHOLqUias4R7ScaV/8HjLMp8arY21exS1Lu
mSaK9eAbtnZFgyNhzzphGvUdfAori+9aJzoXAr/9S/GsdOqIbrOJgUl6AiZR4ckq
8A/jItH0O2V4w9VxCxML7nD4/V0N+WChFeiiFSs4BznNGSN5Ro6GWukHoCyBSBd9
/pJPrmqvc+J0nXuNo5PUFfkHlTAgjCSRsMYuTeGYjGA8TENr34FYhn66oL9R+LjJ
XCProqTPvVUMZ90cOlOksmSUhMFq4hRr0I90rqgsdksWne8FuqsiRLJKOT737qsK
VWIRH2zsgFLtFX5MO/QR4iBYolprYsVO6m0ISLv1tnsmfsSfAv56aah4B/2QTy+N
P+TnQRMGn/FYvJ+/tOBDSMko3ncfVzpF3358Ps4O192rEGQJ2DHhj5G1Jykgz0+i
3SvKlw5/qEaOUF5Mojht3mXArK8MFe2osLm2DhaIFJ0Zn52cDk/N91Yp5LMQS9Cn
cLX8wcC0910bFLGLS5d/5vQPLySHbnFBalWVCyGeZsUaPQndjDMCJSxJKmfBer/G
n8cPxtJk6oK6yStspEm86UTmYG53bg8QUXhYqBe5FrXcvxSjyR21ZoFicY0ICvd5
CrU4F+MkcRv7k35aFOEZG4ECe5/ycoSUn26mQYdenU4QoURb4zif7kRSvu7McPAm
SykwgQOC1q8TEjYGyExUR/iZYh1Fb8YKJE53nNQmCkrhFheihxCL3JUDeWSRItSP
AdhCDVUujnz4arOXCNYnH/BvywCjDBoW2+QSiopX2lXpxK/rSpAtMyAiw/O/EyEt
PPPZpLbsSqN+O6osemksE3nEcZkRj3xuSg6teVqHg8IuQmUwU6arenvoQcBlMJEe
71hJ8q7ew5GyqnWhAwYLN3HCkINr1X2MEPuV9RxD9ciKjaIF/gCs4jsuLALaHLHv
/5mZJAw61bSBpLke9WMF3/2JK0TMLVebHtCu6enpK78AY0jy3YIOVF8sIFoPgsax
SUC2fnkIccgRzYbBJAeWTYppv5RCQ4OgElGsOxTDZOG0ij9EToH+UxKCi0azESIF
tjOjVqZWljDbC5PfcDyIPfPzQdBnSp8T8GshjxxiURGA31v0K1R0Cv8aR7JqOCRM
4WchtRIsIEQ64X4lVR3WQj2jtD+xWZiQT84g7WGfML46UhtvNM2rMbXiGgdM6iCc
9dTfGEybs6leDmsuyyb6Y0jOM2tYYQvHyPE/IUCQdx1qYJWSXtLx227rCc5HUQoc
hNKeOYy/G+YQxoq38OLiyI94t3YIN0vRpOOMwiubXrMR/LdAWshKVOLehKdip//K
nGO3DsOAA+UdIOX2dX/dn/KVv2JvvibBnn7wIa8Hq64AA4tbA5dcVXBO6Y+Tu1JZ
WsNm5vFpyQpQV9mn2XHUsf4eosdA0taPG3DD4ol5xec5IOA4eTrWoaF7v4lTvu55
DpsK/ygq+aARh6KWhK9qWI3BzvVje0au+brpYqjHovQGz3WKNYIpl+hTJ6YIGAYD
ML3wbkOOUYU1D0Foi+5ah2P0RQfFF4xqO8fC8AjPE94VOjcXZMwa3Rz12jhm7R56
TE+ee0qZlaGK402dszjtKgfseHegMWFVsgTFT3OpfqyPD0VnB88qMqYodzWsOyI8
NVHTOVzeSKsYOKXGbWKKXMsTxbOx6E9QFxPuEIH99OiF2N3QTpld3Go58Jcx4QYq
6LAGeZAj0ecVJkem6aLHyCshzThnNnDjMTNaSpPLusqPpSbpuRdeMVkGP7XrowJ+
eBm6T0Jt45jCr0q7Vf2SDshN2oaHZKcee4olZsf6EfsMGj3IYjIqGc0nVy5IIjnu
CVc90PwGZZ9SApJ2IkUVEIMC7iyQSpLNu38TwyFihtF9GoJNwW64nw7M9/49L9FD
UPj4PiprrQa3uelfCkb1NNyDhlJDZpdmPrKwu4cexwltSNuGsJPKSQX4hfWItjax
Wju4SBlDk8EmJsQQ0evkrFoqLolAvkfcPHbGXsowQ8dibuD2qk4rZPRCxp1cxSZe
iH9vPXFVro/P6sM4AWtY/2dqN3klISotGHvv318IKR3M4zHdgMM8NpL3FPbvI+Ex
5CBb4M1nHRYewNyuD3np3DBhOcfjyBpuridgC2+pCte5nyKPRJpLM+vvNPB1Em5G
ELKASDeRoHjj0z6lFM6K530nEI5PEPnlxh0OO9iXpSMQj1mhbu5oPLNZcE4vhTTw
9J/9hRw4Ip2U975GHaC8K657PtOgTm9Uw9i6iGnDzFSMsqHWViXtMuS7AlJz83uE
kGUPL3R/7SqsWxyK2g1RPgB3gpEsoZhSnHOZ38ydXoJLBjNm2Rtv68/T/bDYcWWH
49EwD7I2PC2ODk4MUShRnGjhgHOhslvWGJUr13mBCVeKKp7WKRzIzF+bboRs7evR
XFcZZF/3o1yoMBJArvuxBDid0GwLFbKOGpT1s4lROlC3nHoM1eK03nyhyBiB+AH/
L0/nOnVTxgFs573HUbTFvbqTOyNyKXCE4cEKR7kyU/J9owybq9VbkRTh5qyNOmHq
JJBiNTArA4Ga3anltA7J+tBZmBukHP7xu2nXsfs7GesHq2m39BCdgMVt173VrS6s
9cIkmmJv5jmzmGPquIkO86ocQRnliQyBoleW4JjvCwXN+9TiV9cTgMpjJKGmoiZi
XUhISG10Q4uWs7eeCXHOOUkgIax+VuHTqRgSS1Rsqd5ta6erUJ+AVBEB1WB7hXkr
XD8jsC2cB26wvl0O3F4bJJWejJIe4Oc6+38zi+8+YQ/jgma9IBpnYzizQqZFJv9E
KEoDbE2hR4bV/F1RBU4/mMagSXkejNhQYNxPgFL5X0k2cLKqpnmuCyi2MGdPoMy7
wP3bpApwHG4oWJfp+1xRJmra3qxhPlr/jUJfUujBpzKKHhuJkFpf5rKkhN+u7UFO
2Kg/M3b3Aj1r8TU0lKdzY9FjJcXRB8ey2TFV0yXNXK9fz/+W5O630h/pbIJRvvWg
yLQ7PlQQB3iEatYCWDogs8gZ6IO6RcM+0YzMuRiTAIlpgz5FPjXCuO9nGblJiXhf
N8K1deK/gA6qpB/tbjJKvWEE9ct+q5FQR17HczANAxIJbQDA4ztHDp5pS8WnkR/Y
2EX47s9j2t/9c301vCcf5pFD13tESewrRNoiOUl7af2DcHvk5PftizAxjoXbLtHU
F3IxChZ3liF2gxBVisnmoZt8kYcsDcpWzVK1A5fcGGmMEXpma+zLuPARuH2MQ0jS
KaNG5SNnlzWf2h8fg5gAZsx3ktc3U6QOERhUCuBSyPqrLGoH3Bfg337G1a8i6fLa
DYbhLvf0APcQZkssG6Y+25sHpfLCkIWIs6dpjDvXmKo8YoRgisTBxqjcjvGI68+l
Tq82LvowcTmRPrUSkahFTaK/oy55yUMdP6t++jmHtc1joIxcJaNFz+XRa8Vuf6M0
5WS0c3mQow5rkZOgTLgY27/VS9DhVPUS+xTom80u+LCFNSrZ3xFDST8XV7a7g50g
m7kscEnouPX+ocppWYTDftuwoNuO0VWisqYjTH48ojz71ubYQ1ojumPkOnhJF+4v
r4O0TXyBYwBNLzO6rKk8niVoTmJ8eBHCjg15HBR/3vUDuuJQgeRirjxu8Y4MdT8R
MqpTuxdG7AzXj79Xwe5JOZyg8pHBqxqBjJ3l0DxYWxwUbERdav3W/LRerFnhATEq
7d5F3vpCFg6TxUy9Iujm9dbJgqfVKlE35EFpf6fOH2H2QJeMSZ5vzfFN25qUMQ4A
+3wEYqZwmaR6oLt3qMR7TJ66Ah0x4fo/EVRscF2wYjbAwkNQ8lstH45eeAF4Fj+j
BZbvHiUgYyfgk+mMsJZoenJepFqPxS9BJmR9JsVtV3+H118pfshsEvWlJfAYZIY5
eZ7BjfJ5nhBNJQiq1Ck0H3qM8PKKPd7iNn9a0QzesBkJMdc8neEcvDgztOf65A0J
Y5Hor3GzSQBxfXKXD9gfIObnZM1eap8xo61qgcjhbfil4XHgd5z0Q+p6qlhveohx
ntq76mFRxLRHYsLlhicfr4XMCC8Hs7qFAmM1c3wZR2KOm/ZXEYNrwXmmZLjihK2p
ZLjmlDWBISEqkufly41zpGOeqoqsC74eeO0qpCOH5KsUcgrULv89yDiUIZYCPd8S
dbOn9a0ocJz2cYXm1opeqVv/74c3xtjFFh64RzGagPXLyipgONvQiNZrmGLoVRYZ
egM1het1DX2kD187IgmZOyHk+JGOdHiaBO7ohM6n9JCULSv6DRelIuGfEUzZQWOZ
atv9kBtB+3WZwmjMxTVq1ylyFiFnLGylVbT3+oh1pZizC6udSAkgZy/KY1ZFNXsg
Yjl5UxAyc7gX3MlQ5RXIwGSpQDvflG1psZuYD1TsR/PC2SbIeb3g7sCVntMyupsK
35geZyA9tf1b1yKQWfXrs9uHg/TvZz0cm3diKtEd0Pc2Ii+k0srA0m+PDUVh4EO+
lNy8ZOwyqJK5eaEc4sNnlnadZi0oiJn7ciPIQF/pbZOKlx1sDAoqI35ePNbf6EUU
20Su7IvYxCUkXhX/coVLzHkI/umQRn/ohHzjVOW2wTXoVXsRNE3GgJCvtaFXzlan
kXZyZutFkbias7+FosCMI9wmDAmcUh0/2IVwYLWE8vTXfpZ3N8OUFq4vOzpUQKyg
jL8v55QUpoJTKlS8ZRvXnN8GacwNRlM064dYqXMRjCBcbIewYZfhvyRbW2Ycz8PN
MHinGlXCTI1JKp2lisM4Yb/MUEYReW9kk+tIHJNZjj8hVC083iXXYB0bD/Fj5FTt
8A8k7TFl5SrHk02VO1q3sQccN71JtA+rV/WqsF4HlPTMHZG57JMPzuX05GzxCKL8
G4CbvJKmHMhKJQNPLAbxBCfvQbxkWHLvfVcFJhm0AWntgis8vSVJ6upPjOodcdAo
rMpSDRWaXIWMH3JcN/pXWOLrIVNKnaTFVN6dDa1JPreenxU8WlqsQzcHtpBHv6aa
eeiEwU/jjfD2Iv5w46EEl8Lx3zc/2b+24Ey/ByhP9F3se/zdbOu03b3YTOVSH/Sw
kMziuXo3BP+kFE1bd8AK11DMsPqrN5MIMiI6xW3mXfSNThJVknxWujVX8rtMqN3O
KQBHWpZDfgm8l8axSjAO4lrxn1/O5qZUWOhYahQ0rVtpjjcOeZAA4e/ty2tJ6DF8
uycT68v61oyi68gRvBmI5GgW1ijw3LQqJez0lNUva+2yhUYPd1Y3ge+tkihzZ2lW
QE5zDhotLB3pocU3aehbPv/UzODmfDTPkcN94VsJWrjq+j1U897Hu3PdgdXPv5w8
oqnrq0GjIAFs7h658vLfyij+RvgHzS6f+t357tn+oyl9MAe01TirggXARSpFJ44t
ddTvml5IJlAqVWO3WOMYYvXUR0LXNVb9OvcbKVTVshQaOPRXFS8r2FotAm4ORDwL
nIi2uAADJ61B56MEUEJy/6Tgqg78nxt1lmfrbwK3YaL6HjIRcH/UEuPcqHTTk0H9
SPDWeLiL621yWNjO/eSfNy8EiFK+sfAe3NdP/H0RBM6gqLG8Dni1ScAQ/y46jor2
rbtv7wO7cPOa5eS1K/nbzeZEpddM6pRJwuzXJIkPF5qHnVTCAjaVuz/ClM9HjbNP
DFMhOWEtOjjuqYlcSdynBynMbnNPoSwxiWZs72QZD6LaenC4iRj71ElaPS3MlrB0
qq1Pheczb0BeTzYw9RlgmPA20yz4iQlVdKcfFyF/b5IdhAwSDSTXOvugMKXqWW1e
y4oKmOLCVoY2QRfdA4rlAkBSw0eMdMTRBpmNWB+DeZv08VJKMakaZ51rNqPs+IHU
6GoEbpd7K0xE0sO43oAZxR9Q9XerqXMbTDHA++BFJvzy//RxnKAkU2gzadAFw097
63Iqs/kPAcqDCa16z/unhLl6c1vsB1kbe2EZsBRTNpycgqs9pOqimsYv9OSIlANv
8XeNOYl1nBe0+FAM28ifGppK628/Iv5z7VOSwgXTk6crFYvc8ZWuMU+sXNJluwGc
jrSPbgu4uM2pFBwsO4o+lmCbtTLQuROpYfoPrNZkdXZ9ra/LiKGiZvvl3uDG+DMK
a5qqtx9lZikMYNNdHk/Z92fXFCJOM7wVkNs9zCFkHW3EdPbaxRuQ5N+lU4/2Ordi
21n/FpZEhROqYxmnZdIDJhish/TiZWPznbrbA5+qnNshs0itkiPJpmsiZjtUZ9XS
7Cd6uvskXBqdyizAI4b/p+K2dThNVYsiZnV5RotSrKpNh1VUhRUlWgGzlnD5RhFq
Yb7BXhG9gCCCPu6lP+GQA3jfCMAPNosWcB85/ACU7hFXP5/GnAmimp+0xZqp9kYx
37iUR0H6WwZe1JrK8giPHvV02iYJiZOZZJsMX76dLUlNxd18ju0dGbD/x8XWKcJA
AF4AguaWmKVjRb8BFDJzQau/q0/rNM47JFe+0jORuSF0qQmL9j9StFjEZ1eZWiQa
5Q35v73FMhPTQzUkNRMnqYGbELGnMsN9f7uxIm292s26ZiSIjvpZEnT7ssNcjc85
uM2xZQjVa6srS8FZjF3aa4BW7dC6JRKQFMk2su9C3w66DzZp+bBBvFQ9O2xuwMsY
1pnOFDPT1c+OA47Iwz718TLzy8nr9P6NRnW8d678+Q8cf5SXvaOJBa/EFcEI6jiL
srnHrxYDPV64R/Qn0Ik/ZzA/DYFdoHBsEvlGktmJ1JF6CjEEVCnajKPvo2xaRnq/
NRNu5ekvmGoxRP1ZsayjihIiw7WueC6A4k1iKwAakJBlPzS1dPH/w5pxzrOh/ZES
KH7n/HewzFGSlU6melj92Wferen4wn1ltkaeIVyrliCc8hKdVLt0NAp1MBr6HwVK
ngvai62eDPJAnvf3N7j7xR0hYSdZOvMOUzw0svzSL8SUR8xNFrczWWTBhlIvPnia
s43QNWurKQxikxo03o+F0+uWu6lDiRTJDGJV3uQ13RU9zTrgWRsC5+ykqYXCcg5t
aqFp+kbP1wsGZMR0NskkET9gq49+SMO5wQ/PHik3uhHPeDEDno7+DG6Ogd2+o4eZ
n4v1pUkauKVvlY4Ncr0kv2WvohDSV4oN6vQmP5tvGXl733XkPDLO76NAD/Sq0Ekj
vuCWkaMQns92zknzAJrSzLIt9qOoILchDp1SE9Yn3zG7sP32fRZX6TlDF4qyNaBY
boGUgFoZx+o41nRBmB8PoBTQNGM7FIY6VG36QJ5CS/J3hdvIzxGNEUVvxJm7CvdX
hJ0vnRj9sDeat/BCSpk3dYZAKP3y6GxCekxqsSTE0aFWg/DRn4BpT7/dnj2aLd/x
62T67VMGz89QE53yMnkrN9bIPCxGi49pUPYK+xgyyka9JVtUcrmNNerA9O6OE8cR
yplmKnP4YSx4H8J/X//6jQNNVEz3UcbIg0TDLRRT60BCn6Qiirf7uDsbY0in04WO
rxRtGBEWMukTkFkIbJhkyAGp97VcYXdwskSkXjLT9f+OBcoCH6ls+24g4RZjquPp
XKONrImFgsp1cdjbdu7kqfRBwgb8qG7Rhla6nY1hQWm5QeIVKBP9Bez3iMu+Wyoh
thWQvt5Gr2U3h5VyKjZbDILD3khlBQNKWcCyO+fsNAd08RTahIa3oTvnhmNK+Qmz
UJ93qInqFlIitCFFV+5Zx/ZEG5QjvAt4WPjmfpvpgvqhX+2Eozjom2PySnYYH92B
+Rs/xIVtNbMgsPjkXG/gSgsD8eHDp+iFIw6s3mdR0Uk3S5hpzmSQO8YH5PvRFF4Q
9H8Fuh4t5P7O7/QimlqNV/vRp4lyvsbCkhpz4/YmpiV86x0W5zhzYWteYoZtzYuy
GsZCXWbrASs53c9it1ydV23hvICmoLZuQ92a0CPJKn4CWN1HoIh78ueH9+aT0BuM
JqYRmXctRJgeRA+x5Hxzca3pcG3kDkZYfKSM5MSRdDb+HlCPQW/0ovnVLVO/152I
FBkKfAlwaH5qen8aUVDNI6zaROc//nsLbzVPst1E/9n0Wtt5ewxtRpTF/XW088tW
hyeyLp6ZMAPvYUpepS9NoRWCH7PdQmtp4aN6dUqO0RqXN5rukb9F415cuyUD0iv0
vxFNvbhR4N+AnL/ueX3QSZmiy2FevdrpQM3UW8ECEpszaYpc4outNKJ60o2LArXn
L5+FLWp5sX5p52UuSafDpRrbE/grWpxzhFfmPiK6Z2ykQ5NXYlWlivtO5fl5deyg
rxWciQ4H2dl62cbE9gD9jnVbivI33ZX1Uz39TuH6ZIArkcDSvBmQhCkBuhBOwNeS
u8wUz2/kMeI3uQLj23trfnkgaNriweNj1/EMMHQeXAteQ3eI8wvWBqGaGMqvtGOZ
PYNrovQYXkveCSq601vmV+3soqxFowSeVD9Q8Ad6uAoCIPZDHJ1JiLIvF5gOGqQ9
o66hLvTdBicZXGm3aFF+grNEPNGE11ql1nha9mhJyemr0EnqQsTDpacnA3tBMa7h
lf1llJRaMcCz2PxJtFMDLkFtTz0NY3oexdh/nwK+10jjokfIn7xcsK1hV9tMSjng
fa+NmbFTIPm1ocC89c0OoMGgT3uiJ/y26k14fLjk6IVe7ghSFyGNjXmpVIFK3jT6
J018VeEJytWy6Dl9UGCyMFv7T4/rkVyT2tBs5MfdNPAaR9/lvA/jy/L4fFHCMN+t
Iewb5auXRw3QDhOyjQC69owCCd7cnecqdX4uIb3TchhHVmk8YlXU0mR0qm0+uOx1
9rkkir0u0bEYJDu+xvrdOBhJalV8X8j1fwQpo/DpKutGo5cxSGL4lRjjpaN26VB6
WpqGgDiRC4G6a+OsMsWmPKWkwc3ctUU6bcjSKMjrIt0FRm3Jzo+sfx+uWRx9Fawc
gAEbEoZlyKpwFbo+4x3m7u4rKGtjHvON1dVai+dlCwYnAzgVpmKh/bXXra4agch/
mp7biTVT+yK3jpzX+51EuYWwZSEM3PD5FOXHenITmhezqgo7SyEoP/IhyCT5zika
apuDicZXS4rkMT9E11ZxsUaQpMAu/N51G2x6uC0+5VayvSqziqj5c6NyTwuBJAFt
wrACryi94L3LtiVIpnmKXbKq38PXWRY0QHoHGsqF8K2hN32Qts7dLI7MhlKqQPQo
aLDBoLPNIGY00enK1s3K44InRtgF2+R9LxEGEb1Jcf+xubtS/CUoFb5kBXvHWUql
UDZGWC5h0vfxUG8rs4XNyyzrWIAiB0LdpkUUXJmF78YlsuVrkkbJ8HzKT4NhlOH7
MnKzDaCKeedyLQx7EFoU4InT80NCtST5SUyruZYYtUkihQBduDK4SZ0V8nNLV5nn
2XADrjS4sF8ARAWzJGDmDmrG556DadTmv68McrJh27nRV3Ef6LMy+TLrKdB5Bvnc
qhzoKlUwcfizso7bBka01KzjGd74XFeL892MJDzXfsvmr8GsANOJpUYaBVTduxh+
Nu3KUpW6VwxPNqpsORSpdm55Il1VpmOv9BXb89nq0CTFqlUnWoPbWeOxI8Uq0ntc
UQdb9rh4BsHACUrvMiKbTxJx2fCzeVg31VN6iaLpafj+reH1FpML8X9lAu2JEXiL
Kpd0+WV9QjaTuahsuEwOZqVcYZi+QlZ27hio4Ji1ICGHw10AEZx0ogS1Fl+2LCzS
karM8OiJh+8ojTfYx1HgTjc2wGgm61KuVwMJ5qd+wdt/Wl+XYbrZnARbeSBGkadB
qWYlHs0bhfTo3j2lqnkYlWyXj2jM/sqCVsbkQUNTyI45Kc7yE3H60x6bGqG96XhE
q6c3aFepqeSwMYQ2JWTjZmhnLWy/vt78fVY5eZG+dGZnXTofAfXfJ1YtnFY9XW0f
3+lo7Sd8DNPe72ckAjIVufCTDif2huWSOqapQZH1cITtdkSuy0QyVMGIezZspSOp
kqQNI66d5GFir6NL3bhR9Jn8DryLpNL+bvYAO+ZmckA7QBY0FJp4RrF+BKl4hQOy
Z8PX0RTPwhJBuZTa5ZKAvh/LDti21/NyWUO+b0zcMcBBBQNPTZObqP5II1ON2Zdp
uTwtvwEBuSexbIYW3S8d/KUW2vVioZGMuThexAY1bEeJkzsjW6c2c2tg7PFqVcDK
cB4r+udPvXZIkSokwhqXHlWC7QFao7jpyvhtPBCafS2dEKQcLhmu7Ge49C/mrg1B
bB+GlbnOrmqyND2ef8VKzlyHZvevWwO93huM4Q7m5fTsa+KXfqA3oBCRtTxKzpUh
t1EGhFVMvy8twwjHczqeK4FQhQnHsRSCQK+tp7Ot5/vLNErrvH2RNYWvtKtfFJBU
2HCEyGkTU6EeA5oa8g7qV1XBZ9iWAGW0bhKD8xNOJzZN+JeThqbl+2M0PUd4gkd1
/mvcZduHpcb2F8Vzwg1uHUVlTII9S2Tpn6Db/uWYAVSTnM88Klf2Umv+cMmY6jpM
NCDGQ48OVYtC+xIndXvSBCic/xgMiWpok8COYviM6d4dbhHTdVacWnxrfwGazVUY
MOYi7tigJ/5I4THXYIs/Ugomvyp8lonMSDZ+Gar+V7161zIMsRftkEG2gmg6cFfL
Ls4Dw1bQbCBFg4Kzt97kswa4QEQRzB0eRuhzvWUjoG6KO96hVM+uR/PHqm8qdCeq
tW+C//Q9c1+ohLKQ31VQxESbD8VaYoaqQI3iqme/ShgY9voB46KO6WivWwGbMy0u
34xKknJdyqJ9OdQvUjcbqTv+zMTCYPA8eiGc6peyUB8uJdBw6VyT5Uu/JPqpcqn6
S9NtmRsldqaXJncAdk9mugg8pTJ4QjySHvqL/MVLFr00YiHuqVeaND2xJQczYpjM
DiZ79MRo2fS3ANDFvYdlju76ImuVaXvBhHWJ4rpkmGOKkT7G62/IeVwZUDAqyFxD
SfGiAH4CG4qu16r+hhT8oYxb/vmcxcNU+NLJTswEc7iLL2ZxTtsoV3A82IqY1YJy
D1JGuCa2nZjNwCPdaMGTysLsxvQiko8O35DsxGQpTelF7jyfzPvnvt5P++hPweMY
agyfiYRs4bVXJlQslXeMJ5yw95O1QjHZJeMPBhf99VhlsmHA/NAcJUc6088iEUi5
L2KJkQbrihs1+wIPXSmADPdE6apZPB4cP5kViyWZADnLJzC9k5bwJ2bxKBbXELzz
8puLlIzsmswXnPZm4hJiQ7lO8cCpR7ONofL63RPoVo61o4H1/MAo8AL/AsWkaFH3
HGSR9CguXypnMGRbY9e7XJuFP93a1b0/9RUlKT5+kNZ13bsSef7tts3tDL7twm7r
oRD6fCtD6BemM+WioYNsBzaPa9wxqn1RFHF5I+C/cKavgxdTGDRLYTaPwRlveDWh
hr5kLlUzRXMX2ktWX4ztLpT8OxT7AslE6y5ME+Fmt+RU9ebb1ESeqTTbvrfCdybh
Ie2WXhhUxZfrLqJv4uS+DuPB0zFdggI+eJZ3gm/TCNL+m8+uKEOv7ojvGORZSKMY
8b1DMwxXX3fnOiuzU1TA54YaTgBItIYiAU4sITbxMyWj0v3InwxHfLl137fzzWPE
D8T33wms7OVZXmuKzGAwdHyTJpa/oVA58/3CSm0Wov2LQ5dKC3KotaYKmOmQn0WQ
MjQHzGRLtsFKq8bUalu+F7fo+WwhsOpdjJnRFHbCrLv0iG18xAEEOPflVWiMZKB0
E/WJesj0fedTiyzcLwvWIGlgdlEX9mjEnmxR09PBu/biBDW+Syeb76xqAP+ak0UL
fd/znHjDQw8xJNnZCjSVfg6hpf3sJVZFiMSc86fToEwzgNEH+1QkvtX2PWVksS7c
WHrbeoOmpfmpdsw1nbHfqEDKp7XFQwJJXrVnuKrN6A4UTwBf/5Zbv0eg2pQqp3ma
U1ltYG/7WGfQPM4Y19cSsVSbu7Oke0QoUReT+cBMhRIQppEMv1bjMnL9PETuc/Tq
lVlsFZYE2fdt642CJWv3bCDkpoPzh3uVVuwccjbhGbzUuZUIiDddiz7+4a8LTRmU
TYKJMwtFdcHOBGBS3CJzwItxph6Rn+Ccm5bVwUi9AslknJ69JcbvL/Kc7XQ2W0un
bApb65Z4WjlmeP3ZwS88R7aw/djMbWodiQd8gz1JoLLji50OQUmlNmMKthgqyqYK
i/oD2P9h2pFX0E2c25baXlsoMxyOpwHh8UqzTiYh1RYrOZwh+9E6K1A8CpkuOFgo
X3EnyP3KHP2848ChUAbYd4g35ijjGq93VcNKufYRVDmQg3dk8nlNQPkYLf3a+1LB
OaYAq4xEgUpc9jemsbgf2vxAc+kMQo7cO9/QxMmv2OdZtIzoUtV0UgthMy6MJXpc
9LU8w51NRz2NcTh2utBBxcEta1Fq7CNSzUu75n7nwHBGJtU61jsQNTm+svXPTtf1
IZTpKHsMRi5MO/GEyqZQ+X2E3STPzfh1KqWmcM0bLvWivBDHi0oZXohdaTByiA87
8h39GhhrPdQIEimO2Duhegquc/ETdUJ6O2Kzy2BMOxcsGpA0tSedO7/rM4Efe7Ym
06GXeTFppyHr/Ta9EZZ2AavFxigbH54SfOiHabDoqc3cc9zyO2UfddVGeK4EuE9h
FSbaktgfrON5Kjtp0fJD1oLITHkJ32XOc5Ca2jRFTcnuehAU9TEx4ao0TdJU17Dx
Ucv9pTpWWDMa3/M22j8yba/CCtQwkeQ7wWGyBqA4KPz+scDBrpbEsgY0GeGqNM/D
c6D2bdcdVj5fRQ19jk7ovyRBfiivYduWc1ngfRmLHYyAZ+biz5MaXAXJj52Go4/I
NY58qZjbfA7Uz2TcUAO5G5V43ZykTsEygqsORSipuvnc4kq6cyLsbR6YGgxjaCBY
ntDCqbkVYGQmN8QBpweU+M4jOR80KLrB4/HEToPdoip3r7S4ga9Pe6isiCR2xgmO
+G5qFDYZSWcA1D49GN2fAD9FZvtbOyaiwi2A4Xvcs5YUcfmTkAjnE5BRLQLMxlPt
WDvqdtVuBSDONyHHd8y/t5k82mcw1GKjybI/2g7Q/iBnyQH0UTTsl/qTMF+N2bJt
oYfqp++KJG+cvZkcixyvGgxcOZWaGB64uG6FmrXOUOJZAWpw9Y8cfAc7OZDSEW6W
HROUWaohe3NNHIqH0fyY8tnUAYymouS5CsJl6TWa1HKiQZ91bDmMBV4/BGivK3Nj
BubOeRIzLHSY3kNUP0hwcpjeN0OfCrt1K228lVQG1FhofyNg3FLl5+jswmsjia1Q
td4s/b+MmCgb/s09AqjpRE8Oo1M75ed3urn/+XHAwuWh6i9rvpCeJWj3Y3DR/bVM
4JM0K9wktvTnC8NFb4Qckzgo7ioApV2viqs70R/v+XF7V34SbJu9PUGDEMzL5uZn
vwjUUY0rmfiyVdq7oucIDATg5Y540BpoZdbi8FcjdqEmAOWGCG+6xnw2sEGDrdTv
A4jIrF9EK5GH+z6ItbJURjA48RhucW0nVGgWoXs0szks1M4aw9zrqxOW32Cur97m
DqgcTu9LINcLnIjczbJG21VSzO/VFFinN9aNect5QENcnEE9g4gR1UhqfifSQEFy
rS0mR/Vo94oc47RjuCTxaY0Otc0bJ3CiR+onmq+H9Q3P3aUf9Z0xeEoMoUOwAxGw
cjR5tb9LqaVbn/Ckh728MfX7e3Jd5mQ90kUEboxDPs5EAfTp/r3OTCPzJfCqfecJ
kVtcCFp8XAyc70iR8fQtdHIkiuzr1/M+3xPG4E066BaNJSfauJrJUymL1PlorS77
RQ5sKineIscxqJ0H0ZYIJt5Tupld43ZtYNaCdFTmCnGqhmYX8RWwBs68sXNMTRp+
9w7K+fqUN4NsWmHiA+ACNa1GiGojYPkGxl5X3WMIM/5wUcsJmBfpKhuHCZSLJRNA
YH1CO+OmEHwKrGxhaXhE3vD1+Xq3mP/Edw4ES+uhFNXg1ytNKb4gFCK6F8zQulPc
dDl1JtJpil211cVv5kOHC4U+M4H8Lfs1smzgX2siklzqrBtlNU4QxPWc/hhEbrtH
GbH5rOj2xkq6hmzcCXkTIamrwNep/W/hjtOKLMOytqJ9h0cWwZ8vR/2WkLnq4QJE
GoDd9c/6RyF0ZFE7KvfM/RHPH7CNLtXX1fQT2HpnibgWsGCNxV1+r2vslJtRZ1Ty
lUqsKPVCR9/K6+MYxyMOfg/IHq2991zDMe1rKAzVMF0cKCqBlEbqM7kxSbPWdVrl
yKfiqZBEmhDzQzEoDSULhOZGNzS/xqdI48prtDu93RLujSdEtgm2Uu912XtlmmLb
W3QRm6K2gAgR4qWWZSsdWHbOD/Xej3+s2KbITjnW4EkSEIyBnJVws5FUWDd10rEL
xapCcCjHLZjvg8YQWQVAiqd4zxA1MLDukmneGav1HuH4x/c/Fqj5AxCvSkljk4Ws
gxqRrQJdI9DgghgIpCgg+mC49fHL0s9mh6zs+Tzm5QewrGvLS0ITZtPnpbPN6O6Y
/bw4bqMQT9B2OmOlkG+W8lgmYeCZ50oxeSkYLqVfPiaihNdI5HMZuS4ZqBTiL8YW
KVSoPQIgEv1prqj855gkrSiSY0DSm4nAqB0scVI3SldvsYGbt3J7ds4g9cco4Mrp
EUcmSLPbEXYxS3M8QVppD+6HrDD8CS83HXm/5mV4W2QJihpRIpKhQoipHuUWr4uF
NEIATWtJcVai7BsRtVicY60P8NZ9Xl3Von1QP8HnLfYkI8XBNEWy0lpb2OYj3XKA
4iHRs9v+rkkP4uoSr1u/T8aUJqUxBYXdicWEGMaADwQ/Bq5n7sRT0iF4+fBKGPs1
714U+aOEL58yIYL/I1a7DSSu0jq/+4sn8rJFXfUmVklugT9NxjbtzFyiYGmv9Z2E
3NKqQ5++JISnDcLHukiaKohV/N0q3HBBAgj4ry9Z5cLIQoBrl/xTbu6YKylJcmct
MyjVxbP/go/65OPDnbsrHeCQKZuDWgeKid0hLlLNRGvkCl2iNSyxX4a2hbSkyR5i
RtZP1ZNh9t6UkBMRf/fK8X6uKiWcRNSZ+pTN66RMn3WarZcJpolkjVnz4DFitaK8
XQWf5Jrzt6QlESVs1AKdhRloQpKj3T+BFLgnoGiD+ctYZm3gVDz62+hgFKQw6xMY
H7iXBhCKTxK2PdA5Iu8oxRiP2K6Cg+PeLXuqpmkVK/ceDHEFlNOb271T7erYIRFW
uz3Ub18ezH1Uy3EBKAXgjejFyU1sqZHvJkUuPagjXbUrMJpe+nQe70TC+b4voXA5
tqJCckePSQS4fGv9JyA6HiL5kgUOBf/x/99YkqXuKwwQtZ+0ajeEKiImzoCdTZwz
Qyxg6YMaYICvfBMalPtM7gRMWVEiyRQ4B9CmeeNZ2IaH62BifIoEYC51a7pLol7S
l9g0Q5YQk/GZxFNyPdB8pqA9rRZkINQzGsVTZqL5otCsYhEon5WsaP0YS4P8sRRa
6t3EWQ/9wajxEleixmVf513ttBZixm8hO/giV3IQYaoaKR3THB/dUqVnhYGQVzUt
1pqCU0A3ZN80P+64GBtLSGz27rPBvmILpZwsOSvMf02bFIDSUsSBC6T8iu9HoJV5
NhoMjQ8VEha8g/KvjW1UeA+UBAEeCrq1XjPIte+wEXCdYsFQQgpa/umlOQSQiIVO
4JPqbo0kBYXf7GwH7tpSP9zjP3UJSG9aiOv9kcdsckXVsaMY7HUmQ1uMN+KG5Uib
3lfBRprFFO/23VjPcRDkW62J22b7N/1R0naiLsi8fRe8FEtpJ3TONsuBRSVXBLQj
wxwEwjFh4kX1p/F3OtSuuaND5gFN88egnhPih4TUkxKHtMfbPt9lFP8MiJsieQDp
8HsCOLL0KBDIYlupZkiIkk+zNc97vDq961frDCgqakRzYwxGjnxQA407/1mUyYxg
QO5WOBMkdheZx6S3NWlpnDeB7yS0rBZ5NPYAWXP2irZ5zBle1USK55V+TZbc6Qbp
pZ38iU3uLJ44k3wdKVML2loZWJftbgH3G7QWCuwMYIJV4fB72EUsLjLyyFEdCFWx
0BIDQtBh7/M87r25nlRPYL0JaU/dGh6pNJ1wBkELm+jNspUA6ZrGjOrcxhOsXYBa
tNTmguRnq5apSuagrCrZ+HtqlcTMx44OwzjxlddRtBeuuim0qDicH/iA+jbtUDY0
pn5g8lGxAgh+rxPzqkariipZ9EdQeXs1b/HlWg/RU8pLRjpPPvbGMCd0YD8nkDlQ
BhsSwjtWG0DZgG/7/o24iTdr1Gg/XFm39GZ1EWSDg6NHxYC5rFJ8qDi7Qs2kxmwU
4veBciJ0Pm2jy63fSSxj7tV/ubM/yBCTfd4VqqmS/xJRgr2ZhUaxnlCa8zYQreUV
AW0FWOYBZsBIxQErajWRwEFmwUgspXfqSX8C90eY3sByGkmGSWiLoeN6I8fxJcgj
yux6MZpFu84yPgyjt5pIm65anvTQV17WIMIngktITpfYrjd1t3sayPWZ86cyaDb4
OoGzMDEDYbxKdpak42wOOjr57F1DXIA0/xaBc1WR+dMyieU7lZvVAnbgw9MraOpy
FVWsYdSiz1wi9ro6gJFbn8SeyFcL5cn62m6YKapquYZU2dABq5i9cL75D/1qiyPE
FGYc7XQVK7nmF5XNY59wuAwVRzStrGm198eKrvyQA37Ef/89rqgK8ACgxvn1ApAT
E+nEfItDNHNwnkSqsJaUf+FGuG6yya8b0E2gp3lGfvW9Gq6gGgq38apBQnXjkT+S
johyWCc3zaRdctwLA6WjUunCfKbJzMaD3HVWbu3ZbvvSGymj02XBGHhnb7UsEcrR
SO/ivcsrdMUnbWoChhWaVuj1b8rgQuf1N8R8cq9yFa3S4S6DK5Ssnk2FoJTcP7pL
Uww3RG0I3XFLNV91pB2zajpB4SJARqJntfB+gHvKITLHOC0+meKhMLT1pLVbvU+s
B3yKnbD2iyDq6NY5orb6R9DtOULv5eB8xTrdpB0tOzo7LTmGQpMGUmeU+R5+Ftuh
3s/lWL4cpU8mUDr+5lR30jL8vP0uuLJLTjG0zCyTA6SHRbkHZOY8YYvNT/7PY7JX
voDnoEWjc09HNIT9yYCvyVfaHEA6XWZ7uPVOinaB/UmBAOSFU/GqnGRLi8JnX2az
jWp2J0GioJkv6A/HO4oJGqmQ2YzbLPavfEmS5B+fPLwSLVezwBARp+OuiJsD1GYh
vSdkZV1EBXY3o0Txzo9zSe9AIvFd8Ya3tG6r3wwyzygiKhQrCmWMD9KCcHbz12Mr
3+wo3QIk0Pw9YhGywmwYXsE6ZWPyKI4/ikKaUioPdS8epC6xdQzXZ6iWmNu3v7gR
zIZRtmFRaH2U5fGEWTtIgrQ29VxBrsamIgGkmA8WmMYkLKRpkZqEjWFuOaxun/yL
aUV3eICIkDVE1ZpAuqaWUikaq7EncAV3jKAbNgrqN4fYX6K7L1wGeyUkVYqSRknR
sg99TA+axvlhw/M/vLV67dEc41YFSTJvWrRtHBgryxhfglpyXj4WroZS7BHvgFMU
7IEOyl/ltymVaUAawvZTdkttwrYAfGxWH7PAmEBncP3RDzOv2y7G4i9fthq1SZn9
MgoKlKI8k2Wr12CWPMKPjy0O1x2wWZW684mK2KD5WfDv6RvO0YV+KOb5L+jFSUbU
zPG7rGkn1jhUcOWSFGS+Rii1MZV7Glz7U7ckj563pEpsQ5bvFk5OT2DQUpuwU3m9
pUXL3rCyT7O0tj4L/tkMCn/XWdTEcjRqFH1yQGxDqwCcDzW761HD02gig+63OgHf
Z0mBhvd97YE1fQ1p9yCy2HwbejxG+YrIIWYl8nB9f9Q4tnBpUhCQg+7prXujjsES
PH6KnAV78LCAiANkU6Nc5SqdZSPEc9ydoilgOMacXrZJx/6jy6wVVjv+8M3i3YFy
Ho9VmV/4pWAAKFdf2CZGAtpnTNJbVQOSvOkLkBXqnu+JgYaVKvdbHY6uGjEGLCvQ
mONWiIuG2gk4yax4Auvx5jFFTbyBGpPiCqOlLQoR/umpCvBPOKzP+Kv5Et60ozOK
lo7oVnm3wUXculGFgNeffrpSx3tkTMpdBZ+mjMVpmXn5yJS2AVAJDfjQnRsEHk8T
ehF+Tqyfb9RUtoq9gIcFkzI2ZZc/dXrJwHr+JTTDnfLkUqq5ue6ejNfOfq9jsryt
c2YtPqQu+oZY1XLGy81WECj8iVGO/HxbHZqApRtgd4bEiIG51M5u5RvA8o5nO52R
OWFKZcoX0iCUHQxGXLE/vzoCSDFrZ92kZKID2EZ/IhDgTTgNLd6pymsOY0Vml6we
Qdob5CbAr92hXfOxDyppy6PoX+vxOcsstHgHzhvZm4G3R97T3KezxPANOKRMAU7p
7ZMVAwHHYg4NFvPOp5y3fdvkkd7Vq7XYq6f+RmKa4qxHu3RYn72s+adwqPaPR/Ug
mgJ2gkNzoY3NrAUrd4NVWrTG91qwmFe3octEqX1zOeIsm0F748YGa2w3yYGI+YsG
eK/52Q1gl/729zYEVEENWJFt3UmmV6KqKd5+w0mO7g5+q/EydljsusvQSJosv+vK
BvZp/WUkKI80n9RsCnA9EO0/1C01oXMaA9tn17mwIJqcEqmv7DkCXtzNlBODRWaF
WsSInUAtLNQOX9JIuCDkOBEFWQO2uKOuF9iQ1wI6I1IhFx+do3PSqAhAAqSwRuZX
dAjUrRwr9YTF1VlCPkxAC5JfQmzrDEJAinIwGZt6TMP1Uin9H8U5mWFJDjlhIfR2
1/Jxw8Kd36NxbMRDNkbJnjXT0O64ThwLNNDdd/CPi3BBVYfOx0S40ljBqNvfC3fA
U5HwQ1LC0cQAzR5t0O/GUEuP1mTR/eM7Qb4A/gsgNuio8fepeFYDWrpQDek52z4N
x7SE2WbE66lrvao3H3pEd8pkhBLF9gjBpGbUYtaUVIHxAelmEw7wZT7KE2wr/MgZ
eXhafUuluWHK19WZeNnPmpe8STDalTQAPLbJ0l/YIqk2/u0oIRqbHi2Vc2nO5FD4
A+mCd4Hmy2A2cROh/ov9jyJ03WqwdXHJsLwXg5QMlvouHw4Naegq9qfNIQ1ObI+O
+jYs3nj9poyz/gUGttkCGQqyRXdIafr1TxnWz3MEo6VA7UX/7CpzARrGWYaVS7KT
7k/F+ltzrmfnYo16GCmLWPtp7paxNo5zhusguRuSnrtiAoqhh+b8nVVTBYyT/m6O
YeaaVj51BRPB7iQ85eG3vGeoVAdarsu/dmCJl/WmOvFSs3RLnH9ynbXqencJuLWL
f78NQI3O/FDdiB0Q2Jf3gULiF8QfVIX+dBPvrOI59mgOdbuU9xCQQkV4tx7wjjuu
yOQPMRdhii78juJFYtio93Jzr0lLCGNF7izgnthaNk6KYN4C3hbqF6ejh0HZMdkA
gKAbe7rhZAgMGtCWlwAQXIBNWk+YXycFB1yN2hDXiDWCCDgTuz/fdlCi8Vfp3MlD
FNWE6+JJBlZVEWvWLrNqn/ByngnO8LeArc6pxG/jWtne5jYdPDBoA6BPQmTTsOjx
uSasZiYqGjeS62O6XQnCCmwj4ultKTPg8BasCOj0NYnp4iDjxTgVcchfa5EaBLZP
jsUoMHZoh0Py2sz1mkvbanwuLdeCU0MyxVr9KDfaVyt41P/NmC03qYs/bpyi7F37
iaP0U8drl8A1SB6X4vWHDs3MkplytdKIrMw2ZJeymdxHeYQ/buX2u8dXQnTQTDf1
HSF3W5CdIp5usLUu5dSruNrmzZcFF3MLi5fQg6AlzNc+xpBujFWY3jePAWWy3zPv
DZqjLJoPRhhMr+fagyNddeMWEVwQC3fZrxPnHtRnBw0usSFcqapS3JEap/52K1ZW
JKr+EHDbUPmcYHIcoojCGrS9bm/+qK6QQ2FmuHf0C1Kf1OMPISyvGbfF6zBUXPwn
Tlz3H9KDL/47teT1tEsLPIc7ytEscopnEGx1WW3h1ldjt/6yEDT54u5n+YYUJzp1
LeMZASLDQ4ak7Z3ri7zYeXDS5DLc7s3bfvBBMc0np4XfYesa7coZpdhmNH4bJ1fD
p0OHz0hAM5vi2eY67sKpRRMM6t83g4tS9hqN7UprEo36g4W9OCi4Sp6+SaVtiXBp
G0kRbSwkecFcQViCzlccr+yG9Qd2eHc1wfnktjQhKm66HAbmij1j2Li64YOpkVOc
MU4b5N+RnFWw1X0wPWvlh+CksrIPQ00IGFrK8OXhanHAmR54mAboE0rCfs2Uj82n
LxQWigmrioQcr0hqJTGp0yvZFH33BeKkIMH5QG0tsz53CbS7zAl0Ow4byI15vNFH
kv3idOBUlkCaJjN5QL8lpNHssTPZJh2l5zpmI3rq0dnwdtNuv6LWlIutRxWwJ3/x
4zWRNKvLIEl++8bBKIcLIUOkNfoJNFwFnkKOYAz2SQp07O9kJNELYSBqvKoQQLjm
luMhVjx2uN+iwr4glOagFg3GP6HOQNSWmRS+Om+jKfYboFbU6NjmfAQL9tUDIK0L
UJNimldpWHigzTJLcyz70rFHTYdWYycH1OGuSqUSdkmhP5j33rt9jF+nzv3j7Jyk
f7k6mDq5a+aoVC9co+VHUmhzIK+gmq1rEeOqxV3iOIm0yxfpOB/mznm4N3+AIUMo
nB3dZ4PR4cnkQ4JEytfl41YOP/jAQbPTggpnn+ItZzwyxwsx+3KvUa6b45vb8HyY
ZvOQuTej+7nAJrXFLabW8u9W+ut3PovZ0Stx7Nc3kjVHTcFskHShIE2QPudi3Frg
2YweKEb66DCiY6A40OxV1t4NNQe04WbdnD/Xl7RhIzqkNslI860dfRIGvtEhWnsN
5DhTdAbZn9IGgknq9NkXd4pZIgiwPWuj8rdpXt4cFvMUcjrynLrYecboyY6WruYX
yRojgH9tN1jo+dhH9oXOoVvnLj7Y5VzVkpSgwvbFzgawA+NZE9L2+amOQgJ9QFZB
vK1T24vyu0W6XUCiipM6xApNLL7V0njnAVfL10njuWHPZuPFppwoVy18T2+hTi97
lGjkl/+3yjGMeGS1THGEwO8XFgUjgvNy8kvWbW+lAx/4SE1yaS71jC/FySg5H8Cx
X9cvCTJgZv1Q2jQXTllZCTYBP2+CImUqcwodt8a1OK2CtS51nZPrFskJKK8TMw0L
qE06wXqAgPnv4gKVeiDJEjk9MnjyXI/HaPqF+qz6pxmfo9eHuPpUVG3rfy+H+LgD
U7FsSdVC8CfsMCwzl44GxV/9lj5aYiLggCjgEOczxweqAU4RM9N+aI9qwXv/vOyS
USYdnFTexTwpR5t35fRJj+QpTTWkcl/s+tixP1hWvkJ6IpkFh0PktmXB7P//Ce5+
Rd1jmaZEp17p2PeG0fM9pku5gOY2t9g0F2v9np6veuyjCPsSVUixETTVPmQ7/ej8
OQF0p7q1MThM4R57XDI+dYs8LrIYMQGuXZ/sL8Cp+r81UaxFU2SMrbDIei0i7bbs
Xnj1hBSVFBa8q9nJWTTIW1HssiQF/I3AIUnDFT+JiSVY1UqR65Qj+/rkmwwLbSAE
R1WFX0vL1GMDR+jCtCHFW0IMBkvTTMaastlYh9s31BoG1WwoPwfZuPCZSdBT751E
r+F4SsbfPBbsPK0FFG0oyIkqBEZwjipw3hBhcuzdeJdD8sDY7+U6XkeErqvk72nu
FbT37/pIS4KTx19+Agj+1/dvnNapfqIBlPhsrHtejOg1NMkgV1YDqRitCs/CFf/c
HMZD0m75XBKi5abREzm2fWIIgtCMiZw8Y5azpRqD5zRPvCpDYUJei24jXVVPwlHW
c6ODV91cUXw5is6dddO+t99YIjhXSrNKB+92Y4YNLhmLiOs6Orb7zr9Ade1/p7q4
DutLUEuBXNaZW9FqIug7lebiMW7QhNGoyJ9sPEgNbpzKOgYLg6ZQJZ1yPT3v9PJN
vzxQjut3VP8Mtwmrd0b1IvSSYS/T1tvFAoZ4Qv/hrl/mJk56YS73njY0iENCPQAO
hAfyOS6t/M5Tcifq9khSBcBPCW3jHPIJKB7rIUprLoSVph0QsOwgjpd7waj260En
iD3WSgREIsxkJ8+BzKihIiGwGEsmve0dlXp+m21/Gkb7sCAdrRmGAHtJo07VrH4S
Vrtno+S85IzTk7skSHdiLPRMWhTOMuhtisFMLyVLsR7XOuV0tUeZ3VdyEE4xPvVf
0Bwuu53d8bvTBxtnDt9XIIy2fdCkjjFIxq/HZlRqR0oWKpGtu6uevNGvjNmgHt7d
pRWBkLOgvADFZ4QiV1bizMlZJ+iUjCjo3SMP3HqewuaCPC64lao9+37q4OPGpKs+
2qOdEX/1+W4dFrYxQOLZEp8b7crIs6xaBVvGeHHc2uxRLkqKT7apRmupDnf3JEQT
XBzbp8f3cNTW7d9CGXcKgtigYH6ouvDKrhib6U+iyQgIyrU/alHJg48hDWHT0rQU
q2sebp3utskLekn+fmC4i4csvA2xDCtmep062CVJ6MkGl8NCzIPKQgZkn/2fRMoE
gqLE7f8xpJYWrspQDm7/gzTDKkRV3xBvEA5Lr8MoxBO+NVNovv5do1PBWRquK7IC
daIqQsm22Thve5bODLS12QJhzKg4ak2JPEk5Wr6tIift0hqB6XZOhNwBseNpk+OH
/EkMjjJkU6LrLjgvscldp8bCjZizpaPbLUpgVmPLaEwfzr0FXwAkW2bWJEqxXM+A
mh+HXRcfXJv+KxtYumdHDKVgaf1GbPr2/S05Yrn0su5zLen8z76LuHUcAkcUmApO
FVU/y8cjf84fMlZ0TGTpXQGNVnlDhN1izOaEucw/psIiDfo+M/iv338P6l5eRfoV
GMxwTqBbYbl25bDnKmQMvGBBcAYTLU94WNc/GGlK9NTNxrHzPEwRqIqgKjmlgg6D
kvqOD7EtTYu1swx02TXFGrtmOaB+KkkuIQBv9PQUkdEXJihP0STze97QqaYXSLpJ
oHnY9SA+/RdDsoSyjGIUagudE64LAea3GekH5VlMhE/6nwYomZIC240htDJIlrHw
4ExgWjEqTMNtPXimlw5i7O02Lm7MYB5xsxTgQvRJ+FcMDDKiurSH76Iuy8kB/fpD
q0N+lqO3yblX3DJR0V7s8Wz1W93kmivz6aotfSiQKALLhaP6lTt4msPV/VT/BBMZ
1iPhmmKTNQXYgYVxqbsEII6nQLB7KzAwFHfve09+dRHQE9tRejnzetBcU/wqngzb
veZjPyS8ZUtjHl68ljtccovomsCvjp3CIvL5n6bHPyO9zz7TtKtC0LeqtLvqgx4+
1+DxSBKAYDNkANtgtQ2oPDYDkaH1S3MmU444CTjpAa7sUKDMh711oPVIBmR7avYK
GQaWiVHro4yQVI9/+8PFV+hYhCU8/iFvSbCZuaeFxINIOi+Cu9jrrTKB8UI2OudH
HObFI/0JiJx0MXxXMyNSyDCgSOLXXOdL9kp9+U1gletPg7akcN6oXjIqQ86YsjQl
1OtfprQLatmjMnGwsH6i0r6IK0V3YgamZpBllxo2R9MobCBcZSwoliRBR+ufxZui
W6AmwtWf2ag+4flTqJuNypT1IIvqMmIMFG+315pAYdVbDMtZtlA3/G2LP8prgY+r
Qus+pDLGVcjEcT40jgpF6ofUDutglp+K4U6outVlI+y5BEBm+ye469QV8G2ve6Uj
zNkxOApuAmx4ry6ROULI61l6Ga3Dc82HY5gJbOg5DFvrN0Ifdw7PmPVoNpBkqaGE
sYobALJiiREFc4Vv2Y37/D0L4Z//LCvupdZv5ITruwATaC7tkS+x3Gm4WNuKokqu
SpQn37ezSA/Etst1BD+4wdha1ycKgH5KY1GtHtO89PFFxbykLaJbSqZ4Oo/WNllA
W40xWgOtnARW+sLoIbt8RR3eCi/Ob2D+NcjDiRNOuf/2gfyt9FlZSN8hn6zFSCmM
INxNmIes+3mWYsbIbX5UMCyx7XXTqsqjJmQ4H4m2N1YunLuq/ialIsbAu4bTOnAB
NF9B6V+67KkGIHf6VN/Oyp+TMwPinCqoHs+yhWTPmNCnbKQGfs9JGs8hw1IBS5Kv
5Jv8f1CbeG1lUotAjUfix8ObNt6yq03AYy1BbZ5C4M6gS8YXKYI3+2axAvi112Gi
90JzQ9XCPmsndP0pAhWT/AcTJB5qyuSNIs6Un6SeegeohOvBgIxxvtQlzPMABHmO
cpBSQV4ckPi/gpvpVLqEoNMozgxdqjDeSc11eFV+6wj0xNQ6Z6hiQ8eb9AISnB7v
x03tm2Q5Q4U9m04K0ItlSfB/5ckmWzpHbR/YHpTgLkvceb1YLfKGTMTgVQAeLY/d
dFUe1vgG6DtbN2yB732nlBctP+dlO3+ML+YdkTbmid9q1OEuMC/fh5fWksW17Y66
7GGUutMYPhbDavy3KIvz+r9PQKb2Gk1+XPQUFm/58pAXo7yipP6GltS8VOVyrg9A
iBPNQboXtqslT8abVvix+uGroqdUrxeW10REq1KGejYjPRsbLz12yInNkr71ObgS
JqGRwrmNNcJ3O+nWYYza6aDqU7xTnzzgaouNYPoM8u5MUHud3a4kOUyH6jGdfwJj
mLk3vLNXbqSM+IHmbLEIl/aat1Wfjp+mZ4Yn1j/FSJhSJOHhIzCRz3Fq2a2zRpyb
0IF2Hw4HEjLBGXkTYKwlnyDtSei/tfZjxJ8WIhBAuwKyIW/B68U74zLFSukJcJk6
sbguI88KTZrGsJ3R+ExWxHSLidXH4yxhh3JXzZF2NiVYpModER8kUg+71Sl5SZ+9
YtbwbPH3q8ffZiQTkqN05exHAWDyNGMYSST5x9gEvQcuukt2p5XUk+b7WfRY5vh9
sIOzfBqYiRoIjy8cM3j22KubtsQ8PeJ/XNb5gz1XG78uhKz0Cz9IRx29qHZQL87I
uBwNeXaPvuiinjBY28t1Wqqq2GmrVcex7rqgRhOJZtUdshzkKb629SuF8ZJ5KJFr
JKL2k08xLWILIh5WVkVGys0LdeR/HnpdL0PsZHJ8ktr9zAX9UjDsZdf2p4Cw6oow
J1JCkLxzYF/ekk+u8MonYutTonxuXuOIfWeDYaCS5UKjryygX3gysSE3KrSiDAbW
UL9c4XdOWMwmP2bBcv7nN/ticHaTKzWEgwB2R1kacPGmSaVEytE/zDZcg4Zy5to5
Nom4/AGTZeBNXoiDsu2x77gZzCfjrdyjjZVTF/MflfxF+ybIhTrF2lb3EoYJfAdU
KuVSyUIol9YKWy8R5r7Gro1QxdsByfI2xBqjV7LEYn15LMlFB8kUgsJiokmZvG4S
lgOsMTAWp29IdOEE1bXayKKtlFlxJRwvqtyOJN8Zm0LhWGS5KJYCGdxO+4cAHwY1
A3Ny+i0d0E0MS9tu8fHB3zbcLdxsohbxRQ50EunocClrYtsxNPFTa8RrLEvZPEPR
cEfdQu8+uupUKF5/8eqRpuWQC9PUwjDpMsDtOIW2OJJAZn6bnIRW/4vE2lbObQyC
xgUAGWyimYypzGwn/e1/KxgkcCiz/wIsl+kBCZSvvsplyQRDv+mM5Y7loZcdr+iO
WUWKSUN+w86VhyGkb1CAq3uffoE7FAPyfyaopBcgWWmGJlX8j9uEoPDVVQgdBpFq
FnmfEefQNvLNuKqGM9J9Ozn8XJxvvld0QrGQoIZc6EVZ4LCVXP78KY3ZHwOd/wz6
F/+L7lC7UaDR+KS/59BHaDb6aQwU81qBI6OElEsdeAb/6g8sHEyoshhXTLH4L3G+
f+hDQ+VuLGZLb8FK54xu8Aotxb59YCD1lmje4/HvrcDvaAuzDzyquLcaHvglsi25
+Fd4bFvGdDmK1htRULkndnm640Quc0kVWnxWnCBCObNoyrmx9lvamFnWuRjp/s73
0jRsfuOlGbJ+9+SPI420FEgUXIOrhvjg+IQIP2pRSV1VQrtlQVmO0kMTMn3K0dcU
oMc3p5YczA95evnnjRy8KoVuCwlAdOyae62/8eZEElJRn81XyxXM/2YjbnkXF5ll
7GShl3dYd1Nh2SODCBTa0QCKm3Ax7okC1EjV5MqCvQ+wD6Dm8xQpNd0bhIvopM8v
oPKK0J+iuS3y1foH8qpyrF4vRYs1VhGLGQVjPFdr8yPZhJl+DL3MDZPIvZqIDP0F
6LdQd5cAZHfKJD0VMHFZTx5XJxY2BNVdotduGnD34JailEMPYWzbG3vnmlbvJQzq
8c/71f5qTw+gWf/3KZ8TcehOm09jtSS3R5F1xas7AUFxw42uRWLIUEqe3MGS2PiN
dZpYBGfRHhGgqf3Xqsrgk0i6BINgcUaMTNNcvHcgRalT92TFxKr5Q6zM3XI4a11s
QZFT1+N5Io58e8vS8tzKuyDwRe4gibjU6eHWh/3WfwDDVHASpzy445uD6AOGVwXo
w5FafFWkEZoW0xLnAubOySLnToepxepUrup1ljC9mgAIouWznQ84E0EGFae/+/Du
W74kuIpsgxi8EIVG/jAcMCHjXkfmUpKBpwlvH4qyLkDXP7zSzB73g+wdHv3+voWh
Fr+SucXYCtVoRAf6VDwKaeIKjv9ejyCONzhwARvp66bLMJ9FKUZNXUJTtfKbP5wq
BIUmSrly4vJpnjxhebGJTraBb5gxrIS2dQNGt9ZQ7DLq3AAURFfAMcYpOJb2LNGH
K02+2JQZfBfGLzmtXRAS++bokHnrOpWf6u1LBWAtOM2+sWtn0bqZgOphoYOIhWlO
SC46NigiVrhxrpIhMAIb8HoSMUaQ4/lXGqC7Xf4xRTWJf73vMTqRNxe2iGFz3mrv
xMMlC43u1VROSgIJoQ8hs0V9ic6caWfpl9WWwImChmDD1WaDB6rXcXQO0hrXam6z
j33uOkzCZ8ZmDZPCuMR99wiiqI5pkkcMuT9chnvJUI9QRqYJhdYwexcSp639Zwdw
vEng1rPOteaLchR0a1bE8NUPl8I4ILWTnrLO/B54FWZm/6yewTPDVZz+r7X32rZZ
DjkeZwzjWnz/tMBAOIkJypnGbmP6boXC4CmqKG2xXPrke5ZcKq8nyR7uPYIFaTRj
GpKA+6/IQ99R2JJEFOIVO8R2Rcbk/MLIJolM0UPd/qyIrtv6UA0SIWuicNeHUcEQ
nJY8+niT0vNWrLX5HDHrI+4wyUnvLnZ1SuyAj9tfLdme1CyrQCbA+i29Y8kxB2JW
A44vdQhE1cCzD35C0DwlUnSAPT4mD+YWkDdBPNYvTRaS4fyF6D/RVCoLdp9bcktg
zndHHH3acwR3yaLMZA4//wbxr99DfkxxORt4byS+3uDfAFQWh8e+/29m9VM6TZ59
ZEGo2T1J9SQWOK0rp9Bq58DyUWax1J+EBhCdJCjxugy+oVlsN9HhgOD1CZWizmGv
Mk4nB8hA5hPA0Vq4RtKeUP49c+QeHv8qmwHDSAI13q+1TY4mpQcseAE10GxPI/kC
awAOsBGVcGzbHnwDureH35sKhu6bqEZ7s98CVyVL8di2LAton+poKNRu+dtjpC6P
OF58TYh8uKe8En7VCGRo0HRCmE42r9egfXKXycYSfOOgS3FY2HePhbLS+yS5srDU
OPJwIbmRtUPjeUYmK8zgJ8gZMJt6rX/sGb9izqwK9pjeOITNAuoF11UPJ30GWdZW
fVU/rRrYTXOGva4inA9NvdFrG/DfFFXOyf/UE1grdfUcULp5HrCm+oOW3BwGPaVc
RZ46QQ4H/ott8vJRSlTpd90hlnRqXk7pU7pHMRSb7doTqDjUv17jnKQa/nGbdYRl
hRs0dnaXf2sz/zernFz3afnSip/r37VPULfUqWy2UVeSTR8OEMUdDB+WgqVYlK36
H478LpuBwYTrrYf3JNljnC/46H0vmuI39OUQRcHGa9BulKUnKuIoYUHdxA3T/g2n
91PZrJiEOoqluYQVTbmCxbV+OZXCt8jFUmps7Ycx6uxu7tnv4nNtf7AfdB84no8y
fZc6FtqhvFhrMqHnNNJEbCRShZ5Tu9uLMG351IgTqNI/Lqvau7rSexDHjNC93SwT
V/ur8dQTelqAEShQFoDqs2C1DCv8xpym64TPL829VbaK0AE2IWw0Zh2sacOjzWcZ
fe7gT1W2MYXMQUWUefGb3Swi+CO8JoE4hj7gXn9lex73rXLLaLGkcaKo+a6AAMQ0
687/qTqAlgwM4EBCozX60slX8ueFLC2uQpfJd4FaQBOx1vSEFcV+DzqvDR9SSzb0
yIQ8LmzsDb0Qi5bDsFu8pJkS8NYXQsUMPuNQE0QzEUz3jr5wfPn2y+vyUSNaIKvf
Ztq3oQd+9ieTdw056Dr9mfFdeYUGuXvwFlpMxIyKwcsfDWISTbFAdInodPKyCGaU
nQE7xiungRRqFYroP7q5hgn0D16R8lg7KbhYcfuTO4S2b3n/TAbLLfiKvl/NDBP6
A2BsaLToSwF4LfBgJ2683BCeQR2q9k2zQgtH6isHr+HxofjcBLRo0b8TWe1zH3ZS
eanptMGSj0hieKcLxY7YpYBhpu2mhVAbLPLhMRnQTES6qqz5iCFvLu/v3wa+wuqX
O3Ttgm3XB1x4AUgAS3RjnwAVsqB/bhhjvOFC79JJ4jyy0RaXn57KDf05s9fxyJ41
kbxqxOdJZIQWgd08w9UFHEJPD7JESoPp1zgtNdHBdVpNZ1EECR7ZK+kiggPAnhSu
/oi3LIpQJs/VmAfA2kb0LMDWXTNvqPnSr3es5uMCi833WxEy0J4GYf+7R0VdBnFw
DXge1+g8Ns5x6AbtA2AsKYqKQrMX8DCozgxCrc8TPVv9B2fw5+2qwPY5jURqdEQU
oH+v0yQpYN7g225VucG9hYJBsqNnBP3+N7/nbmR3l4BM35Qwb8koyDVpTkECwBMT
KxUPtGB+oiHSUDGTC6URmPFTiTce7f/Smhy+41CnZw9aMl5+OcVlt9WlWqtjbcX3
ITTT1520GtMdkw0G2VEqpiDqKdSWHU5R2Gi1FbuwaNbVmq6AV3fgSLvLSrFno4j/
BAM/OQtMHHTBnUKXKaMDIUIQL6R3Rt3eeCRbm/rRaMNtH1ypNiMHO/sfyJJRgjkz
JWYOLvZFebS7heURwe6DNzejLeEtfY8XqORUwswStTGLRbhMkoxuTxfcDHcQnCBS
j4oywLr/WgjQ1438AQeaS49tfC0sAXpD7RkY9LzhpjRviAjsfLDi26GwvC4hEbAE
WmtrfAAYRpNW0bHdk27MoGWBIcIxAHPnz1m5WvNl/oqBUdPeAMkbKUrJpv2dkzL4
vBoTzd+VpZmdaHfMMmHpUFuQo6WeeGNStAvUTujirmD+IJ5/WcjY34XKJt1jy1o3
H/TF1cU0ZJddAhBdRpMuDHlzUicI3+szaF2Znu8d5SG6VUSz+5Drr907GFX6GVAt
zCp5m3p5+lFGSjz3TOuPrcn809HmjEv0UmPh1UsbtONKlPpMJEAt+phUGKVQ7Ydr
Dn3rjJC5UTtsYtmIz94O0UTbwhG+ZDlpCCz0WmTEYUm8n75OCsLzJrXNFm4mQdcA
dnL9sm/3eSLGk+vMXvHSIls5Cw87bWiqjVeqqNWTZ4MgFYg7eSZYJGkI79SwRHa7
SHIu4vtaMr5Oqq2m5vXFKGgKPR9dKENoDThUJlXeMldeB6ixH9BbnsPlz3j/PC0q
5V+ylQ2YRnidtB8HBQ5oH0ksK8LePR/129JCin+H5l7VoGRseKkMYSiPOUghqdYy
oAe4hqNCORCpUdnQu/vTC7ygBFKOqyVeTihGSDAGtz2mJXEhMQXnQqV+vfC/GuXB
Yufxzgvbqr2RyX3M7s56fcIitbc173dnJQkMsGLL4bR/zoCeBQJtF9etXAXc21f2
kavdrKNy/VpCW7yYQ5wJX95y06hiej2MSL2v5pWO6pSoisG1rKoRUAUXYlw7xLvT
/Ld9WqiBUDbxW12F/JFy1k4YOgg9z3/ps003WC5EVYniJuD9i6kZiu3H2bFard8G
emx9MXB8Sx0+jzAqHFgvnyi7SX9cmFhOa7WRfIgcGJ18SqfJRJiXahYdMdLkPUYw
7Pm9ouKAFa8gaqfecsZfONG6sUIjJE9Cah5eXF58bCIx3SL+0/UzZ4k1rcAZ/ygb
pAY5h8jLfyiSVIvEBPl9STY0bQVj8es0/SipIS3pWYDhvfXJB7Njpolu8D9nRc2T
8dOQ3uBoCuuusAYwBPzaya+XF4XBBZEUgzOTn1prkxODdRq+aD5vNK/C1lcipHNJ
l3d1cRy/0KbGr4TsAC01F5i/XKL3HBeqtpy6hnrbTBmuSdWEx/2j1n3iXfNI6lYS
9SXkRa4ztjQKNHUTxtHZujvmyuGQ5MtCIQm6muazJzojVFYR9fzjMfiiXVWDpI6m
OIuy6G/+MIx5jIk2Lo0kNrPm76L8yxGYZPYPQ0PwyjOAb96Wfl4JaWTOuB+X/ZgZ
ea84Bd8oUChsRBPw2ChrS3n0g04FJQUXnXxbP7SjTVmo3YteoeT+zlLOIhNa0suq
4hfU0EJZj1m607selDMjkkRkr6bygayJOT7o3Uu1nxNPnyce6K8ZswE/SA8sDwlI
tVRd6KbpYW2AzM9hOA/kOL5RIjmgAjzKsaoyfd0+TzaoR93CNgDVID3VwbrD83C4
E5xna6/DgMK0QxgkN+XaffmPF/GRMpLbmTjGLQ5SBVl6U5TRAAdzMFzRaciptr0o
txCEYIBsclKDGMuzJ/l1TSdX6Cbv6LdROv62WNZQU/Mn5TsJnykiMNNDxNV1y2Mb
eh2N6pRH6wPMzmaXYujiTPFcz7FS5my1hVTGXgYkx/mQUO5ghMoCEaDzmOANjvCy
2EABEjA07agTjAw/NZlFo2MiITyFC3BdIVuITFCOyURIxO337bBx8iQu0kiEZ0HB
sBXzamN3iNMQwPvzdv/81P32zq0dhUu0c7EjwuVD5k4yESaFEH/qG4FxHGIkviz0
cGaUnLM3RZGXW1k2pkv+BfRLMGwcSh/MX9unXcFuj6mzGMC2vZ0F9rtBQvdO0Al8
SwB3LBPbiQVDq2vVhMDNX2J+6nVgoKEW3t8InKdL+OQfHqEbf8CYV97spLdG70oZ
aruP5RXkURuQd5kxf9609LU02u/4X04fkO4nGqKtRV3JqOZy4ipP+Y4hdVRyMAmQ
t0qAchCX8+JGS8/pY4qfkH27BU2P8Act0GQUBdeeAq8xz06pozL7YMNd60JiWJ0X
WUhdlgANLDS4+WCzZHeq7KcT79VWO+u8lhkJKtv4DHJweI6LqukHOb4M1LCyZC5V
lbMmtGWYa6RHtyEfFr0sshSgfkNa5o2RHQZ3GmQbKJXyEjz7AAoKLx+1jDB+6jSr
r332efKBNKn1yi68b4iuAOy59i2IZ8sDunaTBBSrJtc+8gMLJIABk7cXaBKNfY6f
IzSfDSvgJ44cvX0cfIpMGUl8d4uZ/yrd6WcVLtHEiOx5Ckar4FSwC+pw0GAPudmn
8XIV/TUAu2awwg9B9uV7BYjucyhsYv0GDPJuPinnWulCbfwSa4LCvCCLz6m4EhL0
7zP9D4TPUHhIVmmTeeW8efsg+HxCBsNwLL38M6AH+N3C5oLM8qABmh0Stq5zQ7V8
ydtq/qf2mO9O6fvpNiq5eXToN5L7LVup1CKUuMfhhTwhbinr7nLo5CggZfvIfEIm
ijIHgpCZ/55/xLeHKUO4NkCqEGastS07RX4rxUtS7TG4Ok90/n9uT9yB1ojvmDBr
fzL9CiSQLez+OJcShfk1Pvc3wH1OMSIWL09MU2Jc0Xh20bhluWWhGGY5NmvVpo6y
EdQWCU9hDRF6AbE3Jt+IeL8jIp9hZBPbryJOlF+nASNRR2004oGJo1cLgP+fEt1L
smEZh5WxY1PnGYwUsm+8NoZL2iJF17giOXXjfUnZTOTdtVuOb9MxLPjyvD+vK9/1
KjUhjCWghE3Ybf0cpQYo/JpBSRF3L/YG3Tu9yxFYKBCJ8z935tfMKQkKZO2gDO6Q
E91YBvADK0XF5AQsycXB5M41RLacKGaUDG/rAKos0MvgcZBMpjVC0Ogu590+m5Xt
gnUdcGvd8uCF7czAy48k/eGE74P+Z8aeP+ml4EId0ixloJsaLmFxnL92tb18hWl0
iaUOz/QFzUcYxI/uhR2FzaTs2+0yHrftDZCR8iYNAPfdX5C3I8xqrnjG8M2cbrBc
kFFt0aBd3FJhPAnlLo2jlHlnVdpd6R6x5DJTP/z9pzNUnV4y3pJEFwwVxQEIjzEN
vDRXeLY7aSTiXsg7QcsBa6S4sCyWWeTZzsxzHz/NFDNdkw85lc8rZfaYAfR/58zx
5oQ2sasZI3HGd1Zw4GtUjiWnaYwbYrlP1FaeNAVyZz8d23Q2mf4x0neA8tQfC+7R
BJ9z4I3eGhlKkIQ+sW48hgWIlTmmkKgAEeKEo7PSBt2WAKA1lFkWOXNjWnNL79IC
QS1i9KEx7C31Zw2wuVbqU/473s1pohtJFbKP7/ZRq5sFztq25v6e1obUbONEuFmT
ga2HYIw5LepORCriiZpbwHkE1/VqZ9xjfzpDxDFIJTjfJjsm6DRUIIH/jPojfyU+
OQ/tPR8WOx52lR+IMy8XmSPZ9sigRYJ07K4aGS/HTzdNpViqGH9WRz3SdmC8OUf+
azGF34zJUif7PXVUAXQYD5PTDlmyDo2xCUhj1B4RUkrreDvrhlt1DWGMiNyGMpAR
/3KP0U8YXbOIueF2IY/0FrbyPLO+kWoTNke2JVN0+vI84rCGHo4a0RqNz8eeFO2H
XczKgsOITvaduNQ3VCtgwZbociBFYUGLoyAjy2sa08eK3A8egKvqLwZHXN3xcVqL
os7IUCYoaPiFHNj0k2mv+KB6LNq5hLOQFaV+l92sTZ2rHo9blhaqS9ZKR7lWcn0+
AjCDq2oYZojckiPHavrSiJDMyKhRHivofMNX1rcpJdM9dRGLcrgLvW/U/spnCwiI
EuC4t+nyCGlGgublcSemofoTsjRjpvj1zEK9gN/0uGVegv1q2u1eGW857+uVv4S8
NuNiKLWa01Nc1NP1OkexwqhqvWERke/Qyyrb8RPUkPoKLIAQFOd5aYcFF9ZB3YgK
Y8H4ickc7iLNryAYMjD9PFCaBHuakaSfYzSMb4OIoT0Jg22NXyzzTjITgrwGi0o4
cblKsC7ojWZQMorVT409+kIHW3MvF37nts/wllFpJIgvXOaOjdO25forI1PIkmcG
ffJssFrKnC38z3K/YKWxcOWk/PGmpqEHkPzUuASaDBLB2xLkFSTnYV2n3imL15g1
2EYTbURStrph4ApC0mkmdpQvlr2p4Owu7NwiGF0z6wa+bUQajJSbkqYyrmPbvNQg
D5y1KBQQjDlMMB0JxtVjkfg2jX+5MSFTUBoEGuBAJSNwMKtz0BzaFJscw7YxZOpA
0nYU3X/7sHhN5zCHMqjWiSd3CSOUG45AgYUjQcOO39De+U1rNezwfVniWoPa5hax
L0j1a4oP9z+JicaF8MwPYnGoQmIPns8uD2yI49kLnCmBOz01xtfO925TzHoDDku+
uTWLPFA3mGGxBoXPMG8EjdX5x1okyypplZc4tFXgoBX3bEkkaYHX9WctMoYpH6Xe
TPWFYgdY8nJsl8hqyRPwsIFFBdfWs/b6jj74e/HoLdIiWoLfLD/YcsRyLFYelulK
oe7ZsTCFl1Sd6QtGK+eA6ExD7pKuZ7DLFoB4Rk7t6zFx87FU+uis8ewuVdlc6K3r
w/X80JLjZLmTY/MFNXbajAHCO8YdAZpeMGBJgQH6wr1+VukyoUTHJ/bML2F8T4b1
YvhjWbTuJUA/BE70nkrspqxLfisq8g/a8nklsgiZ307678Ek4M6blK7uQGpC2LBt
z4zMCyLtOqOpjqi4wzAdUQF2QlHVMhb5VWcrVfuwLDYfb3psXcT+jidA2TnqPVW9
q7Ftc7g7NI1sAsAx+jIj1C/4iy+056AWheBWVIBvPYORSClKTsQASFlxWQzs3XG3
CmjMYu1VlMN2H6Ii703DDybt7MAoNH8v460ygM8W9qFDXZz5faKfNgoQGAu6PdDJ
aFpf6BjChOX9HcGrEvkgZii7M9k+xhBkLZYPcRhbqInl8aobKtqPvOpxMUlJvFEQ
t61SGDN3DBOyGo2nUD8T2F3MX+fESc4efye11CLbMtzqM7+/pH7IxB0SSw/M9/HG
wq9t/6WWvmvSvpqnO0vIdzaxO71kmw1xlnAR6UlrjLLFLPiHcJel41f0SXMg4he/
qIywwrt2JqMaARN1g8+WHi4nDML1rn1+j7JQEY1Rk1snGwfX3CcO6w88TwXcRe+A
oSD2W4RBtMw2Ph+2TprNRQ/HHSccoUtrbmYA9MB/D8Xm0wf6cUbdoO09IFWO8jlp
/mMYfn7oDLf5nrbO6I7A/RP+KBuPUo2CuAuC4unzD50by67GYz/X9BFprr/co1nZ
cKD1kSkqqSrZefA9lKeVyG5E/uGrnh+Ei4z/CyxSDOUrNaoHyrfL9VUm8QTLUfAg
gItuPF/qtWYFHv1xrczEoXXf2pEhVgX4XYZp2nRwQxmCoJ+GuXvhCfzY2xTI2wq3
UAgYTfKRGZsnza0Nh3B7gJhVfZUKKi5tcexmLcfCyJJUvFP5a9ASRqKSsMcf5euy
Rd5qdwRqX/j8lFlbelXn1te8QVWuXPTjrtG+V1fiWKF6P0VYsdx/YrG5qnWPemk1
b6HDNr+/wekh6py16AgtJ345ojTAKXXN8yABmRZKnLRBxdP5sfYPKHHcMoiRwHLa
5+vBiC9eMzX7aBVDdNjjULgm9EiCmSKAlwksW3Jz81VIiOPrbBOFUpGrA7wD2Sil
xnzU9ObyQWzc0likYKzbcyYywATQ3gFCvWY6PkfUhhYtMlyom/HBz5qsXwBqLFgO
bsL+hCccp6KjOCYrmfwEMduHSgp1RcWiazcJqLigQXR7xDG6/xQGAnF0XT0pc4oL
yLVb0yOrOpHqcBb/WaM+CH52TeaWqh6fivh/T5jBPQV36asdJqKPPnsL+Q1Bdqyl
7Ey7bg6hmnZKtNgBYorhQ2A08oHciAC5IYIkFtvVAaymIVAf0Fvfj1+oG6RuPTKr
yQ+0N082x30FjAhHJI5jkR/KYnA+7+FxTq2S4nHt9bpFxtllzUGCbq0p9t1FTZWi
WU12j9NxqKH+tLoYP3Aq3zmj2zxOgtp7n+PJXAxbuEY4qxno71/3c9ARS2EKeMus
OptdT1Z+A72YuOYuGjqZVycfPS/aCBxqvUpu4va9m+j/3oD9Lca/GJPMxe281TRD
d6Zz0Sy9ZGa5/4Rf1fivKcq2gk57j7bKtfO5ugTH82I8UklvNhXJ9l5klCq9GASB
bcbHmRndT3u8HNFNrl9C+3gjayrsX1e97Laj3LhiKGg5wzTFFElb9rG9dVltj3Sn
lGaLwJBS3Wfofd/R6WDgSO6nJK6Y7ZRh203pc64pGjlsKawEOav4jBFKriXCNIeS
SNiUexBBLxd31O7JTf6EMaWnjkJTVVIaT3BkMECe4EgHgI7q1x9RzljU3yqgqFLm
5bEwT9gWrhuwNzUh8GdaNumW1DL+2ui5y0iT10kyHSqT9M/QX1vWsL//tQvvUcrn
9uKKLK0dNPSpn11KDfwALTgW05xqzFII/DljcaK73zGRXY7/EAbPXWSCNQnBiUTe
0UsEgAT211vKvN+9SqaGkFbvbdYkHpncMyCaC2Swuys+uS43nWziLHzNXUWnX6uD
hiiP13XOuD+NWgZ+GPbX8MEV7yg1Sr1Jy5/ho615L5lYwAGojlGYJo7xqw8tgEZt
zvTJJ/eKEmzCcjAPfbqTko1ozmD7BqXmzT3uUlagXQJyqm+y7ogF1sMsxU53Q8Zb
JtjZO3D/EqpGgEED4//8lmL1VyG7OvswhGYj7gI6Y80xZiKGRgEmkg0TDJggkgBU
QY6YEN7V9khOV1olmmHgiAKLQIYbFiFIKnVjJv3QjfgOH8iOaGSHGgaWJrn41wtK
KuOXJB92hvYXXvey4iiRTEHqEBEdU9YF02+bkV4b2idTc3NqyeqIQxDc/pjz5BTo
Uxd8hw+X/H3Lt7VqjuziK8c+xcSD+eCY6OuhHIOgF08uLIE7IhLnnbes2cRgi3Zg
0dyISyiSE6+CxJXAtwkJ+VTOk/tZQAMcpnHMF6VXsB/obx1foqZYxVEQy6jnFpHe
8+8mlCw1BCX8QWrRrYCxM5fa+pn63YHFfYQFvCwt1cahWBN0s9h3r8FGJBkstlkO
Gm7RV47OMld2TJaAsh0xaKEFsJCM60QJfP3vPV/bUM9h4s882k+LuWIU8BXuVdtc
wYQmjJ66MaS8WLpjWP71xrTwSQaQC2EQjkkMPyZ37qqniPvfualHYdIpnFInAifL
8Vu6wI3NV23mh2lmsEVXPY3ay1penN/w/NTnUkWBlGUAAN+bCPkCnI31hd4rqBZd
jNWwTyLYf8CoT+ZVCn8I7IVi8IG9UK+niFS07xyOBdUbIoBvCaZ719eHDiepVoct
lGt181DDw85Sb08dXqyXjkvn4H2s4FFmhBA688mtjythZumNBDwLvlSGkCF0xzK+
4sTicwWeeT+ztb+7cCjHvA2ZxLnHntLp1I7wQMsj31NvFG0RUW8gvkW+6u9AB1xv
pzRXfL2HkYN4ZlZXIFjvMe+ItoMVHAl5//WoQzqWVQBRKp9eWQZJ35qp67J/Pwkj
fBskj+hU3FgmQonlWdRCJS99WyuR1yZLHosUAOYxlCwmp0T7x5qBWkUPggykxl9A
++be4OUs881ItDubJ98OgJi1KVGDemf4vJHryyHPz5p+dncBqouz+JbjzqLcNk1d
nJ14KgXbD7Fcx0K3ClNKGZZtU82OL6vYBdzkkazFsI47Frtq4EOwWGcR87y0FKUX
OwXtAps1IQrm7VJs1UYc2zK5JR1hdCSM5AI1weKLgQtKPvwT/x5quzXiZ+Fz80m4
fC5jSAD0GUC9ESj3Wx6XMFAd0SVTPohkX4dPf5Sp9jsxsrFGWTVucsaYx+YehbzC
PSocEIZ2mofoy7cwWjmg61xBJ8kpaydovwJJYBIe5JKKS/wfgvwEFLbq7UP5GUlL
1cvrn3FiPYRxjThvzrJjFYgDHoECoYPXhmpkyue6JCX0A3gzf9QCah9AwWeELYvU
UMCECSi2VVYDwrqpCI7UeOG6fMy4Z6vM64Z+Usm6xORrnz5zlWYRAtqQ8JkUgHeB
qGVu9zNIhfwhp15hhbyMoGWRU7RtgVEPzP31GyvrfiyWAnOb6SisQqevgplHWFYb
rto0SYIcrM8059HFHzfzDJ5D0Kn3pvfFl2LsxjrAc7GBgd9+SVAshmH0HxTMZOKP
+gWo1FptGrEa3dI7DLRk6xDr7eAyvHrVMkKpDMnD6lx+81e3fQPL9umFek8lV6M2
F0TQTMM5BIwuAKQVTSK5pDbK1Vp5qucG85u3h49p3gYgP1T3NpJi3oj/uhG+gfX5
Fw8Gb1B/u5MybrZA6zvE9EnIzNBt5cKOxe3Z9xTomB1NOPj96QgqfWNIzE4Ef/Oi
nA/7i2jkbXygJnwN0QcQUUNxExbw55vcYV5wGRMm7aliiAOtImf0N0iVWxJHw3tx
FNBMfan8rTLmReM/XuAwsqgzqUWlyL7mt0NbKq6UnP7OWfXZ4HUOJKgjHLRj2IZx
iuNg69WugHyLeclDMV1+m0z0Y96zlmvOEkOqdsK/x9NWGpZG9kOwASuOd3yi4qXN
j1SUPHGSThBAtP9Anj9mWF/MAlJfrrkNLtYyP5ihL1PviGbveP1CyJL6R0BKSe/h
SsxkmUG2B6KwhTMU8if9J5Yah75S9xKddkHbsWCY+GEhX55dTSCSkMoclL3sy+hh
vhewS5vyZEiSteDFGa+MQjqSz5bFcycEeJH7PyGwlvFnre67ny2zV1bpLB/Hgusg
4OI4fp+Gz4bsD+7VYOtzCXsQQw7TUHeuycgnRV2s3uLOaR+iA2uoNd+4SBYZNbdv
ZlxPVPskQFvc8nrHVijPLv3VxY+3Y38QIxnhqxZehDzx/ucPpzWa4WEexAM962yl
bEEMD73YZPQRzyIHtagh/butQKTEmAaNymp2TNoDECC+H3G1ICFgKkPgDEZ5VTu1
KDV7NXxmFOohHrWuK/S76FtFwTJ1cloXD00YkGxOlYtLObRwDj/lugHfz+jfq1N8
wR/1kPv/GflTHOChmLKlaycAkq8s+y9cRXcl3ie6Cb8VwuUPGacGbZUoCTAS950q
YTFCJz47DLcXlixI38XSlXWFr4tZzuHOdsJDysHwYeUzH62uTb+XTy5LHg/42Xdb
gPXFOevbs6A1i5sbuDcT+7+hdV3Qxlpwu1UlP5QqnLb6HRuTvYqgvPEeMhqqNIvc
Apxrpa3VFj8lIjKyQAqA1b6joj4fp8x6n5dqHQHTm+E2kXFbloQSlX8J723N02OE
sHNEljJNnNlpG7u6jnEsGjceNrvleI3D6qc1oV8wswdkHcKq0PNuHdj4gE0vpx6g
qSmLq9Std6mHbOugtG96X0UOXYN/S7b35UrjWW3J+dpZH3FiiHarg9PDs1qlY43Q
VpReSMqxd083g5FMRbj1cW9htQb/VXj5M9hYWC1uyv224V4uzW/PmDyum3UBc7dY
d+ag46AeatCOwpsNkcNOolypSrGGKwu9wR/sfdlyJoZlzXqiGbDimKAtF9vVMEjw
1sW0SbynATi6TUrxUzIWKQE3fIDCldZwGGgEITiPS0EhGcfXhESvkRhPj8D2Q6vw
XV8A5n2fnDwrG5daDMK5sOgMa8rB2POKyGGgrIbmUArALThabbP5JzHnF1HrePUt
262+zPmN7hT9sy1ueudW7mhpBYUOpa7NG0mTerUJxW7Po3uNdgHUTbYwy8hM9Yxq
1WSfHl6349ujIBCcGYeysQVX8ScR6/DcUnNhQohfGR5b8sSrxo8tm9qYLZPEqnYC
oHjxuyqfRVNRd+fV8IVuXmGxsMHmmRGvJ57IuAkAfLjM3qN1OAjtrQfRt6ewR163
zp8J3+7DmT+w8+0UV3JeKhXKM/7+x4Qc9A+lxXHBwV6cDe1fS+wG6qOxLetHFGFk
I1CyX6E4k4cor+oNbiPf1Z1kJgpoJNQ8L/RR4fWx07tCHi4McTL1SHU8ScX6FxZe
lwGKZV3VhEcWmpxWidnls6nSedMRj0x0t/bLF2hx9qCv6lDYrFLM/zgcXIsB4wKl
alLdKx0tnofr5Aj7Rvfl5WpDu9qc9gP+H9WvQl2H5EOn3nx6FENKCl8s0OIOe94c
b0iZ12fQYgXyq4Aop/kV2xgsxfaAPQOpjjJtxa0mKrCIZM6fSykrqUVJ/JrsNLEK
khchWzwqWlbA+gPx+vzHTO1C1bqkewmPVajhDFGDr3m2Fb4dGfh/pMqXQvZjUCKs
QuN8ypgRnr+pMxQYlgbNGztFCiCt5Yb8krJM8WWcaQL3QcLBMck7GU5uZcCuaEEN
MhsCsjq057D9+qSYqc4HDA6G6dtCzMQAdY3UrVRwkopGD9u2UTTqdU8P/UUldnVc
Wr9dViouXOMRNrdJD9k9YQ3SIMr1fHH00Sq6KxFVJr9nvqcBcZkjF5sgHLI/iUSt
Vwo6mw8JI2N4PKeGV+WKoc5xStCk7TgOEp6sTxh+TIHhcOIFAqUjXIH/d2PSyXru
6XYWSzLT6tIlhthrqLuDZi7aR2LYu/5Zc2hamXV4n5CIZOzxkI1sDtTNkn4EsXkM
yJTYDEECWaqC4RqFFxMNtVBtrCvX0g1dUXEkvf0gti3pVFMfYmPL+hHosa/Y9v8y
Hc8ni4XeOlpH7KJBGSyqiZswV5Zv85Jv7a13nH7TSNXTeVQjFeJFBm6J+Xxz52hR
3eyRb73xFFbn9OTxapabbuMXykXi4HjlHNL5rfJc7N28v98uGF7K+tx5cr9seDnd
grIKxqFyNE46SlNPwdCIaw9xt2OWY03rA0KtoxKDTcgt34fAZwU+EC/F1wKQudCE
USn6W6y6B6mFcUi0f062Zd3vWS3uGo60rsw4pkfx+J1i/9RaClGvo8qr0iPeYKME
pyTDI11FMP4R+vA1p8Slu4qjCejQ1FHrl1L6nmcBDjZyXFoTsPeld4D5/4A7S5cg
b5zwWMJKDZABBXsdEqJGMdwY7ZHaB7+Fmi4mi4XDo/yD+l5C3vs/ZupwXE2R1NWE
TSKumBqyMgNurmtk6bREXkEzBTaj+pP/lkbMzCaeqL4rgk7P+oY4UfqacHzAD4+o
jPi9bdAI1PAuL/+7Ll/PFFw4j4G3ecXIjs0WlakCLDdBBT3FhLE3xz3sqYzowzhY
Gne7Hfx2NMIqCjzQIsAtCmwf85pyEIfzxuvi/sA41XTtNSV8e/gIkMV9hXx0QvPA
hMUqFf4eIj6q+xoUrden93EAYt4roeUCiZb3EIzEl0ry2Ve1zMJ5WCh5qhoA5esd
DRy8clG6rdfhY1iJ+gJs9WczmghAeHb8yvuykR6U9hM9XLmDsUpWwJmSB5EdeKGT
Z90g5KjOAk1h3GLDNyBFlRUv+PLo2u71F8bPeTZQ7rXz9Awmt8p60JDIuUXOBerm
uwpcdkgWl7ljB2y1x601+raylyVUnC1RRVJxZp9Joj+MdmdnWZ1ZGCI5SWlXxlSh
33XCVYsj7S7g4hVM3CZQZc7O3+Lapc9LNHOK8LlHN1ZxyscoRv/Pqnz1kCbYPl4Q
gPZE81SqrqcKlWEtnBQFlj2lk3wtUpPanThgFwoOkOsM4DPu24jZZSaiZutU0iwx
CcYbMPwBrod+wRe1fxrNJUItS3L+3s4KPNUxpCtiNvfhx/70rWrsvgSXeV5XAMAb
z4wWjMLiQu2tyDwqu93RNgiSSqhRnDLDlcHts1GtNtuuGYvWNPELlGoriODiVERz
MK6yV3O38YLql/lcasIWfkqK1d8oOhSqzYCUhBhX4Cln81KCWHGtv91LWO+C8tLd
Pasi3NEt2oTdHaz3SGTvsXmwuAF8nuBetaBZRIOw3opHPM4Gy3KVBDjA2F02rr/g
DFYDbK0J1LtBw9Y0mZS4ObhC3bRtWFFdCxnhL1TCXEcxYgq5gfxIAQN7U8kR/sqW
yD/G+B1GBcS1e+cTl9jG7LndCu87hxz3aWtblXo3nJH9fXYeWIFMbAXjtZ6ndkcG
7fTI+wV56tnNggnGV8qDxQMxdGxG7ijoYSoiQqQbLDPzdyXUqKj5EydV2PMgtqi6
BwaY0gK+F/Z/86m/d0D4LTO5bXgs5efy6gDgTLDLPq325GlCatvWhXWWiTkPecjy
l20bTVBthbpX9LajayGfc/VzVsyVBiFpK9s7o76UrKfY0rYeoZAp03NzeN5RElsF
rc9cAERCcPaLG4GsG70GMzS4f9RQpNLP5hQRjNHT3D7WVsGZZIDLezUJL0xIH6MD
p8hvn13wMf3Qfo48MWRznbJysCtxZBMiJ1CbQKawa/xohGzMyQWq5IQpm2RVlU1+
13MHh7uIKF6xdoKq/t2SXGMJpWZqQnroBs435/3Dc2TD728EYmeykEf9Eu6Q0kXz
+eLXoQ8RLHMsqbdJ01tF24IqWfBqmAMfVmwpKP1oeGTVUdaCfkl8zLhHC01UwP8V
FmuvoDM+yPZZCXtKD+llyJcvUDHJakEuzKvNnSKQedTSyesCA0NfHvGjboMvwruF
t2HKTokziKbRSxcv7MpTJC46oaK6hJUYKv/S659fkyNGa8f7dbByM3MdjDnIyzYu
05r3yoVWqrIUiRFUsZVWnoRm0vsG+Xo+IIN+vBxWjvOz6pmmJkp90aJ/dif0W+0k
EeurF/bGkogXG+CRLguTvh2rRBuOp4CijLwvSNyTc2a7nxqDASWcsLP/5ufr1T2E
XHbQlRqurw3UfXd6FwhX2ctdLmi+hloDNsAH1N6VFvZMmykszbTIrX3Sz5UpIgl/
xfU0jMi5JcTrziQqb1A7N/gAN8dSf7pk+jZaBhBC2EHLKEBCCxrHfLBRCmf3WaJ2
0XIrUZ10Fzj8X3209VvJ+vB8brekQ9Yz68g+gP106ESY2IhqN2m4B6ELqZJpNu3Y
nWdmGa+7j4+scNzmnSIc+sHW/fz9z9Ydcz6NnNBMV17O021epYOWoUhS7wnB/Zm+
haakjAeAJy3oQuF9ZQR+GIf0WikOaokHNmb07H3YF8eKvnZ47VTqoUt6u704uZ+a
sTPptMszPzF7NXTR2fK6Kl1okXpX3ZJS1vf1QLTRZzYvlCu0qfofiK0FDGYH0zSi
oOkMZ7n79mq8eiFfglQs4n5ANrpjDtCCfebWFGQL15Teq4SEN8QabdDiUphPqW+H
g9g2pXtuD/ADB5sH9E4StGFAucaO9uWH9UkKbM1DHLaz3AdNI65jWeSWLu9NDQ6/
koaq0MyiJNBM2vD3yuKQRey5UQRXTJL46QeobVmRrcvubOFQ+5YB5OVnDKgqcTzM
pC4LvQsmxMvyrFWJO3/GzPmxeZg51CUmOAo2Ol5jhoqacJxHaAix2WqrJVg5eN+A
5OEAzHkH02eLmTlgdKXMLobq/jeJh6Lm3Q3mM0HysiHqCdjGZ8pqzjrtCwP0wjrm
/Skd2qWogKr7J64azUqn20pK5Cqtybm1DkMCfRptfTgPxR2cAE69QiB3mcpLbh+m
ZJ3ghGrefGGpxbjPa9p++k2V5d2HS/zfo9XI++Pvu8xjsxSH/3qN2B8mZ3TzCaQA
Czfl4y2Rqr5i2tqQV5zJ6DVNVrQmr47I1qAPi0L+cH97aHKfFcHooHA2gCYD5fC3
R1vaI0gGfHVkz87dj+jXhgttk16IwO7SB/5a7OvaFSf341bQER2f2ANQImCU798l
i2iiQjt04v1Bq3LzI7XaJSVWd1bCPFQ8CXtswLDLbZTv9szTkmB4nc7bkKodYgYy
JwwOKd/u1cg8VMmMM9yk5b3mEO85nXfc16EinGPM/rQ8AUjQPacTtkBPFn1qk794
Y5zRxG6HXDtfy5UkoLD5aTEBixX29YtiylS3qUzRdC8sJGJ/IAVOTcHvy1oeEGpw
hSsQ20rwyoVKIyBI3+MUrdTdtqkIlxZGx4L8SHL9yoEHAmqinasOHQFHkJ4mx/C3
Ayb2SJJ5zBiWu9uL21mCrUc+HIuWVpfLjXPVwdjy7kKR7GSIe45ytCi3A2dnqoiZ
cGMy4SKNwqDs3iSqFoiK0s4o+WQblGyoJKRzg7p+LvUAvTwjt7/7YEgQT1Tq0e6v
85JAM0BWJBYvSUBAV10/rL53h97sEHYpKMNBrwnjmJOXfbLNirdIgjqh5c5kYVzj
kRojULixpZ/DjCWbOmihucxT/BR0tc3JwfivB2mQcXNCC7B6YiZFNvm9OkxkATT6
6nht4oH08sLbSxB0KPRz9Y8Qz2s8xZvzpZ2MuWUX6YH5ZhL2/fUHLXRy7R7HPLIr
7MnbddCDKeT61V4ijaFuJjPA0LObWy4gR5dyU7MZfqmcmEvQ7+GIgIK50CpL8GkB
pS5ZU3aI8YDqfXLw82bFX5KU0B4CAdldRXxpUAQgLUK1pO7gwCM79Ta74BSGBJQ+
JCKHeo8kBsbHDjslVf5bhKCcK0Cai9e7QeYlGvnCNWS7W8Yq7dYNpyBmZkqSpvuB
Phd1L1tRx6fNr9TRfH0cwhvSliA9mX8GydnOoLfamqSHt+uG4/oiFB7CLcvw1++Y
dB9RXgMLSQTg0xZttPVLrGynrzhLW4iKheRtTncYs5K0DG58dJPdNifOwufVKJCJ
PObHWmT3uyZPlZ5yDN0VIq+R4VJGVmEUj2x/bpEo/I8ShCNaxbzW4b7mxxhw7/oP
RheD7+p6OZGlBaLinz5y8qKJ0pxLX37vSH7APkSze5sLwMR+f4aivZWNg0Rj0hGN
zMZjbDlH1Juoxb2r8z9zmHRukFcsvNIHrX5eIsJnsJ/sCWrBN7+DKB3+Rf8AzswX
wkUU7UZLnIoaKTg61R8eO15QiVDPa9088j4orSqShxgpzFzkY7746UqrnHSTqh65
qQyP0XOgr8W9G+gB2NjGo/zD4o1w7VXc7vDY7Y5lXISGfkIdEyPoDDbwM/u4YgO0
cpfm7D0lbBnoPwTBUNLVwINJtS9ygbVIx95CT8IeFnHG2PQpNbYgKelIfkHKj+xr
eNFz+ShztnGGQHXKT5dtwiml5mRt+h3FJuLq0gTHEmw6lE53wRUszs+kBP0kou9c
ig3/0KcKi63u+eUJF8K1wWnoCgkdTmO10jwoelwAHA/f4OJWag9DIeq5WmwT99mt
/XMjvxUDwNKTtmXGQ5FpXRUtHc6oMUFtuYfU4bdJ7u7ftw2IvA8SbCSU58AIgotw
TJbohPu0ZAhtwCkobWfY9dSeYK4uf/D+9excsQk01deMXissPKvkupMSymFwFW+e
AuWz1swyKbpaypCxD1l6Y5ATyXrG9lU2ZLUe1aSR3RkkMvEoyg+BPPGW69PLC0G2
EA+LsGGEfwjcevO0j4EXRgtDXWkMNoQ0HLEGijBbQnKhciIgdV0t5UngtFec8Ayt
cNS9zciJJt/HWEwjsHCZ7HEj2IaK2W2anas6Oc/mgm+2EA6IIhoFT7XG1FbCfFUY
7gOaM8YE3G7Qm157PwK54qwCibsNvh/KgPNVe5ZNZcZoBUYplSA7h1x4ieJpOGIV
Pd5MIsXUjx5ohH+jAEfRuxOcYHdVIGjG2hHgDmky/tGkFnQSvETYS7tCPkVEWUHc
5k6QWPsMgbOEgbyYu8KFj1PLXUicMo5eOEJES6db84i57zHHhxUuLxjX/eVXGMpW
tsO9ZqXPDuvTPc6CxJgwyEVUmcp9bD7nLAvBYLGrj/QElEVNimEtinhAxIEkSmcG
S/TiqWbCTQgPBLAgpRdb5M+ROnfdF/WmNpwyyk8OxSfGYsZ6myLynCAl9tfHtsVC
hrqKOl319bPeT+5lNWK4v71eFHlI4juCKplsCz2JtDSrml62IhGsUL5KYm9bMnUF
/teZ63hGQPsO2MaLbZRAbKDS1mZvGIf4aLWQ5BzpwARJwTNFCfee5gQ2cfqve1jJ
lZYlePAqtMb0WwRCOBVBdAX6ZIR3F12V/caCLW+2YtLNXOOFarHvxdSMQdE50b0+
3hid4AmIXh1Md+rCUj6Acikecna0F3jiGvtSWdl4CsJi5tkbiPRrtEr318tznQiQ
HGfywjk+OXklX8piljSyctV8Zc6lIP3vaLoS3gcgd6J6G5C96/9JlRtQzXBezejq
m6uIuarNvlPS0cPg97kp0eRU7zY1tXUoXcItYLzsKkg55W9UPa92kh3zuLHe3QFz
2MDgzZXKzYjkjWUMKbWxsiLuN9bCiOjrlouMDivGDFT5KK4zQyN1j2A3kseu2N8z
1VsRT5AFeyEAKaPUsa9e/2SY2X+R3FTbuNx6uhaK6PthJrtKRo6k4kNCY7yDPnWl
DGwFYXbY38RaYcm0LRqbeamBNtlXIyyQL4ACg9zIdlALK0v/+RT47j83jlfVaT+G
vdB+bi7Vmxebi6CTpfng96ybn9GkhM4dNi1+9MBOKFBsjhu++l+nctsZ5V/CGxJZ
1jUvj6ogpypF3jMi2Gq64bVZvSJCar3NpBt7X8WX6WD5hTYUvDIlFFC4Tg2tw8GE
AK0JFatwktMqVIxZ++/pnRcs2NTACpC4D6A8WUYqvW2Ol5n4MNHpTSPEB8XSAwxj
jwxbpfAAQeyG4pW9ywvso+mUZR5jbQM+Ck2xXrBVMWQGCHWPPStj3oaqkEX+AJpj
KDhH2nyfow0+8Un96m1XqJc8TQwLIH/NrlAwzChJh648sdNkK6mKsG/EGnbox3Pv
+PHsECxI0eUDJUDogbJSkvaGZwuV8xG4fNeVDLOi7u1N/qelb5tVh/ZBunRCN3UN
mQ3m3W1c0vLQatOwy0sL4BuGnon4tBhm2hXLUDu01KNlg4AFEZceLqOm45rMWWMl
LTyd9UHi7r7D7CO/f6M6hc1sY9l4sExq0+ZpK5xmvWD7IS4LwAuspzvX07qE5NzZ
y+OicM5Jf0lCpga+kkzZsCZw8jkOiCs43k3vft5XMgV2n1CJFz8lAKrL6sD5Gqzw
uY+OQ6grp3W6TDn89hIN9IQbfr5UOoroSDwoiM5cN51cQckvk1wxqe3QywSOpZfS
nhgK7yj9EeTE84Y9sswB4xnILs/eS1OawQdkU2VnSeSR44HO2rnlcP89H2/Akv7s
xoTUesgG5qNrzR+6cGTsGXXUpFBtBD8pxA0xkrohgTUomhwFCFTlKUOpENddMr4c
US8DlsyAm3poYhGye7K6lcKaoVFeBMg57gcoJySp5hGLvi9SPP9p0mVMUEx2wf+f
kVoFyZJe+ARR1vvcN+VO0hXIIXTgvSUw2+/7MW/I5pCiRqHMV42tTjznUCE+yWFf
6BG0eTUQsbG7rASStqP/6rEd8VkwPMv523N6Tw157Q4swkut/dSzlSILwsOSjmfC
y/iDWvYEgRCW+qUQPj8PUr/z61lyg+lcajfBXn54y66hKB3rNmEb9T6tHQV8arLv
celtlLi7IZVyO8Mxbw7s8OAjz6EXyBWJcFy+7QC2rmCi8zemeqmFFR1Z3Fc6nVam
zUKZSHI0ZnpJ5V434lRuZsY4zx8s7BoopkifyrrEySxMu/u4zX2vyGXgZ6oL15JZ
9CyRQmbugC2baAKUQrwbRoqT/vIyxHdGEka/z6vsExV4r+6F74GoGmovaLI53gv1
QDG7KxG1cJRJsGNZ6z+qdUAFZsseo4iFLk1XfOHl7OexNZHkv07lsDd9+Rq4xAjo
ItieEdrCX+IGkebeUg/uyEuCAvC/h6H+d84/VRWHR7NIip1963LfYCpJP5jvey08
Z9riKvqVzdCCdkJAH2owRzJvq3HbHrXoGCwyMJ6rRAZmrBZ4v2H3HYV2dmT5D17M
3bNTpfEAbF6NoE55ZlzdLSlmV9RuxKlMuz+pODif4sRZMU1HufN2h/HGGGJrdVCa
sF+OcNXfOT7qP2gdFYoGP/is7gdwQpvpQxif1p/h0OZ1Zszju+1mLxBpIwYFq6k6
I8bEUZludZvkYei9eqPOYk4+mbUZtykmZXVViuNaLmXEPGAYRHKx1coOgjhJzHQh
EVx9FOEGA9y/Nm+YJOp9MB8tpdP7RWeiF4+mdHb0EMRc72kxvNp1ZLIVXi+HhX7c
8f53H6+Gmw7tjIjYOXWpOdUwh8EliDOV6sgHUPjmd7d1mAKRzqWERSoafN/DXmhw
BxxOy7/TISiKjS5/R2GFgPrAJseuOPCIErh3qSxY+lFljWTzdrIA9QerzCAG96Jr
KhuRedth4YMYaxtVQMLf7qo/hihLe533a1/5sVXpqBviQEwo20ey39haFYoKKu0x
mn/DzrYn4h8rYXrvzmf5Z8EeiycG2fGdalDp8NbYOxSHAl5urI9s5yucCSEPKP3I
4aT0/SxTCNN3rzBq9wnMdM6DdveoXYYCEbVYEpAjz07MtkIis5sKGKYW3tYPWVXT
AycdTvAGFLzwwbSb5pDzNtYTxSn8X/ALLLIEyLjEFkLBZT/2uF/Rk1CW/+LnWDTZ
08BE/lr6ZWaJyTbKokZAfTk+/XzKtGhdQ6sGg/vhURnYaBIR+/eZvGsQDG3w8TQu
NM5NF7FF6czjPbH77TmkqTUm0tE/ueTTcghPXHa2/fGYveaBzh5ZQVNm04onJQIN
RjPLyANkVM85yjq0QgZSU/DmInrw6WDc3iWqvL0i8AU4QK0VzMWkp/btRcegFpAo
QUPREiEE/LLOBC6ltZqMxSD6ghOTprqA9gbkZf0zLhapLT10ZRfDPZCWr+kdMKtA
h+RutwxDi50JoQXMPnxLUon1rhxjH6cC8nKIQ0sCxpXcpBoOHqH53FalCelm3Ow/
hHEvLpL+YfE0H2U7kU6PQtXgR7LobvQ1dePPNoS2V73Mc5M6ei7NcaRf7GVCIIos
8CM3aXgSzX835KlYf3rf1KPy2D/FO6nxxCsdWRTvqNCBc9jrGdVI+kWybUTPwq/I
7woLq57rJ/wNIQxCRdVwWrpBYtiqAdOt7CjCcA8c21ufbQVIk4E87IMiJv/z1ySy
vrkoJHB2jnX7fG2DAZMpFk2pcV4dawnII9v0FaVHI3dD0xDsheNPOM/UxKcwoA9q
z5dDjZyG24hgab2QVFil8g/M7SAIK9u+sNqMKDu9zCxPB2ppoWcPfZzdxqym7TZz
KRVPjQ6o3NBFcER5Ijflnpwrwbckg+wyXqomjtitoTIlgYsnNjkqSVACSgAEKGga
9xxcn02y70D3DmJTdi93n62rYGPSYzUJxDfO69m9qccBNPmcfP9n6+f7iExaKwL3
2WXYmylyCEGaEeQiAtU36f3VxRBsvvk4+hKVZF3ViEFR2qWHThLTp217QPwdCEIE
H4REgB8+NFhYIEu4SB2jM5IP5WpGSB5iz8MaM8WQCyDbHyN2x7w0yGgkiZcDDcg0
BAgvXYHCWHHhA2q2IjvCgE1DyTuPavnbyXm4iljXOC8VoaFlLEH+FC6JXSlFjBJE
5GIELuzlU4zAVWBzgOq9UbRUHJrqBAiQHX61bBwP7SG5/TlCYP0kWuC70hGE8nY8
mIswwTSPgFsFC2PM+lSB9F1AI0gtntJBnO96Bs8bwcQYyvFwTE9LLgrYNFlvM9RW
VAKtKJE2Oh8nocg3l5tc4or6Na83mUWiTC3Hn2PN4AvYVQF8WyvH0COQEwaYtWW7
2q49D4L+TaR5DmQFhj2xtM/AUfo2ktC/tdsUMtxRjK3dXvqRAfUXlWz7yqXswi2R
VJRQaVSELxHhgL75KRbx+Ghi8Rhz9B+RPdlInMLff1d9wg5ZI6tA+jz52Xt4cQJ3
4dLIm0xWsKCU5zxHuDBwQ+UDs/jH+B/0a71Yy8sTOVz8zMR2KvU+78nT3QmdfQMQ
MziqbnRsoUSAEXoR4sd29qaPWHjkIUerQS4IufdpZ6RtLGH/1dBiOMOt9ersjYRt
n0tE/TsC1xgSWiXGWN6VH9ndDsX6ww254F2ovxcT+brGqQM1FPMqhgkcD8yEUlib
YQSI9wR4qXHx1j3SvWdueW/eoxG7jnAKoxCkH389M79KYwEOvxxJwbZSibJQpkwA
iB+BFC6U2NoI7boXDuC7iU/rzrEryn7VdEE2CGsYMiho+8RDTtbCroUUGB0a/eMo
74KqBdLQGah5Piyt4+DWfj8kanrRc3aZldm4pp11GgRHSTkvXZ0/KHPzc/MEkslG
VhGXuc2YZFylzCKbCr4iYB5VDFYp/FV/TSTPYk0agmrjKltaSitkbQ+c24obQfgV
9RNA7wYCJG+OA27nwJx24sLXTL8hv4kCmORLfldRCxUyBy/c8SOA49B4rlxHjP6N
+OsPRFtoPH7+qDnjZjlZAtUbrA065oo9n2L526Ekmshk0VUJMo4MhxuXEkF8pZQ3
4TgU7ukp+0iuo5cdjyY44Z3QBajLuv2v3l4TJXhT9/vg6lfRqW+yRDjGj32qIRRy
Ak6xhsB15kvs5yWDeE/5Bg7UWc8/AlnE0ey76JkKHPJ5dlD5k2rfdOia2MyXvYVc
NDB3D6gYU3q8hRa7zmAuCQGhDHySW7o0z2baRzaEzVtJzcpW0JXd2DfqXtB/M0aE
4CAsAS6590gL0veHtir3BMkPmHov9aOk22jRvZ9fyppwRp2y7QNsB8f/H3hRW1Hx
+fJ07w3yOVLGoS9uK02ymx2x8jBuuza7+fhsxZ1IewUM5eAgt+cOcxvqble9d55a
K6ztlBiW804NakgImwMlqLpb/LZSD/75P/dyZQecggpVflgvNYdXNHAHG/+HRVgn
6hB7faPtqIoq+3dVxxv1eHTfVPQyOcCZWX2RiyLlFmhEDHp+oenyggpWbybjPFZ4
KdpIUY17MPwKdEpK/OqgbEejIzxyrQcAvdOrPCejCDLoOoHemjt89eoNtu+z7UOa
dyKZFtwfvzdSoLCaQDakScln74eozxBiNdSVLHBPoDuBMubb25BxtHu65ckidrb0
m/oPhnEdKCXRG4HXtGUh/N3mnr3B1wooyYd+xI2cbheozTL7kPfyaV2uwk7qip6a
dtkT4ZVW8Xm+TkAXF6WiNFKFvxR/ZZhD4Trx4DVwPrF5q5822C534ZxZEQ6B9xSo
iNT25tfyovovR41aU8hhJnuzOz7fkfYABnbP0VTsTcxSInXDy9aP/b9/9glBvid3
8H7l/QnNspviRmT8W/kxjXoU7RVgpf0A7rewQIvt9QUxJzS3Zhg54vQTWvDQKS5Q
1F/zlxPSzSorNdeQbm0cldGfHL7fg/xv91BXIs75Gf7/Vl7AJviJB5w5BoJS6uCw
6UTF7tFFYTYp6gBdx2xy+W/coVE6RgkgvMHtBFuWj/rSu/oDtCe6IYIfd++SX3nt
FM8Bvbm5ERuI2lyzK3z90b3KPf/KQs1cluZ5d1Z57J5Y9GcbJqmjQml8C5ILwqkD
s8zUzmF1NM1ptsRpZUmJPxgCYCMDUfGZsCNFpc7zoA6VoQIkqukNgvSIlmkxXQRB
IKxV0p3fjObcHks/bNDwq3JBS9vJ+3Cp7gZemd3//jDPRdo17Aw7CXXnaZs2fOMA
MS0Jzl2bImVKtvShD80qEl6pVYYzggWNtGe7oyrj/L0GqW7WoazmTtW3OgmkEGsN
hxpWrnS4/HsHPyNWRLgQZQhRlbF5AdfiNzvvQTUThJgwmTytb7F7cuh4E928wAC6
0Ok//ZopgrotBFRMNeg9AlZcyJKAxwNjwgoBSIHTDGoQz4ceB9E+JYjEanvE50Qf
cBFMt6LWYg3H4tBTEdEJBmlRqTCcOJLjIjhlOTh+o++2iQdUWRzCJYnitTGv0tf+
fICeD3z701egFCiEuNlY95vGsjIbDjG1VUl+RqiJaeZ+OpNOuTN5KHCbSs1w6zdK
P0f28mYLwrGzTf2+6gcNGwCUqwxe+yh5tV+Oeog+/xuOeQuR2WUHBJyVsGOIROZP
Ip4N5QmIPCPbtJ1cX9tLGtONFhuX2b/pY5QmQyHOofVqokkY6cy1ooCvXtk2NjMr
p2FKV7rDJoEI6d9ruF2UNnH51Edhuih6TVkrzJX5+nKZEuNtzLwFMlF3ftJo7ukk
gIAk+beSBUKgfTdFL/f6oPAYJgd5sO2BA68QWdzPQCNecwnL7GcQr+08Yj+Gd1kT
GxK1ZgZPtVewoeWNc5ALFjJHb57gz1rh9LmOv+d7oGYGZahhjSqfcqF47LnDLJvc
vFaSOPrs7xXrSFJzhefmlub6BumVHN+ilnPK+Dvqwt0dnCTn7QVErfgBl/vXHMaD
wf1FRxkrFs2popkoYL9OXcQRXoFbyVDJXS9EX/wTagUEMAKi2JrUZ4tonsj+yQ+G
4DEYBSta9q2OCF360pS6/WTs9xpqqcdPA4TUsaCcXYZNCJN2AO2GCjHEIBVWfKN4
jaXaEXwvha7uHOroBpeBpA7nDFTkAfAU1fhrEsr0ZDVIF4ZysfpHnqHYtVYz0r7Y
jfn1yiaFe4KjSLF5vT2Y5H0vY/+l961Hu3u4rpWOhH8ZSWaKu4PmDNGa5gEt62lk
CIuL1MHzM7Kbejbnrhi7H/isA1fxjCgQOG8swoIX4B/NAQn2pGFE7JNBwUNedOHm
D6Q4V/+xq4IyRC7v2EJ/BtmtGmglhQD2tYYR3rGl5oFXcaw0yYOUMdPIePhJGhBV
UBHlRRB50zPLCohIsDug4PPse7liDAwz/xzgGXsSC186/B4Eo98zOlxXTl1L18+S
jkIYNkmmpJNhksEVSl5xrNT/NBqYh88NvapAoxhDzi/UeD2pkVUnu8DsaY56yzn4
E9BpH0IGxM+DcE3qifLLqFTfImZx8p/WGuqeNose+wFCsNO/+pExBCY8GG+aaw3J
m+tc8MrBIkS2PF1QGZUmO8lSGcx9E/XcllBHVQJC9RIAwRxP2l9m4p39WxxKy58M
c/Ci5yTrPox7bMoGedvRP08XkAS80mtGprJjI5p3vpLLWz6QqUIXr3SykxP8M8aV
81h7R46ga1WeivHn9CFrxGtQWqhSBzcqIpHDGlUujZElc13PIQiKM5UJKFmme16w
rtsCFDlH0V8CxuXxNSJgOV0vAGFvaL0D34reN4hI7mepbwQTc7aKlLfkks9U2uVl
SOC3lI1LG4PJXqp7e4dXIoZJV90qZm4ZZ58Pw+jyDxOcAvWs9jb0vy2Z/jvDKQAq
Zh6LkSzaMOuDcwnpXeRqeF6LDcJV1mLo0NSP0pI7zIi9B7j4ddWYZnfs4CBUFZa9
xbYOKXjx2IsZQ70vYTUjrfyHVTRN6/3v5pClfBp5zxLLih7uQ8j4cnNAkrgJoeCv
YrjG2I155IyNyEvHY2yTC33HClPH4ExM/wCDVvHSwgxZnhIun62osRZi3tgZEkuT
WuOxhSXnBFMF1SuROhFT8mRSZhweVvAWiCV9fzx/dkIURzkac09MzmCyCvGctp88
47KwfQQ8PaHmRWBcQ+8XsNAEwotN2ToY9WnQPPzw6IHdPvRdgWTwoVCo8HagRsur
oMmxX6M0+4Pzf4puJR4VLqkLUTzF08vKQCs+SZb6dweJZiyCYE59UFZintc9CV4B
w25Wltf7preqZWTBBPkqTAvfbFBuVaNBrz6StezOBRgorbvF2qv+VJ582tTbimHy
gliJm07M3R8HrLTUGhaR4+5vXYgXy95HHlB1WmHDq9abXMw1YFKkZRjPJfJTCsDO
pA2DGTEGgFhql7ZYl8shCJM6pV2euCsn4JajU0QHCWOvjZwxuGj90P3mqTYNrgpD
HwgCjllr3c8JvXgp18wwWSsrYHt4gvHrbx1OVnkhP9Hl3fQ3EJQiyhS0hFsP03Lv
pOkWCc84WdaH0xx8uD8QFj43AzhDW8AutFWwpM9sjUczv2cTzA8K5YCaXVQRMtVw
39noJRRew8Z4HvoLm9A4UAARj0K28G9BqXfaHu86gQ5jFo6ga48RTu4GaleA1Sq7
CDQjqAeyIYX2HvZMrcNbvgSIEsCKFi5fxBzSD1LgFxpo54li6W8rosbyJZf2DP1r
3C+Zai9eY1DJJQFldNIqAknp2+NDohiJXPOuFNglQRM4yXUTzHxplPTHw/uqq6Xx
vTqgCVRyturKlAixKPif+yE9aqY6jQENRNwBb9oFrdI0rrPCBd4BhZw/LeJsK/gB
c9QkczXUYVgHuCKtHESUQpB4ACAFEuXAznW8f93y1RCqFXeFd7kpzibGprwogsJp
7tYQnrjxbtdFoVBSvxT98NVWQoBo79N2OWdfNMCcEYsfNokpOoDNVqPidOUbLsKD
SCMz4uP1gUMHrxdKrHGza6rbJOoXqsQVxHv4t9MNyhYWQ9N5dUI2HqQfpyP2U+uw
zPKPpL/tKh6yzqJgK+7V/lNb7GgmM3FH08OCmqcFaAjAkJlxjW1fuLW4fJCS3b2M
DpYeLddA5ATVwtigHMkfgn+iOPIaGzXQEnghxGKPpdLgmpUITPDpD5L1NBhMOaiz
5b1yemMrpleFH4v009cM9bQnvshIni0f7FCPmAwdZRve79vq7F/jRYU65ELnBuUK
pB11WpZI9HqzlVTGojVxitAXyQqs2nq23ZVLHZROWpg+4bQCx8AEDVX40sr9GrBD
F2Aj9u9C99W6/7bzz8qgnvoLLUVIEBVOEbl/AAhS1uOxsCQs9EPZSmRMNwNqg8cB
AtFzigi/Li6NBZ3aKzelV3d+H2Mn6Pys/YGflEYHmG+jzB6cOXmYjBtyCTtjWu44
WTVXEacIeaRqibXgSl7GR0CyOEkLll1n9DIqZaQ18u+ZFDDi1EJmR4PnTKbnoiqm
OVSWh76Tq358SQTxdcFYRxe116DWqmyPEf9FzOMSBmwz8muCiNhqweF5jKAOzipf
8uNy4Xz6k2b+ZS+/l3qLmik16zb+VSlZdihRvsNtfkNJs/Ml9l8af0r+7nsCH3Y3
lIoJDb2mwJGD8N9XlAu+mtI/+iK/RKn4m9I6gbVZi78BmK77axXkCDqwyOm5NQ24
E2NzHDf6zmFDPJg1KRMRBhGHEuoq4DruJle5MModmEiZS8ZgK7V0RNzRIFlHW9vu
b98u3pA8vXZ6HzUQEFkSjXoH2qBua/LlfTROmvcd8k7JTvqeGBDj1cwcJ9QaSFbD
IjPnDoZ9+ghvID9lbcvLUy+a/HVY92skfXj40YI1qhDnYAWf1+35WATKK/oWU/N8
zX/V8C2gaXQCgYZZxgiFwsBW7lbuV5kKvMZ+xU4SGfsWXi+6McQwhwdHXI57X66C
uGzN8/Onc64pO+q/111DwdbNHAQHAV+yrdUG51azA/ocy07n1++Y9O6kY6xyTQ4J
E+Po2ITmI6UwnCY/wayCuzO4NsnF52+/WD3N1XOopMnWKqx/qheL4N+2UoOD6XUq
Nb3zlKj3+eW/GV85+Ei4NPQAqAiKuOhS8vvWrE+HuFyXQ6OA8fUZTi560PvxSATl
noeGJp6FhPVS0bV0K+mDM7xxYkwFLq/1VrkYZvm1cEJrLUqXYLAQymDTQoagEj/S
RqlutPUmrrb1XDQyHQ9voA4W/yu+EqjxmUHd/6IscZV8K7MHsgOIS4WMWV1JH+YS
rSL7JfmRGZhMLzc+bVdSU4WgnwakuAxUp7EEDvmwFb1fVhawnl7BkheNyQHV3YFV
wMTnCcmdHRdP8Xxg/I9rFBhbL1Xjrh4975al2+ESK/3uxlQEzSBNGxzLsHvXHMCZ
5R0rpklg+k1EX/W3v9pprLu/yAzviPM2vko8fHyqmypnGmwT0dQYtf0ATnLOK3ib
vkCZ7qo92QMn1WozkBVXznJGfni/+UCFKGmlOcYMuXrlfpzKFBtABgYDoLR7voJx
EbAPmfsFbwvrDvskt254getMci/bqKTGBW/j1No5MWnTV4aMIzxHwfNEmdA1g5c2
wBLzVP4ERvlbB/Qk0nMP9ESgGb0h4YMYNk/UNYW42XnNj2i2QVLnr5CLtQOlZeLj
RVTwx25NldZWLhSD+DHL9Fuq4b8LIiaK8LZamUuLUnLhm4F169lMAxcnMGyw0mzG
HpAQTZMyu8wtzxYhsqY4vWVFgiIAmQMmY4kMrbJfPGiZqqBmRyl3bE/NNqev9GwF
gKSTqZGn+4Hgxga4IRf8xzvnuRUTiJKJpaYrXknuyCkzKq/ff+Tjm32nTUGKkOzb
Qzo2Udc4IBUV3i9A1usR0GJIOOJD8A76w/3z1G2lQuMXMqbkoDT3UhnObNNb15ut
Nr/yUT3FveS5pxz+EcOshFjlcNh1sHd9Y4QvZBLUjL8BblZ4b99rDLUDaHam5WGg
YuxW1EbRIfEG2ljtL7UjFM1REdajakLpyvXYZwEDkj9LRUimrUOzOYztQuT5N9se
7h5+V49kKHnkaRXwGr9OM36NCZEMeOIKeicASJp9Oy/0eOAtoOLHPehk3gugCL85
t340vtxlEalKXyCiupanlvScrGXpouncj4N31306NZLMEEczmiBgz4XLykcF64FK
MXRheGr99AxOIeW4yEG4FHX/IXuS3aILGmhTkRGClXrU4KseM29r17iQ3YedOMnJ
JEVoAYbD7TlP0wQ9gwYt75SWzJRH1cIYoc0SiJLaWNUrUgH0oqY7pFWuZudGxXgC
+TS3uL+4Et5i/VXf3N+VquhhACxqQXykO+/I3Hp2mX61+h3nDes84nGscbPje4qH
XHc6dyOeRHqZY+4r3Qd9gyuVywakjTo75H0ap7ZIJMhk6eULYEuDa7g1SGx6suaG
/B6QaRXH9r++7i1ffDeGsZ3RzoejrHT2oL0Eoy1acnMbYcPJi4oNeHD3aQCa2jcY
iRcjU/Y1atQIdl4tNwsNtp3LDUwB5QtgfoCZmFaPIof/KtJwf7GYclZU7sR2PwHh
3soGbUuSTLMpQ0ce+ys+UKNNyBNMCjiwe9DGox33EaLpJFinmdNWN0fMyBVuSopd
4LEwiJHD5ewZpP8T1sxHvACplqUUWPbF/sygxzh5RikVT+mS5a1lvPm5cQFPd7v3
C4TqwO00gfk+kYiNmZWJS8wEZgGlR37LNex83xKJtculWBFaCikvSYmgJdrJyYeQ
NKVC6dPvo09gRSlcrZr/vNcgRCkirdi/KFkiLaa6X9Yv+B1M03IS0qz53+u/omfQ
q/9x40N2bRyNle/pGskwbHWFcbe4JYdKwLel6fc33XgmkvD9nU4nI+D1cAn6CpL+
7mTBMUeFk2TVpvegyWT1Twc56Utsh/NLkno5e8zxaW9L+UUn9dt+FVUffAgt6nFe
vTNqzpL5d1ATMZz3XrAMTmTzfIlWhBRgME3b7QtXy52tUFDJY8hQcMkiTsb36Riy
0xULQodUmx28Cy0cSeG4bHdq0VLMGluM3c4KJgtbIukysWIuJmGtYlqqzXxrJASi
eDSv0OU8XNuZBz2sdPmgs745U5mVr2kI2pRB5VPz9cTxRz2AiHiEw+SiyIk9TZD6
eP02HGopY+8cv96eNA4pm5CR6RHviNQ8qyaDmbxV4P+XoAaeAGmzIgL8UpEoChK8
ytt1cAqz8A8cFMjbm867QtQRpCroQHjmPpxFXjjVGkkyA4igLk+hd5FAfepI+d+H
QEV1H1NoOtLr3qHXBy83oqOTUDG6JpbVG8nL/OwuMe7rsDxjI7fgPJguHxJ3GBIP
lcmBaVGz/LqbKk2wwhpiNi3QQd+8BCvOjT9/hpOXRBDHzaNZDhSO3jL0VjULTaWz
8JQFsi/blS0LVeNXEyAn73V8eSoLjMrv8agNMVtUXWMSWpMde8BfEV8opOiFipwI
K+25DQo/k2xGKYlHZos4C2Dhytr9UJ/UuFeYXJQzZwo13omG2bxe/pWb2VbQzZz5
7EYiTfJkD5KOy8LdwDUb4DUe7yK3IRCJ8wwAriygW+idYqNZm6v13eZrP49VTefG
dplnAbCENLyugvN0Eah1jzguhWt0yVg+FslVmaQNUWsjVyvucxP5x1LKuW5lgzCW
ZjVljtWTrfQqJHuoC/xTA+SxPyN/uHzGd4enyadiYAQttaErrzgml+lC35cE1T8K
wMPMXZcaKoOa+rcRTZxFPIbVueI9njfhEAVcf7hHJ78VAnpo7Q10OEZrYSTDVP/Q
LpvvsLeq5dxrywGnwlklKNltbOdqAim1azbPUG0dKI1qsw+OjRLXkBQqfo7lscrO
zAyQXErJISchDffKZOkLRMs97ngLXKncwyTUbNnPD6QLagb8oAcJq3wvBOEUBMr0
91Tksix8QYC/bcoktB9UAJVs2Q/2JrwHoqANwG5EGfRFsLBEubGpUb2rtNP2cZj5
9jP93//3C5LgHmFCcJccO3JfJ2AM2KeZQjgUiSZTiiyLjM1jrX3YfLCmOdee4eG4
/Q1P1HEllvOLuXmmfFEoo1MYdiWDcPxq0IVAF3shY3JjPnCrmIRPOgDgzQfIA4mq
we3f3sBWFydmt81n1f54GwzSbi5w8uhtLryk6ohSqZae5odt9I0VKt3pQoJGYojJ
NrXSaulGg3EjNzhLaoKIgMXfSHJGN4go4fODAXQawXRm6SwGecSimx899/YQAaBC
pa2bFEz1y0R192XvZY49DXLkNyS6qYlHId0EYnbo66oCDthONdis37OMGNUageNO
NXX7U9FckrI6gpdfxJLaynhRWr+I0eTUO7hPgwcl6Mrg0N/xMtrV5z5oFmNdkrmt
YBxMpULut1FFrleMlt2PLEC24M91EE0/LfHMsr9vDEuBGfIiMK6jQvZdZwv5HmC2
eHvP/SICj2ySYg51GBZK16CF2AqeRMNnCjZo0cU2F+lKFGsVTHAAv9k1ur0eKDqJ
5euwmIiRStzlYjdw8yO+Y73eFBpdbmebAOkrs6RNW4cm2p0ZsWRAbwsCEY8ZDn5m
rBdbZu7pX7FTNddCxHX+v/oLuMUFTpTmXDX+7zd9EkQo+q98C1VEosa4UCR/T8aW
9cUqtp7mBW9LwbSVKxzK3J33e3Qf6PPtqv2l1V3H4PnHlPSmSO6dLrWAyVktnyUI
bYJ0XvI6s2atQIaJKHAjeRmCvAjhwLunEV1faJqp+lDYSjIeue4RDZ+gPXOMcwtq
jmUlpzeKBNtgioq7UrDx3vrU49QbX9f+s1OrAE9kFDt/LFcQvt4e2Be39Y1pTt1L
t1orO6CRzsAKyI078ynu55pNDG9MXxHxAjwwzRk7pTZFL5oxDeTRNDUcuidjvePP
j42mIEIfMq00NqNbBVks2J1KHeORXsRym6TZduYrV8KHNOtqLcAEr3+/FbT8iaE0
nJZO+ZmankdABfNGNIVv8gsfBKEAuaeJ2hhdYghssEQQvJfWw690WIMfabtPwY4k
aTTfzxaLsPFI/X4oInq8ww8EugLU6LfbptTpY5cjNuW8P9F9gZEzJCnjmQvINae3
/xMhY5xf1XPpKOF04DNqM5sbAHH9Zu+fIOLiiiA5pzjno1L5uxJSwdJKLP0X41yV
PNMuBdhesolcUvSCiXPa8lF3olkv1p1IKqQOmCWCSJOo6VkTtpAmCXphHr0XKkvl
s5ncf4mbaKsbaQ7I+MsObkONH+o39FBwh5oaJu/7HzWRDPJ2RpBkDUV7S5YDFWCt
uJGNPHt09561+KC0acLXUlitkGYASPssLmUQycTRmmrao/v//AGeBBxSQWOKPklW
IIYZ0Fp/KPij+LvDAhRsr5O6b8wxW9FV0pjR7bx+l5lympZB4xOcw8BZ9eSenD/4
7TCpBhEIbmekrlyo0ZjYoL8QYs0yTIY5n0shXNV7Yrp4UdjEIMaeN3DmFemLF5ne
+9+TW4+/C2VXt9lsjLUuRvj5z0peeIW66m8Qh6qbXKX88rTHAt8m14Y8y8U6GV/D
Rap/oUoK5p7LddQ1sgu/Ic1XwCrueS5dwrGn6med2OArCaXMnMV1e+++im0LOy/A
idjhi+NzcWkq7/VAJExpNpmVejKb1xPmxEkspevvi00Zv0n+X6eHBe3pv0wwT3ha
Tt2GEhnMoQ01eTGgMvRGVUTr64D3jr797WeXB2eED2+NfilpwqCCZFJYPFimafAn
ULvU1vGLZ+IP5LY2nbclllbKgVR0teIL+T2bgwFR/VlDeJTqenfs0gwpSFNX7WSq
XZPnQtEH5lhtUHnj9ikkaJzpLsOsYOj8JvUJlaERnxKkDgLWJx0hXJh65HwRYzxX
qfIYF7QgvoVbSXO/B3I0rCmShKPpcz1q4TNxlEZJ7mFCXhI/nbvuxTkv2Ujpcy+t
cOmlOPyKbUqeE4afkDWiORXC2wf78JwbxMsFKay6b0CILaraaP5RTxuDPpXToXC9
aAKbjyPv7TNeYdYpXYjYLKJLCyAIx6fiGxozToiBQgYxYGT+XI4CWlxIZFRsfapW
Dqi7/VeKbiZiChoaTersyU5cjK4jhGyEUzS97Ux1SkVjNuhEhZbOs+JnUOv6yUbw
6ia/mAKrGNuAbl2GOXHVnDaiaCtG1XdTCtaYmJOH2F3faJIP1iBo7+FMIe8htgop
CTo73TbyakPM50Kp2Jzc3LQGfff2Hp98/m9yzllmEqGfCXoc5jOchQq31kEkCHoT
raOZQp2dB5jUCxtAJTQmnNLrn792MCINcyLpcy3zNkrZPI0/7qTczTfFYobpjVZJ
jXCOdCnlDJH8wEmLwaKx1+ZSzq1NBe1nrHMO03FW88u9ge3PIFOVs0XFI3naVqnE
VyrhLzgJSLFe/vqkItYUtdrpyEa4Yf0Cu54DgaUo6pyYTHDqn4sGoPa0kckZR2Mu
tosn44J2TJ2g17F5zTm7Tqt5jP0fvEbeN/GSJZhbMeXyiViaHtXJlDzSHfE/6/ih
1QZj+l2MggCjH9J4acpqzt90suSETyxTzJ4Np/YQSgm8DvsHWnNXd2f7P/jxyw2v
YfOgpy7EUqimNbEQKH7YXzQ09w+6CPIIauIRRuOKtmOy/vBlgVU4pZfKPKvHDct1
9DrQLXdyALIRbMxboBdjFPQo4DDGVii7dQPMnsKgQrTaAGyRSW0YuZGVLJ1KWi36
W7Yzrix3sh9yE3scXUuZWb9lFaOlDhDUD95wQHGVuLJELXyUXz/tMhuXyReyd5NV
rdiPtLK+V8vY/VUbb0LaS06EXCMJEtX+2I1XY1w+i35gmtrjyCSssE8KCKZuWDRg
cIIzjdemUji905XPdyAJtKbGzDA54MyziNlT4o+B0paYS9DVGSmzNm08+g+YfDeh
HVoaMVeq7DghpWkWXFkoBA96Gs7Vh1X9rQoLvsRELlCb2VQC/rOonWXgC8+398AA
iROxZ5bvTD/cypfaEPyAbZU5cjTPiDSDSDXDoEPrvC17aswNidtE+Vb2LTx/yjjV
d7TOAikjs4XAUBtGmjGSQLZtUVsT5ecsoNpn5XH5Mho1+Sdf85TZGJS9+qu89tXX
E95wt7VzwQvPrqBxLz1T08aQSPDtPehQUZkTjgPGaOeBQBFaxi8MpVFGdEBqMIfY
VqjBcapjLaHwzNrfecsz+vOQtP7NKilDt2d1MqpLmbHnPyNJgfqActOpmTFIPh8X
55CwUcf0DO4huSCQe13IDSMArmfsXjYQh6SDIPpQiMxmAzhSFKWtV4qn2tcmBrgy
NeBHygzZ/HYnvLmI6146BbD/65MT36DMZGZCwACZPNIwZaiqi6peA3ITof8z/d/x
7nnNL98Cv1Imd4bK1nCox5Eypa/4HnEFSj2OwiQnq17pwhQXBsTTu6Sp6q7jYq8r
y3e8YON3OoQdDkMEcDpwQJewY50CCJid+EZHjEvYYp2aNFjyl03UCXKLpEgoWGx0
5WYz4QxRgYX/nnsctJQ29Wph5ajujPsOfBDATcGPHaBbYdh1yyg3Qg/n8By+XCgO
fIiAU4t00UqPxuA5J1GzcrTdGL1LovHHqePdpgJJXLQJvE9J+6DyUH99xBkGJ/7K
1viJo6d2zz/ANpK45dQdNfAyhVcPMx413XBlSXnxlIha5BgxZEaLsoikDt+kai5+
7fCW8Ffu74l/UN/ALOHRmYe82XoMoNoT6a30SL+R93YpxirSEkS94JmMFZzwGvId
S5xvb0Xv+GGe9iygNhaJdMoyb3/CwCp2HCEBj4ipdzj1V39lK5l8fhC60k/HLbBM
8u71bxZKSp5tyhDXJiOuVP3jD/SvStI9DVI1hz9nsXUV1bU8/2/f/qfPxRCwn643
fi3Z3e8RWsk6iqtqpqF05RX5o226Jpv3KF2TjIu+A1Bw/I9/7fsqVz7RKbNUslHg
4rOPDXPuC9lFalvLooUBkZvNJO+OWkhfutrv+6GsHWr56lf+whm5QBGpG662OYCD
3FgTcRAYBlcjtBRJeTRYGeHHd5GJHqGOX++vCnsDlVtkrb9cEOjWSLVAYheApFp2
RrfZahk6WI02Yb7mR6GEf/ylXrgS6xqGayihot4TC/I55wWWVdy+u7/qSSaQO2OO
DpnmJw23/XfvMzIMZPf3e85QRpMLr3AaS0sMh+/gyfuYE+GOthS5Sj7DpbjrsQxd
sT2SmgwDzrCc05g+3K4gsbfMLVSNNTP7cc3j7/7RmWOH1qcORM+aWdJq+NjxspZa
+UM9Wyq0ePXSuokURKTLIwN1AW3DZheYc7N93SyHnXPPNUxfBCzu9a1IfgvdB7Dj
UTOLZf/yfAZJQyzmISdDaelgMFCdOKFtC+ijlpVkNVvmJDna1aDqaxt9+1nO8VCH
0Ab9/f+v7va2UuGQQgm2PMCgTk/Ee9X6ivYnH2ptsp7vA1Rj3jlO20H0gLgyxFSe
MusPlc/WapaXgMqqFCMF1cTnODs+O+5Rn9EWd4IvN5WpYHbb3BmztrYRX0H6RSxF
tiwNLKq5h/D6fEtfVUM204smvmBUxHI+iCaux/6FCjTRrG+UBhuLI6LMrm0ZI3jd
cyOy2xQS6Sh5GC+RJpi0KH/Nw5vGBNrTCqNwNxSM1FWF4BqbfRiqNVAdLisoUNN4
KMPLfGCqUMofCwz/90lnZHn7MQmeE2HfdL7eafm1zIeuSM/tP2ko9+icXQLQWmA+
vpD96cMOcoUZT2SyQ09UgWwFFdhbeVpbMlBKL9wckAsNtrCv2+oi5EJ5P0YJA3E5
nGenDMz7SGYV+uzT8316RnaEwQvw6YKu7IpMDppJWn0WLaVDBA72K8llx5TPIfdk
aOjD6W+aU2NWcUdJQx8z/jggXe+OxCXBzeGTD9H35o42etNRpHwFu+LQPHpuBeqY
5bn3uD29RTiZ02VAnIcxrYpjsSS/ezKxs7HeQF5APAcJOYWLOGPd97uTc4lqTKWO
VS8vXUWDOvSYY6bfuCsw90qF+DzvHCd9X1KNs9pd6ahccwQs6OnFeGWGdFZXlz2q
yDsqG8OWIHysvl03aAJtJwC91mh60SzrqdMfZQ5n09EB4jbMl8JQHSTtW6uFkWt8
NHX7Xnh9AIUPre9c+mSkdHh9KWajwn4AHUS8U1Z8WeXo5f/oEDbiy11Fk+50ybgC
3OdrzKQJpG2k5R3q3q7ORs0HcJX9+wfSnlyEeMQZAt+P1xW6T0o5kaeSzeEUXKEC
gYc726U0iyL6/g0uUW7KLuoJAPYlB2Bk3p2IocVfTwcAozdebsMcJbFqvccmxPR8
T/jAUUokqX0Dyy0H4QvsNG4JEf46L4FCVeSKvjeA+xVugKbAL1XN6BrXfe8ajcxq
GFzkAeujed2mx9edW5676J+70eo6DXf3Ha4ANDQvGz+4fMMF7PXfoolw3x0XICgt
oYX0AK/rrMffjONujODN+2NHkEYaeylaa8HJCuM9r7pdd8RDGxFZw5HWIgpenysn
o8aEG/JT+7ke+5CxqENeEEvIVbjLcwQv1SM3kOLe+fn/ZS6VkY8zoNMriX1Xb/Cm
Gyn6bzKvpadm5LSdiG99tiWiIhkcFvZSf5NhIMQJzIyPzP7zq81HVLSsRfr5C8ch
23M4L1mgQ/lU+J8TyPB+2krfYf8KeepgIiQrCfSqDJkHGP5EzfjfVkfZ030pavCE
HKawuyacXcCeOgV4Bl/KN7iev1Sm3kOH8Di2plxLtZcIdMa1JrrbTOsAAYt2Ntrn
U5MTX5R7Cfh7RMDEKrSI6wnX/wkjJA+XNG/xmbusD5HT8sRmEA5R+vvJfOpltoTy
TXdrx3qd6a/Qk7cumvTIV1OhyOC79VmocIqn6PsJBlFx33WC/n3/J3JMIj6uQUbL
jFDZ2Lfh5rdDfA2fjkzK9mrWZy5Gpb9zwEVWWFbkGlhQ31PxOGGgHRcG2QxgJi23
vIflI1ozVF8Kgkvt+GAuQg1PTRB5tGHCQ9NjIY4ggRyeJX6yRzMgaEcfxiY0UQ1t
0kZ+xLpoVl6Umb2N6aS8cz4sBtnHA57hnXQFox4GdBjfvci7zPP90dOjDrZpseXA
hPT+kta8cTMQjDJPsxt8hzcHnCk+Iek6SvjSnFJvrj5riwz2anpc03sXEwqJhPIh
5IltQEjlOyEineOykBWtn/NLdt769Pvpj3RRRwnROH6DGe+5QHtXxss5mDhQV90r
8YQNuOvPrCKAItpxAidVwTCvqZkzbyQgOR9csK9PjQVJC4n56H1eY+yjmUy8p3qa
PubnCdF4XHC+CWIFl0P73jLb83SsLdRv7+wccKgVpV7hvnTxTuYfgU2RM1j9wycb
MMk/FepCEl9jc2t0mVgaF0xAO3vWidPLkMp1ncjXw34JDq7gewNcP5Ui+G9UVJ0X
Diueam3vgoVQzeU9sMv1Vn6XqwwJlqb+xfn881GKvH0TyqxrSbh1FWl/Pvl/iCqz
4lLjPrFH5HOGR8cdY+Eeb/9XWnUNu7g7V0N6GOjAA5Ki3t9U/SZXRbFcgxazALVg
B4Tl3zEWnjNFmNvF4I4WOzTbLMlv3DSXITttscdfY6NXq32KjzAJ6nWd2uuguQ0v
FmaL/PPw2fu2nwUfxubj1f28CE3lk0qiU73y8vnPtlh6vmIZb4QFb5cs08WbZQ7P
gzkyDxSMs4obGNieplhQE5TjzTBHsYQ4fjfL8+tq0WCBcNohUEoXH+hCKqZRLz5+
NDfhbLg3QEooO+MRm8knDiwvHB65x78wS2c5cTEPqnl2I+Rwryjxz6ZMPcAxlKsC
h1Cst9+rsw0doekwvr0eEyeYpcDO60PXBfZ6gPOOwqTfBl6W35f+VzxT4XekPaCn
WxOXDVSyJqy2WwX063WECf6xRSwFqCDL4614JCyeBIbfUGFlzlXHPPHFHz/cod5o
30nSJlFB5RWbWK2p3JLUwVcqMBgGwRsKaOCr02o4nYseLUm8vP9w6i/+SgQj69NU
geI7g2ZF+qkDGgJTAkh3tS9S3jO6PN7lhpCyQoL/muCw7uj0ltuByR8Ia+rfTJYQ
RweL3qtl3hiIQnP6SLG6WSprKIA0esArIzeYLXyKeS+U6wu/va30NtMznFGabBdo
s9aUbfGAvj+Eo3M2ROPeA6v7E6w+1aPx6n70FFBVy1535De7X1pe9Nw/ZJp/9Dci
biF+xenlqwmvY+2ZyJog1RXU3xpC8wpyNzzTEBv09skIgcGwzjnBwQifxl9Ebkp1
dqZcjA+DZF59vEhXNDh4A2uXRp+2FINkZPYx8OtVrq+j2oWqEq5ug66zDEw1kaAH
iFnE8c+xGCyXee9laR+LPOWt280r/qyyOqgqOLeORsYUo/CwrkyUBIKzXLNRXI23
CQKDJZcYJl1/8uEekWsWnVsnv8gjAMwhdW/PGGGIL3TUgUYAzMsDO1TCxldTG/f4
bPELfF4G/0phyOj8aj2bk7GkHYS7+T4UO6UWhoePl+Lc4DE0szomIbCM8O9Du3xV
i5kDYsvAE1/8YLoSAgfb7Ek2zzDp0aXYBcNV430s6eSPPZ9wE5M8Remqia/jYaXF
u3tbovS/OT5EX+omIpzyeQXj5tjZNjWAaqnXAywnr8+3MS3xNaSaKx7eDplWPJ/0
ZWu+Y67uhEySxg/aKVYNzOnW6NBytIwAc5yAcr3jueipq3pZTeVcZrkqlA4IMfVL
VhbQAOpp7JAd8/74vnCajOkv4lItpyj8mXt/V0KFKKr6Y6Be0TUm9wjha7qSDZXs
BTu76eU2nZ4UVWCM+c4DLSab5riAgT101c8fv4XP/Iz0WcR/Wze1XLvh6xAhPALV
x8fnBzr1PTV6ygRAHYTHenoCqa2rpWEVkTBxBs0C20rTyWyONe/d/uIJd+cAw7c2
t7oIvr0WSCGVfxNCouydok/d1aPw9x6zdMxUC+jLpr6k492PfSKpBLfwJR2/4KBw
M4iCicSowgqIx6R1wNwlxFS5l+2cVAS28nvly4nhkiRpkRldlYR3N89Yg8FsVTmU
yHEIPbcik/ww2r5lAARN/TBTIi6qjExVgqjOhtZ+hyFCZ8xNSN9kCVGcPTNWd9wM
DQKnb6wkTz4wzpCMtb3eIZJaYiGAnmtvIo7pJ8mgEqJgGz3kL0hKaHWkB8lXei3A
eWrpGZAMA/0czh8373jNM4mL8/kHqCjC4gCvaYTZWsku2ePUm8PpOFY99FJAkXFl
7+k6Q4O8mqcMS8gSeWZ402sXfHoYkx7qCR2uFr3EJPooM5UF+Dcvueix5aPooQZJ
+Fctg7rgRGVnKt71UUZw+DGnaPDM96r7zYf6V3PRlkr3rtCgJN3LFLJAIbqBKbBb
u7vzg8mBgX9GJ2LiGZf0Grd/ZM48OdRD8k8toPEGyKaKESANWFU70vuvg3lskD+P
W/JRIjn3PTtw9VWi+acVeFa0jkkff8saVAVk8oW2x9rqrf0ubA1mjVLJN4Q3Hu2T
l/32yRS9Tnh+H7y0/rruxCdvYsmnNkrS5LfJKD2hujMa3+sF4MB90sbyJDHY5vna
7c6drN0r7fA7hHOtFGWhmJ7mlbg07QUHv8U26d0guNEmHgWktOO1t1U7WuAMML4J
mGU4WLUROgX4yMDKCWW+kdx5T32ET2uU6P2U/IUk1lCsPjVJB/aeFvzxmc+QT9vq
yXrf3FgUhPlF8SEcYHYVWunOWdaEmEvRty0jLVRyPOHxf92T3Tzbf/mC9fJa0yqh
LvKd0PdoOdBRXIbVakS8KHG5D5RUrWdmzH3zUpHzkGunMthhN3Agg9WfT7D18fAx
s2ccwfVUyLADXaL7ZkP4iCUJ8T+EIyZW7FW2iFNrx3vv7jYvUq+fcE+O2yAhLQDg
NjvJVIroDie+CpCrl4AXm9SPbFwzluKWbWWV7EHfErUNEsqJKAlfx1NAsr2L2flc
H03SJXPpO8HrjV86mkk3YXiR86VzTrwG+rmm3QCx6NDKyKsjOGYhqtyI3pTCgKGq
D21Hodfw8wvBTrpT3azKuDJgXGl5gMMx3BsYCdNYrENwDo59Bxo0uyxUldi9LgE7
sB+tqZzvwVkco+yN1k6ce8H/g1w4zQCxHmTs7pvXghxXtTN10u6zwwC1LQmSJssF
DyI0ZlOTq1kjPaBYZAwNkTghAMTkXTJikUL16s9zSWogSyBFd+nUR6T1v7R7WxOM
jnaHDbbFCUisJuH1KSafPlGyNOgykX0YBXhXxfhPtq4PYl6RNT57iGx7llZNbWGV
lFj3SzNi1Ov2R0ek6uqKTergZ4TJEf/UePacOsM3MeFh94kcyc9OZiAxHilb864Z
GMrIB9464y3stVNM3tYWZsolTiWApQD6l1P2sKW5jCb3XrMqSww1AuIZ9pw/qxjE
MuEIt2923XPnQt6sBqLE9PeLnYkGohbTD+5IonSouyic8IFO07F80lUsTtLzoCCS
fBhr+w4NSyA9UrZQXf8/XqEAF2vbsTLsavOHpJec9RYohNuOnsmN4vyXT9MZjlLY
Lt27p8tYTZtswrLuFyo3gDD5wV5mPNWAcZ8OYZVCwV/WBXpPDiTbbqphzbV6yLX6
63X60aJk5eA0hLJGm7f21YKdt4BcS8luLia2hFpHrrNg+Udu5FjVdkfBMlK0vogI
ZlVs4VrgjAgsYR0h/CdDvKVOR3P7XVwj84mRLV0gh7dUSv660KM8PjnhgqqQtSGJ
5xEt6VlYwfXfpUQswvgvf+T/S5fvJlvQ+OkxDniIbgXIU3tHEegv5MA+5+Uh95WR
IcxgjZ08zdUAUR9KpdUors66rJJMow/2dnTvWSmEU/1USwBd/sW/hlDuL8Iap1hR
APJRhwnrFwpQL97cp8KHAH2T68c2ECO8/HmB1X2HjTAn6oCqbPQx7QIlzDuLrZbe
6n6hmhB6kw+i3VVugte16u8g8dPYE4F+33BJMmf1aInMEqFepWzdQxAtLpR42sSf
1CRcTAN4C57xVpMlTPWfYF5/9edFpZ1O1YYxOOfvcckgr4JV+ns+yNVtaq/4X1Zl
9/wmPv6pmQbstGbsVyjvmKv59hK/IUqK91CcmzYhYvPrKZuuJ0V0de3W52vUe+z9
lsU5TQNzwZFpRq1JKkh6M7IrRMKWOv6Vl4F/GNudCruj589F8evqtNeJwT9QPWRZ
6uJGijczvb6rHXKc/bodQABoixRwWz8KyFlY0xkJfAMtPMPc93Lq3iPgpusM1CO3
9B4TLjvkH06uHodUkIwcRMPHEsokQ8yVZhbrLR7nMTY3tgVGeIXGCXZyQsWaepsw
Cb3Q409pY/+hB7hGPPEj1qTlWP8LIJw3EwpbVTtqf5UFdwBB2hV0NRh2EQbddUaM
UAWkf0luJak6o5jRQPHo5PDLzb5yUUzvRt3Uwc4SdZNdZJhD1qdjiKg4+T1ecRHJ
OfKh2KjxFH9tme9GaOML3cciycb87EwT9JyoGQWF0mzdXc8L4odkSMGGCD620JJH
SJra+z85PAhxaBdC4lDbOkZrEQuNr0R1Qr7MSgpSIiP3k2CRh9NzFdZ0Hsejpi7M
R1YbuhVbpNe5EZrEVXRuekaetf4VWdx6DyoBRhUG0PINA9KKnbqH+mUrOtvU0sgn
2QamFNuOX1GZtyJFqMV8QL0APM8MlIhlkERy83w1uT0q8j3N/abE3bmEnTtiX7FX
mVSrwLJcSFGiQBSV7zZDP+PzgkzePvqnjAW0YurNP9mampZwruv9If1gndJ/ACzF
+IDnbm1PClN1l08r3NNQJ8cEMGOlYRn7AcIYPZsc6DzMXSjF/1Eea54D2/vJyYxk
xy5CohN/fUmEr3EA7X7amJs8V1NUDywYdb4NFWd98ePTRxmDxLsRcf42ieW7H1jP
rgKVMpzJip51QTOp8lFSd4H4rarf3+4P4Yqc9M54DKD8LP1wYjuCL+JCp+nsWOoE
j3mwvY0lh+EQe/t6yCY0VrgcAP0rTXqk6szff/OKFkSMcgS3gHRfrizeDKHh6PtL
UD79KdCjMp201L/KomC8DbqTk/qxtvyi7BFjSX7p4NCn4ideoc9pNOLkpUTqxyRk
jAxb4OWgAa9/W4ZCsJDf+eWXNUEB4iqDB6o0mrNk7GaLvpTl4PuTLXujxiVPwa1M
3b7jklUZZWbTi335O4H4mW40gus6dGUTv2Ihz0eKPupcASniHd37bSaHk5YdJb3t
UdeCEqnOOdV2GpyJEv1S6cU/MbBZSaRbBpvbAbLOx3hbHUxXRu8jIJyd0CpTfZHq
MwZO4kru8RxtSPAwRGaMxIyhV0W7jL5mrS81WhLynqcRHV+5RNVlfnu7cl5kDLiS
FP2XyUTpHO+jbnKWrDriuvNTyppc5nyayYenB3f1oJidF8k1x1ib0qo5vPWM72qj
1R+vcpe3pU6V7NBgqzVhXY+WYX+V9RB3yxRlQfmoQNdj4Sk2jQgMQMXq/ygPhgCU
yPHl7js7hvtAFUPM5H5qfV2wMSRQOZ9OViB/gF/I1CK5Qmcp9IZW4Vce8km4kqTb
dR7eilNkrb3TCpb09UYnEGjmrGmdb7A41D1vdacQbtzIfGftrEkozDt2sjS84/IY
wWBYF9J6lcFQNcGceBnzGFrwx7EZbW0SsK5Wm115M9hOvy1oDrWqTgW39usSpRkd
VXYhY0lqIiHq9nwxwvuiaR+UVRZJ/ty3u9Kv8SlLOH1TQIykg3AvMmilmGq/lnWp
1Q0rCmxquZH1s23f2jg1q9e5oDi1QKehrbpNwPX+APwzc8cm5sfo/YsZwSSuwt1p
kfIU3JpLstTueYeeLWWLMmkCHnuFaPWEEV7+Z2BCWAs+rP57uu4hmQSf6Cb9B/0b
Ovk1dwwQaCzbqWogcZnSDQCMwykAsySrHRb0a2x1tovPqZe6FBIzs/KFzgskVjvI
G3hAkGe8CqHc5Uu6I3VXLF4sSj8wP3xU+iCj2y8L716oqgpahIATZDUurSJgeYFG
v2PZVT1dcJCq6n6BLA7U2sEau5aJxJCskjUcrW17ZyDAgEmaC657feJuUqjeTFXV
Y6SxQSt+sGdnGENxVZmFg8wi1GgzoR3v78ONRxkkPV6B5K8T+We9qCYej4l14Npw
B54q3BBY/66NyvJf1KvCXVCnHpj56ZOgvDsP382wXPWP5ErosViIKnsFnVl6K/sV
2wDfmqKfnkKmn17fVqsQWlp7DTOBj803ewQybZjlZu2QOXrqVzbAn+ThICd6I9ln
o2m5i9KeYRe4ZXd7E+hpOQo4v91zl5Mxed7tHTbi0MjoFQHNt+4qQYOrmdtuN9F1
/jdiNpTAEqqj6b79uiEZcoq1ZH4IOcWFtxHGXcIKtkM471W/kTq+0PUw4ma9mGF1
woC3dbjZbKNot8cW3+O3/bU5j8QcNlKJocp0fRIm6g99s1xOLqExvgH3w9YQWAWp
Vc2cgVcvzEYXmBveDR/4pQrnAZdWizjdhxSLxFw6FTNgRTvTvwTozc2vGlubJ4fj
rFre0JKQdUVIiqBxV6w/CnzRvebZ4vHqUkt4F6No93qXuRAOW1zFqUXev18YvMRa
rvckRRb87ujgaMATC/EBJBFwLYXhqOxTMyXGALdqhfD61yHmvOyNL5WBefVHZ4Wa
KTJ/Vt8s1UTVdPM6v+aNqrBhXLjHQagvRZtfq8YFm/RYX/0EthS/aAn02Py2csDV
mQCJv2y+meYmCWc1L0aTQ+aBYm+89QpvZ/yUpA7uSetDkMBecyiySHKc256gcI5m
l4KvLOhuMEDKeJyDnTSrLTous5dzVmqdG9gwihhjblzouLyg8OUCGwnTPbzhEh0H
MOhbTvbC7p17Gofeep85hhMcPH4R9jS4rrVc/43cLojnZOGkE+QDKcVXBO2dLJdA
/kL38YSbnIUUN8x1VpIqq5x6KszTSxPgmDNsNsqAn+XO3mJ5N4L1vYjHGubrVmPN
ibrYCm5sp8tiHs3iFuH2jl0C3tbLSM1wRz0UqZ+pg2nwBbPkhXqpvfTv6Un5wQWs
Y7a+Uhg8ac2QzpRzkDVLgUuBlUNK5EVsTfw99Uswf+z2qDNQuEmGB6c3DdTJXIb+
D7qYkNTLaXJ87ad+rKplGfWdItZXUo6F8xp1zBUGWb6FGfcOtDpT/dWMoWSx2oJ2
jwM2IZfTKwjZwtN5nh4ypl8lDaKRBMpJkbLpiFhwvUaIQ0JUHNpg1OKH/2HwUUfX
HNMiZP2gk2hhZSGeYjSoBTzFRiYIztsp4dU+7YerUmDZWm661RTVsB5chatuo3iq
EYvIbBgDvt5u7uOwSMCsVEMPE0BMPO4fM2FjgmdRvrY6TmGhRGvi9PcDRqatcLtI
Dnlxwlu37V0OJ1oG6vu+6rQG/IuqKqnM/mbLhk+t5CNVuY+u4ZBhqLSBnzSi1SOT
HaBHU4+gsYr6PTxz+US7UBxKZogeyfgDB48Wu6pAbGNc9GEKd/5FCBngdrx7aDH4
CBMwRldHOaT9ZxPzG34G0QmS1eYx2m/pCsiObAShzhB6Y8ZDg6m09/w6Mz7RkRcU
CK2WYNFJTbbKVPUNnzHkFyeMHfErwM9ppm8qvBkmuScYT39nlqmClVDwzdFuIb3U
bYpasVx0Eq3fXeYD3yL3yVuubpIDMNiJk43AiEY+JZWFtchVxOGz0NwRroArCUgB
QFUMndzt8lKHi1daej9RwyiAiltPQK8UzjCUpj2f/s0oPF4tg14dSE0vxGyjvUsr
lMitKx2MvlGI0z45sYWJXqYzxA2mlWjWKwxBN61RtNLyTqPToqJnzBlkxxaPvwIa
1HIKO7Vyjb9w5SA4Jc2G8qfHrSb20ZmcHZY3Li79lI+50nCtUr4zX4m06stoesvz
KQff/jkBOyeS8iuu6hI45a+KF5qRyxCf0r0K3Fs5pR+YVo6G0GNlW8PiqQ4gO3f8
zD8kbEAAPHpVY9zd42iNAVVgqbDwrZD/J1Q2X3UdMFSESP/arPe4dltehJ51YrMU
3PmLoAQ0nMNdtXzoYFjPGr6lrmAb5k2i2HnLhN8scsVBrnlvfp3TZTE3sRuELVQU
J63PcOfpOQNpkWYTLJjxtRS5+m02F05cZSXfUL3ZwLmNsF1qwNhDERMlQB1xE+FL
uExgikFXtMkyG3Cim9EjfcUjiuQA2leliyvNpk+oQEhgSZZkXBKnjIbcD2Hwmg6Y
byPZFiSQwTq6ir2RjSY9S9Zowo66GqYSBQzHXVR0jWVVNPEkigWM/Iu4M5LqUiXL
TmA64osPTSSJ0i2IR33v6kEhB06jTEH1PacwxcyV3ElfBA0zYjs8ZkC5wzKJ3eFc
GvTTT/gbVwW0aezfRKFzhpcEjohTkWWPKABuHBMDZwGKFg6bmgFUUwfqRYuhMZNM
jPOx9vyBIMQMpu6UcWd+8kCnZlyKLGIurcnyIu8aShU/Z1CLte+ZWSe7t0Kb0Zgt
/Py95BPcZsKChTMIo6Z0NhyET+d1N/PdIV++hya0x9elZC18//nOTGnAcTgeLmlR
7lAyZqRnvj0g6t7W0kdwVZNmf0EMeog5exzthOXHrcluEpV+j7CL6iPzJVkxrb3c
AgAaoIEadrELV4xnkJYegrXccAJCCws6d3jz3dnvT9bUf2Ui7LFwWnALy4mjl4rJ
AX7xjCTDPWxbaPQWM9bwifJSUSOxcQrhhs13b08uVE+mIJNqC6DYiVvmYGkvQ1iU
EtzunJmn9qIuMxoJPZ/9eNRIRNCqHHui0wT474u+vFKpv4BHmfcpNZ5CS66VK07h
jICR4M1ddmbqsjQafaDYqaBHHtNSHw4sEK6I2FjtPAm1zUGVf/v6OZxOCJ2cKykz
swz7d5cKqAKTKyg6xwyt2gtn4VV0pk4euMoufwb5HMAIegG8eu2EY8q3XCqAp8o3
tsb66JpJRVUsiXxIGF0HcPSCpDRH6dgZxOIPkNu3ogl31wrGOLIgk/GpQbNiPSeE
v8RBn09WsmsbbsfpJk4e9LMt3suR7pPiQIHTB75VTuXl8PIPx9C38uei7N8jiaXB
whSq/+pPfXhFGr/mR9H162p5bhuy745HU0fD+pCb6Ej+5onY+v5rSZdjSbnKcMkC
KCd4ijXBUwzxCTqmnlnSivanYGi1/3NknFcgao9phd4t4EyAIsIwtn0Wp8+GXrlB
uGBrNL2xdUuenKKfUqZik9gNk8cgffD01smXdPCndYapkh9i5UsVPYvJQkBbW4NK
sV7nOqhDvuFBApVxSw6Fv67GGlG8SmfWTvYA6BPm4IG68k0+kFbJ5LiPEMFfrm8M
FtCkLJrULkWF/8Sv5Ils0Nl5YR3RLtfX76QCJOokLEOguH8cBF090h0RAy+HP9Fg
h3qzV4kaoGrsUXVxCLDEq7FxzPqhupojfZ7m/UhKfU9DdoM7WxtILwxw4Lhe6FYl
G0PbJ/oeiVmkQ7+no3a+tKJhE9F+ZWFIBl00ULTa0xjzkEAWjNx+sH9aSN8XV0CB
2N2dqJs8nD4aY2yHPDQiC3RnKfElw879sznIfWacJHu17zq4xdjizTdniNvGowya
gY72XR0iSYF1h0h0zCX1gLOTMEF9/D6F8c6Qu/xfmLB9rPO+k3HFR3tmqHhNrb1l
uhoV3bc11HTxvZrNY2SgVC+rF7tbzB40gIBfr718yJrTS3xgZTzVK5pq8L+MMGsa
mccF1bHzDFNC8YzIk1zbu9g1Q/cXai24y9TbEezTnLlZfCgGrNXvvt9VLmcjrcSg
O2Mc4BFQExWK3dyN6cqaSn+AQWRor0FmPMqvCn+Z54VROvMsbZtnRqEQMt91Yx+l
Zj2lSy1sqcXdw/el8E9KDYoSCnyIZIAKpVMMg/nug3SJTij0obc4xBdGqH2yX7gW
JiFncPYwC4gnkDh6gLEbmXkCxN4S6JtI770ponSGIPv2VZzB/vpqcuQ+JoBjHdrn
9KsBQjN/r6vj2CP3IzKZ2DkxQVvaAfs4LRS0sbFVGQYuPaPt7AAMmqrpEjw7doPb
l0MJ5UiCChskmVeikSkvG537LwdHscPpSV3/9WrZvc9FJ4QJhUQG2tp27HDDzv1T
EEj0MOSD5j0oAmsz4QtolSvEl7pnCrDj6YLYNGpnYGGVF4HX4UoUbJjrEhhLMxMG
36OHurCs2+7BpTGveyRwnD4qY1jrnbQP1st3Dt79vnaiV3UpHs+tU2qDgGobpIKa
A+GVt9HZZuAF4uXocGcku2l4dJtiOqUPokfrEtTDJcHnbLI8NhnR9jUMEAWe2Eyh
9ZF4HS1m+HYqpaoie3KGqqLAYR921S+lRiFQ6aknvh8eVyNq9xOS/rWTqwf3HMoq
htE2M/3z+APGcHXBbHaahHpEDrhUp4vdyOAUoE0DE6A71WmuTs8k1qlUQOPvDpAR
g+PZhtXmDp3q69sKANiDDyGQbmwx14rq41jDIgTQjiJgrRT0GCY+UqbR0e/IdRdb
DaIc9zAvPzPwsi9sty8OYsnOgFf3j0AMT1kBQObP8nOm+nAOjsJLvJZuDZ0+Bsge
crxaigQ8IM/Y4cH6yWS74H2ANXr+mek32bQ4pdwFI/eeuVdOc5VFHCA+wDEXNPB6
rhT3aiDAm0Jk9syEcNGhwm3Ocb7sgKGSeCS4+vatfmeMNYMcX0soJSA1eRqHLssq
fD4fumroS0KbSPFhmSGYNzKUjsLWhTnLx2o295nmMSoBW/qSYud4OFBedipUXGZv
6pHRDbnLNn3RzT+pxu/rHdzzwyCZMW+JXljh7mejoP1ljBtZbhLn+54esp3H3QUI
6NePSTrz/E0owTGciEJ4lRaPrzKoMheOt6Eatv9BjRmxz6JdjB77K6ExOHjEHBw/
oxFt9fuy5K1jKHORK/fodtiCJUTaTGUVZQMm6fgLT6VEZBjb5FpXNCd7t58xh33E
d75m+Cb4IChCd32bnaLPvZxZ9rFiOj7vRDX6zcv8dL0ZppeEb631UuXy566KnLns
csMQpreEJlo6cMOwEqZyF0itaWW/msM8jmz2GtXitH8Vp/rZotCyiQARb+pubwvx
oa08dC35Cv9kT8F0fk3kvG4e6pUFN5M+eNdUfUwgJzBq4QooSwiD11M/IDkihU9E
KAiXFZn/YOB6ihxkF52Ib7aQZRIkSo701tjyFyF4zeAQNKBEo1M4CJ7vPR+xbr48
l5iVUpEp+3cLfOyl9i0GXTfXgZIagD0UOc+SsRzEE75DMn1s7EKj1PYRREs1GoHI
JHzMA0U0SqWOTd4I1tJzyuWNGXhyE+ECkhz7zgEZFqzpkAYQbIGC/Ozx4aFMkS66
kUsB49Mb4SimWpNXXuVg96ey1A23hUl16WW0y7SupjUz+WEOJpRLe9PRT8/d2krq
YIts/HwcjdmLMBVazZzj0uwzH7Zz396keLI/ZgchqlLiG8zWJQlijXH3Y6Ixk0rH
Ip5S88pSjTzV5dkGiQvwfwjkrLnroT2yAEV9j/GlMgKEJFXNjmIv6HKXsIl/cU1z
GQia79sdhLn9Qf0sJiTPfc3SHpTlEq5igLyR0WvWgM65ti6ngMADoj1wc6o0AstB
vSJRwY40A5E8t/dAkPjundAM9noGnkSgasuK9A0UUU1+vnkjlblY84zvuPLlOgzo
jywbMri4lNdCli/0KZsdhQjFFptwW8mLQNIFT/JT3CZCRciROMetRM4yExv0Qd1r
FWKOkYjOWI5UdjVV/389McsBpey9288x+p8lR5s+ZDs/qwGq2/u6iFwh2CD3Bg9O
C4tYR+4LeQtT2friaNS1QAESTs5Pi/fir/k67x2zWlUf2qHW3iZmhqkJzvD4Q+Tx
Nj9LpZmUBgwE8o1jkE62XaH/5plomDPGxoszdcLYKPojy9GhfOgtVbd7lB5fiqY5
efY6K3eJa5aEhy4DJ1JvxUTmoU2QoubyvoDXtmBxdfuBYccZgiiLKTjAgH3ddfA0
8mKiJvQp800aXyky+T3X+bjPokXiuXMbSl4p2i7A2Wd1yDJKvXev1libfPqQPPPR
fhUNr4+mPNctIaFP/S4mvW9haHfrHPGxIBnPlQuAmqRL2gsEBTepxc4j/ify2F7j
NxcA6aHmMxQnKbmoGO5kNenSxB/06GjQ5kZm3gu1HO4ueSc1xUcT46yrrqVAGFNW
nICBWsoRHeE3lc4gp4EHTIFCqk2TryrGJP3HtiYQuhzba2f8ldZuoodxSHN3RW48
3H/fW4MPxZHQhQHAYXBG+vJR0JqfCG6jThokf1F0JVUtq7wwUZ6TSpBZ51Pfs48b
2fJhPIxrFe7deG4VkwSjTahr3ebspT28WP2RMgQDObqil4GhsB17Sz2thR71f4QF
GIhjglca7xl7Sz4WPxhie/7RXlkOuGI86auRawVseTkRA25Jboyk2toIqrq632dK
a0dCuZgfXGkJjnF/whVcpPgnNSBq1rCwV6D2gTGBeAFJtUyc3bqff2aRWmNjPj0T
YwNo9HU5YWfo2bNTexC2QctGSb9vLqdrt/cyDZYbuoE+tLeijzLnr0DRiTVA8uhO
3RruMFtH7tQcstqEYv9aHQERik2ZMAuOTp1TYosJ6L84JsZv7S6IqvLOus9/aV5x
KADi/07sHEBDRbUeTyKJiY26QRxQUVqC1ClvQZCIPk4RygFLJqOJCsNXRfPOsNyr
yhxVjVKoFBBRwlJPi9T5x2/88iSlKCyOJJoqIuFaxfCstp3LaY7i9SrKUWaS9/fx
5XcTkluXDBVk1qWe/XBEY8du/1KbcClpaEJOOqgPYA3EZ7d3aNCF19zXUSnG8lrm
ayixRQ1T9ZwvWQJ+Q3bnvFzQQybtrvsGIrI9H/3Ov2DUI0knH07J6FqD27KTW6aE
kLsZ/3k04MsGEkyxiACASmUbBcrtm1fe6dBZV1B5/g7IH0r2/OX4kRDPLM/a4DxD
m51tYX175RrVoL4VBxvQO89Vi00YiN0+a3fpAeLO9YaExJCYDdkqkQ0RvFHtp3rw
XdcfAoCzJsY9KZWXrWws3WlfJBIwHPEroMuI4sg4GXQLMw5I8AVqVwCd/H9IuNA2
Y+r5SU00zRBDyldZolaehjmMST6R5PAxOjmHIaMR9c+lR86I67D0K4w5aYXDngv5
MTduXcOt8emSxc6lMMtS1V8DN++dtT0+u4hGbPT2nEhaTtUvPphbHJkDN34ymOTt
m01lqOKs1auN/OjMd6HWKlgeIy7OLLoVdxM6VJ3byo19iwrLHyz8pY1SEmeqGGSf
r60/J0O8GR89kCpUrsRw2hH4l74GyhRI+H6nbfHk0ipgiyPvtoJdwj6MNir2ZiAR
gmmM7N+VHGpbFPwY0NcSKQm/hDoIxinMr2ukIgvvwV7tosCn253x7Y3YWLXGAmQM
gDsSRkizmxqZ+EoDIYz4Pei0hkXT7b9CB4LMdyGUiM1eu4n8UgAe1PtfJ5NuhvZK
SCylk93KGFSH/JBlQQGG/D2+Hpwj5CJJ7dJmxXhlBY/FeC+SAaBzohPxuBOA+FWu
SsfKU3R5KJTUgukof3KBbHEyRWEH3hrQ4KMDyNPmavDhLm/+RP71Bgs2OEp8PL2d
K8mAd7+TXD+e2EfzQMbDwQUL3DyK8M7OLQ14KmW/lX3QMnmB8XaM33ri26nkxSXu
vY1w39c1uSdjO6CatcV8cFIjzj7EThEBRdAQdebzHh+F4HQR1zMtE0k0ANHj6OvD
vJY/HNZvDRM6xvRQLmFz9iqx9d9OYKHruCXQa8rUyDJn2rSyABejmyteaLdHP52A
+2YDzfYViSzw1eP/KODt0oW8uaL20ey/mTTF7v1DHZGxcS2Ert450yz/8hpFlQ3D
Z1ynag3YGUcq/vJ1OA/UXLX7uix/TbjBn6HLadDLF/WDeUfqwhLRBFUTpDRJ+jt8
H5XPIQqWPgiyL/fvTabLZswtyZkCW4OpQ54HUrX711y2f56ADoNiNnBgQP2RhzQT
zAt2qVa7nYl6T7h7mCR0zxDdee8+YOFDxA9hZoTGPJHlduMJCv8gGLqihqtcLRW1
1yG7xkJZzlDQ5n/mef8+oy9D3Ru6uznqVWwhlxQSj9AqRvUJWYmHdMhJpbGDmYx6
AeKUc111iHCpQDFesO2RkqFzqVUvgjixO9ZZVhxkEXDiKveX7G+O0iMwEGb4h15w
jaGBCv2IAQt9nH0PX7wKoHhFLQyuG9k0EzEbMMA5eC+cCTd+6XspdMODLlbjJj+o
fyg8o4cdkaJqUESeLTJZR7hOxyoTN3kgZ8OYhgvrdZCtRAskmxarbMGP2enTLMNf
61f7ll9Om3RgsB4fwCfHnHTgf6CBT3RdGSMWfA0E7ApxZumGvkpKENyUYnx0W4O9
Pa0BCt72m2DwArkSggQi+EYr7eqZWdYUoZzoeJKO9LqsR7Ip2ELEEKhlDngBwz+j
crZoLe1g0KzygrIYOUnJEjMmUUIUpWUGKv9OB+2idSyb1Q6v4/Jl8VN/OjFIsctM
4ojX6LJ1PJdqlJOAEA595x0J8T7tI06yG9TUUlz2w7lXeUjj4B2HAQfFzNghh5mN
DIUJyiNODB9cJdt0RLPKjPc68TLrw4p6XFATTNGm3zUSETsSy9QDNqFoNAtvimli
VytUkN5I/o+pMiUvcw9nGOqoo0IZC46j3YAnAOvYV9k778V34vZHbAHQUF1omzPU
ha2BAyFzAX5QBtTRz0MRqJBmc2qtFKitl1jizz3LV18JWDC/IRfFIe4bR0Je4Fo+
1/9hQ43lfYO2KDAp2Sx9iVCPeZFr6ZI38H2XHgj8DV+1a3GlbnMMGvuex6kg/x10
F52cDtRo4bcWlQwOgFZ5F423Eu8s86DTUE1c1BV0mXhNiV9bsUy0IMidg/UfcDeE
mvCX5VEo0AnuMNcc1SoKG8/HXF+y3fo7sNsRRKFTW1A2lBt/xP/qrzcfBLgbqJSQ
W9xz1+Xu2Q2xSpegYFXyKrm2Y0kjX/0B9cpX1LhitxYsGyIIhMh1msED1quNYELl
ZpkUHhmonXSG8cJ3TPN9nfiWfy6sUQqqa/9PlIIAHB2yVt385tz76ouJU510PolS
2VuqshahIE0MXprrrrCEluchZ/QHMe6B/+UnkoLW9rCzBi5AOh9GbG7giyDeVFpy
dwyKxoK1V0BBfu9dZzDbkao15IUOoyWTrtvoGME6/HF6+8bf9q3HoEqOc8p4yx1q
TFKXfRzl7AOK7p/vNBfGu9hOtrF7ZTglwQJH7jbCWdJ7tw3YqjRRG5LVizG/upXJ
pbogb1+FEl59S5tVcD0ZeLqfCxy8JQ+bW40KcrEW3vKpTeGICGu98iUsuS20bsu+
+npartQUIq/AY3dE9bNrCod8Tmu7vP1aKPZuYnELE06oejh6MyM8Cj9+RqG9xIyI
DjUww3gDOrCiXks7yriEA4xt4Hk+9QxE1gROWN+lLlu/sffCMpf7qEBDM2q4ZRl9
Zw4RAzqAYUrE5upGAWYX5VFkMy/3L3tKRzh8kVrO6/cMYs/nc2tVnqj98VJn6eBh
rZELjLrJOl9y8uz7Zx2tpQHhZIWgDm90YRtBl/4kttlWGRXds1Z733z1vv9c4SxS
mY/fh/eTFOEL5Ka58aeXfrfww4CHTBm9+3lrbeIqC1ojYMZ+CT8Ff8PerDUd/dHX
W0eeF1mwWWwpDivfhrzRh/PaYb+MiRCTvFoSKYxwFSrx8er+y/I1igMS4If3i3kI
iyYeolSopceUGmC1hNrSBKWoPQGKBwt52DbUe/tMUA+HOO+FpyiIwtkWd6EOQYrP
Qs3C9I11uQXRkw/6d3lDjoIoVLBThjww9iTtPeIln8huJRXBVmYbAKx5JVNhDzX5
+uErX+ZBjo1HDd3pHg71OBy8iPp/v24Q0FPxli8P9DTVimMCUYDTsfyKE56qODDt
Zk8SaLsos4NST26a6KP5rSOVPRaVMTFKPb/eZFLQWlS2dmoLlRel4Ux4E0OT/ue0
taLdfQpqeV4K7q5hLzWGL8i63UIDTtJfg7NqzjpPhFPPKN++QpOtKQsxpdg2MhWV
/XpcGn4GxMLmQ390lK9+angemy5SnTwHe2E/C00M2oIxHSPhpgvTSfx4IpXXVA74
ukBxl1x94dq0/qwEvBDmxTkNi79uQKn2i2ewTzEqvLQ9/FS1QMXVAjAc1fDW6p/t
X235Ww8k0AnSXizmJtAHjJPqf5xRjpn9T2u57NxL8URXhPFOHHRpp8YibTF56SrI
Vw8bClFJ5T2J1v0uttwXeQao6mPlf9zFNGnMTBbbg3IrL4cCjhd6XRNhB2WBRbud
qQ5zoBbdEGzkAC5UYyMypyalrbTBQ+L+px1F48cWw47Tu34xbtj4/CyunhhuAhlb
DD0fr4MUOAajNX4e2GZp0tusIRh0ooqG5a3bOGKr5f5JkqY5qnC4CWXEtp72pOWB
yz0WBdpL7HxMBdWvPpncT8E+vij8gDQV9xcflq1s6I9DIgkKEQ1D6wQ0y1HFV+S8
NHyGhPI1u9hav91hUrySFuJ1duGHCEeIGMK/1VNQPQhFaJVR8es1ZSOQnYxgsy3J
9JbP9bAC6p8YNYXI1Y4C6FXb3/mRsRRzBpFbwnZkcibKTUG2pW1EYt6JZf14OLeS
Yhj+gtykl5QcwtPZXTQooVM0MLe8balRUC391cHQ0/5V3VNZHQvnhBnIt3EkKOGT
p6ZXxdjbRqhdMUsaHs2sGxemjKCgCUrlzUh+2naA61Bmm2SNHayHjvfwR3KScsS9
6OOIhMqi348QWGYTRITBpsDuhmnHkrG8UhIsO/UJe0sMqD9OHIBHV6qaVmeOWSLW
hpcP/eixvs2zzsYKuYnWT2BfzJaiHbKGZG92YM2CKjflr6sOjsq/TN9zg19N2zB8
CD16DMU8OCLF7SwDCyF8jKgI3oUIOOsQqsA8lyhpD4eecwZfm24djP5SYx4pKUnr
xrvXcQayDKYqYygMZ9UomlkOFuQ8+iVCRJolbMOT1sqBRWMSxJLvT1FMqZkP5yuL
OiypS276PBxoUoizu9FYi83hYwM0wwzA46XYJWnFWkjexmj7Wov1Q64FuITJfP1v
c1fHoCw5CEzLUILYJVfYG5XWocx8PiMFYjvGcsqoI+wkaJOtkqRbW/Jge4KtGqJg
xenKl+TyhA1XzeCqjJqYIOgaseTiBkDzDHRNPF3+C1UM9WnmjEg7A2gfd9MijC7G
mDfKRQyvdAnXRXwOaoRiupxEDTg7mmgQoclE2jXf1w4CIiHhwWj1afkc0RvxNImV
Kvi9zX2WpAPWOhVz+RYWQhVOC7LPNX13yv3ixihErysrpRRCzRGVOJ0mNq/JysLN
ckfdJ1swaYZLXJZgCJLOFFViTZsclawQbC2ZjM7NzPI6qq+vCCDcVLZJyc7PM3TT
9pu2gDh0qQgDoA8Fbb9RoORrjFiBZB1jY0wfQVNJhYq+9s2zmyU2l0pq4wvi4mDv
s70ghMGMILz8pytCHrp6VgnBXdZv7/tDPmrknaouuOtbXs5BUzNHJvEn33phYFQs
0Ef4JCVcrrJO8UHXgnDrm+Rt+pvdd742D6s88eitpZkFvA/lr+PUdRDa8Btg1z9x
7gdTkcloUXow5CcFnfclL+V4haaw0aTgJeL2G70Wu+AOeK9nLIzSlc4eli4qNGQg
ec4w/E/5PwA9TdUKy/0sgV+ljCOSQ0ks+tMTdFF5nIwpyWGvjEmjWwPzXWZ8VNUM
wdCoztEZSXfSJmiDMx1rq3Om7XFrHoVg7KnjL1twPUbWJesYx0KEf+6H2xmwgcQ9
YJadb4UunTPfwe7NeNsygbs31MGCc5AbTJnTMfTHyhNKQwSS0OQELm5H9fJVGCTN
sIKLvbakp9KQZ4Ohp/oUmwJcm3Dlp0UNyUzZnhPKzYEdYxS8dkd1siGojOeE+EWH
iaqPasPLzbkXkoBPoDKxKT01899uEXXRyEjsRwNheN85rzLapEsS/Q+1sWFaD8ye
+jm4/W1m8BpvYv2Rodya5sv7wZ7TJX+X1VAK4K1UqMdIixD7A/PAgQ6wd3RGyMC5
U+d9GDDVYpW+ZlX5+lwWgKP6svSPgNWAoiL6gLTRVOZ08Lm/tTaHwe5C9oSc1LmL
o9vmBxB35JWtH+aARydRGuVp1JvK16NGnzL+OWr4Q75tgrfEx+e5CCde/dJZ6cTy
Sp8XfNrnPlMJh2ITgdEIQi0X67ehzNEN/YinFJtcwNGUJWtE+G125rIXLswicdib
OK4yCfD7KC3L4ABamYzA+nd/I3NsbTw111u4t5Hw5EKmL4xm23cBT27H9GsY/3gi
c5aQZvqOrJDSiu7uEWSeLa0U4a2qdmgeZ0Ris2uIqsh3HOfhv5TThr0Pk82lZFr/
5JNOoNB4C//an8iEjm8nvpVdaBU0KzfkwU4r5Mwo6tJp0QnswAQXhzcIh8bM6TjH
IyqitoOtVA2RGXTbuMVrUnoEaEjXeSOrT09u8hSQqiVprsuOiGsWst4+zBwF+eMD
5NtoQR8+8vY+0rU5ETZ4qeryt/U3I3HCvIVKC/ri4Ra1x9caTj0g0ngby61nS6Vb
8xZ14t6KLTU6E58IGg+SJtiSuorIgtPgc8Y/JKnJxNrvCpcVO4HpjYIJbYaF8BfF
x/pPjdEoOO3nWX+u7SnTUxdW1nGC4EyijjhMHuXkoXkVXjTSxR5pEw527n+cJtf3
j0zxKyzNeYnd9pv/UULxF7OUb8vyw3YVReEt59FgQNeGWJx148gtPBmlGzmB5RDB
5HvgyS0UpUbjvBpJQTXE5pk/VUTZfGer2BOVZ3vE6SvtucUA+4NUlzkEUhS3mKrf
tWN3ZdLDvpazfVb4xZHwZP8VABfot2SDUZvtfSkcxcFDx6zq93ODUPbhOQVBQYPp
pnglc6kAqADGKkiWK85dyZs9eqNYsRRSpSjqboboyNRs/2ZzQ+j80J1rMSZKNCrc
OL08JmDSAxanmnlbv2TSOjnX9FKAUpnzJizcldRoO9qoIM99JF20wBUKDpdDn0m6
TiCXNzvkCn6L9UMTFHvNuFUnKf1qv+XYKRq58LsclB9QDNJtP3lnyBLFingGVLZk
2JOT/leGaIG7dlRrBzXSknI1Q/p6Q6eQLWM5NeOewTKLHc4R8qY94cN+oMqQpGsC
psQLeCUonzenoRnBgF9MgQeNRRqDQrHYxFc2NmlJWsyrGibewzw1rDhhvNsjz2JN
zP8uCw3s0ncoHi/1sKC1v2AHaGauo7kmEMeuLq2agKFx7NaJQvy3dTulxeLXXqhZ
mCJNcEPbTLOpRYfG0K2ePhwzVORS/TJmhChNAgatRWNiRLdzdSn2t1SM8OTKY05x
hnoeeSauwC6UkHoZEmEsip+mEDW5f4kTBYe1ElbdjysB+hqpsbnvdn+LbX7lgXxA
UgWgFEntccrFeDi0GxzuKgLhkwCOeUVsT9AyZOuRqS+eR48HOzCQEDlibUiLr8hz
nT1ZlZBRRfys4sQkbN1r7obgxUJXlBdvAmgF4/oeR/eH8ls4Bk8XAZD3aRyduT7X
yWTVy2wQUdJMSZuHZvHySWrUFfTFsVTD4ZLlM7xLqPvmbIL18aH4R9sgznsfBh4l
++BglckEOT3Cn4WWCtXpy4269gF+X2WJRKoCQpXgmopnt0HZ8Ae8m+gqKUgc43fj
ojj/uJaX8suE+LAjIyU1S5DKS/U6ixbOaNBjBiTnseJd71cX08LclvAiTdcJM3XO
phrypUiiP0pCM6a5yWwBgCzigIcMPlnhcSBLIp4jDU7zKxFQfdrrKgiZrQX7OMcZ
SGQU6aDZAhFT+WU4Fac0tSIR7idY3rfl/dCWeYqWpnfldb+djAOjFOJ98V2thsLR
5UmWg8rD6ZiuQB50Jd2haIXRUVnkvK5F2PjzcxT8tdyBGExyJP3Mrce0MkJ4piow
xJlx2FQkXY7VErLizTLJ2+AQF6YUYu1a7MsTnyx2/fmPLjD64t52zMAruVBum44I
PNpMU9PqqUjGF+XFzuMepygC6hzsP0A0vgY1yMcqgxXbIdWJ0HZBjxDyp1a/cWkb
3HI6ygrmcbH769AlL/LcnaG//xujnTtmvvThMk2GSOen1sx/zTWCm0Io6ndwVfoM
QfjvzNn3gAZsYsOIsgbgSgIH+pBva/XflVYJZcnwzL+Fc/Wz80Y8LMyDbDhKKUWQ
F+pEwyZnFNssWLvg2yJJCBxxkmUJsEczm9u2Uxr1OsOiZqAOT5TOEe2X1kx6spSK
/Mt8zs0wNlGckITD+NPmwndGKVEHloRM7TRt2127RstDZMuZ3UfVnU8BvpJBvbWC
0qiUA4v3TKiX6J8VuSkv/1obGQJ/rXi2cjE6lT2zTB4HAhnXHqyoIY37lDcvyvDR
3ZgsAlw7tMw/yW8Zb5o+79LZzRW/GErKvkVfrixvZyTpuEAY5b4rb4D4SSM2HBu9
CntqXf1iAGJbiY8fv9wu7IxaHl7LTa/31ekLozC4d5cinJoFZwx/5gzxP1vrGaff
nSV75PXex2DRGAd/n0I4Otc97Rl3J3aFT8cfceQzImq6lcGFEizRzO1WTaflsHOO
Qd3kSm+OW6gQKqyT+EfhYXG2F7m4GqOYW7NOjsd6CeBVKXn2NNLB1S2QC0nQxnsG
RzDj3/qOmLwLRz0bgxXwX7Od/5sfIWTC5GNFZBDsR9acdbsiUBkpHhRcquois0mF
LM+herLmZAnQHfRDoSj8BOeAIzQWz3ZzTViWWaFn7Iv5nNWo8Zs9+xX6y7N20gK7
l2HIiN4M4ZrRKfzezIqhSkbynTcsQQcq9TRp0Z9WyAuhe5DbRA/DJ1narfGAmuOF
e4XvJNc8xUUOdax1TBJEsoYvroNBs5Ic037FHStoT+ymzloBXkkDBcV3ndulfZD8
amcK9ABdx+b3GCJmOZIfX/M6BXdh7sCJ/5OXh40UIv/ttc/bGKwf+0iG9q+XQXDD
9Zv2GpdCy9ks7nMhqlA13VBhgFzlpj6jp2zQEJ0x7wxJ2ErzYjCx+R3k1Sd7MnHE
J54y6uOjcc7ZeRQsSS+a8o2H/M1ZXKTpTZTwrRewzwN71VHdMinAwZxRpJHarrgA
/gY3gSNOFjNep3ZRsk0QqDOXfSBn2t5LIr5Yawm1ySq9Konvzmn8IBCS7I1Vvr7p
y/vMiQzUWgF8Z6ML6dwK4k7HJpsAsqAt5uediB4NlkpJzTIHNOS4BUUGz+v/gbXt
mksGPbTPU7lPpDYitSuGZwDkU5TW/1808GQnfLYeUa99/NYHZIrinV0c6/aJ5D/A
QsLnfahgGItesmWsbOx3V0AwbIiT2bZO/3eq1ZJBtoPuOvZ7eWcG6eOiGcciS7lf
NZJUfd/6s/Nu5hU/U3zvPzvo/Xp51rnTo3QMNkIurhet+YxQ2KTOyCoIj+5FsAUU
vRUipggJv7nD/VZLA8MHO99MWr4l0rFzyKNWrHO/w1ittVAYphhWD/1wf3BvHTQy
QaA6C2RGyVZyKkfOlUe6IRLBI6woh3NjBzYGvVqHhESxNmHrO+aj6hlWIf/WmoSs
AGAsdZDsMziIxSwnq717QXe3Ud8ioocsZ7htmhcncuF8kOGj6mlgt+PqR7+xX7SE
pO5HN+MVNzDvTF4cIzgW/1a5H2J2WQA2Y2zuxffPprNAKh0xu+vDxNL67a/jGIaY
rTWQWFPN7nTtZCKgWuJvhGpo4GG0I6aQzKSeSW5QmKAjGJQqs2EgKMuJtdIpq4m+
I9ym90xxegRaa6YZAzKwhSgItEjZyrsnojR7+8Wl7ueWXa3wv2RArTMTddCFDj4G
v5dmelE1S4/xuQV312FgKe8MnlVFi75jij+OJRB9RSne9odAeCBbNP72KOZZFfyi
icUZzIyouWJVEtMVeIbUiyDDh4zNKq6+3nHfQgtV5ak3ALdWQYZOTBdyVAAelCIe
owCeA7Ljz7XwTLVGWr5gg7fTwN7bjF+VY1CPWkZ71KzyrVUSsJAC/N8g0eHU6RJW
hdmljk0MaiDb7kAjl0wFJziAVOcdTfuyWCBvR61eAsDwHz7A4CfUo0bl2HxJCz2y
oUHEigdUEil+Iiec6a+UX4YRCePqP5H62H2N3qM30pwxgIEQCszZh5GiTa2eAHb4
IU/Sxq5zGJUx+YLIRzX3z/cYXeI/p71AK1ENUDzjZIG0qwuSIsnNPnMORdeEn/if
M5gCwnCXvjTZ5KS4ZA7DE3I4m/+msI1fmJ8Ia6HwiMOsiniHOxXalC1jxpxlV4qs
EYZYA4W3m9pcZfCnxXsL1NKJlpkuJK3Hr2ukWPWfexNtShdtUqYIlyoo1aJw6ysA
sGFpCIHXRC8dbyqcV2y3byLqaVimOvQ18FkGY125xkqqqV7oKs27GDZm/UQHgDvh
kkoevScX066Y4ZfGN7rZyuY+H7HzrUEbVWKLH4epWU+YOw8O6V3tD+OrlNqSkDSl
nXug/bAFR04ju1yC3IQY+UdACm+U8J7MT7fdI4I2YFBBBkRDsZoDZ15roAD9QYf7
KKgV9q5gB1okvFOWCddVrqm4wBPtwdnLn/hM60G94SdYOWE4EXLkE10bYEThF/zF
2mYFsx2olayn9vZo+RBz/Ve+d63ZxIJVhOjW5GZl4/HwtgxDDXb2E0NmdJVRWR9Y
8zSc6Jl4cxDxi/fAiRnxaYrGM51/C4R0j7crk4h+b9rASlv2mcasPYMSd/BUKv0J
A+hVvxAetRRnjQn59ChdX00KFhHIf2NDg6RmE4UdpCqZAB1rspgUEBiBQwZ4A6A1
wKOg5DgV/75IrnJQapNV0qv60pqOQdRXw+kfyXmx6Ru3UxBv2/etoeFMBHhmXTl5
rXt98chqUKY2LDlJi1lR5NSNkNTw6wBaG7e7veQdyQzJVmHktmlaGKpmqkywMapc
4qIF4r6kxYzsR9fZH1X6BliC3PRipJKBuiG0LVcwE3wxkOBBJh/csB6nN+/zoeId
aN3MU+REMIRUHhxcbQsaHeFOpVjoWfXFbfe+7Ttgw36Nmb4pNNePNr1G1EweTM5Q
LCrXqxDdg9UESgFKijFEh0oBYzjmC+wcM2soQmi0kWgeFV8YcrsERlS1sCkAvPdz
QX2MayvXX3QgiJnzxeY1AxHaeCCYNhQss+cxF1TWrlh5sBV06GxU6k4niI1TZrTx
ySpLG32JOQSUDCR7MKgFAbTrIT7lRRQ6Uq4B3j4Vjm3A9duNx9V1jczpAP3uad4K
GvpTi/nlTfCWeFJXjcjdrx4kF1h3FHhFDZjISdh2ZTGP7q5rxrpkFoolXKyo+Iyb
xPk1UXABIuAbaOT9iB9K1imA/Cs68gkvzsbxQEgbrIHpd7cDRP+ZpETpMtT6tnnn
fLZlmL3KRvSWED0/cOcBMWPEdf0SYQSA7ZNh8O994kiFh2xVws2p623X9+pNSMaH
CdGR6vrOSP/cG3XEiaTVxGifcFe1AgDdPkiTE/MEbclCxEKHjbyXjZHlu31zBrCN
IMq5nldX0TIF/UEJf4ysH80cMu/uShrNXghOq/apIJwR6r5XzQkJMa2P3OrTYic1
SoqNIfwyd9j668RZ6lUTuN0dU5Z7V/j2F31l733pViJaGj6V6DQpGNDQ9sFs8UAq
8gm27vVeLXF3K+QlRp/mZZCEkaD2CfkB962Zz9QcW/OCafrdIql7H5G3FV9xUvhi
HGW0RCUSa61vMQRtYcM+B/nB7oLKfYQIy0ZK0gHRqThDanux9HLKJIoOcUAU+BK/
QT0c5540HdxEebi2ocLb4gI2o7ud/mbrO5GHWLCBNtH5rix2gk9mXTHVzNL1lZ9R
gpN9M7NQvDtHMv7r/xXjrLEVG2wj3Ew1Og+HrMYHZnRQBv0ZIRTgu//72g+zx+ZU
SKKXu4a4apA01ELKim08DBDe1gqjqG2+iMOAU65Vo4pHHfSvwTPCVnOO0vqv9lin
5Bipr/nEVQXGe+SRmnEE5B+jmt//CpZ4XycxRiXevhtLrlKDgB/hUiC7qX/mHIZh
i0kN1aWd3h1E6MvbQgiqui/jp77Kq7XsulUL/Ehm1Cd+x4kF/KHsFpnxWS+3hXtq
yNfbNL19eOXDRf4Ol3/gsQ81SH15Vc1uzz4vmni8WgRggm60wDQnkWC2HgemYLy4
k6YQlpwvX6xRh37S+yD4vMbtjHkq0WoIRE16H5gYHXVAOb9pKeMROo6uK0VE3Tn3
K3nVA8sGhfBdwVZ6VTXZt+1TpQDEgq5QpVf29XORjsPb9M/znFhL3dffRaMqMDtC
tcguOgmShNvNflSDBoVbcj79C1qPYp4Y0rElp6d2tzm/j9TWbOCsdI9geZaCRlS7
iFczDbNfkOcRjNnMAq4HBV95M6IWdEBqHyVsHPrH39OTSXspcUqxxkkAOFwRdaTd
VN7qXV1uzq+jKt7pB42u1jO7QV/AhNPMOhAytCHrg1zuoZOPUiXnl+oFbRuybjSM
XJmp7mIgTr7as0QEHxHQ7d0vNzN521ua9x7f2E7iAUg6043Iubzukps5uEuMc4tL
mW4wS7mZEJei6ozW9Tw50ilTaDAw/HeyF0wcuAOYRxrOO5wi16gb6tF6ZlGa7emo
ec4wsVURwRYlTmLBhdzrUZ+DfDZwUcGrN757Zdwz3qXzrQrBfkWsWo0oW+boQ4rZ
q+iNNtbemS4HdhizNkt4l5+VA35rxY/Ro0fHEr0q5SQ/6xW8QWNd9bGLGtoxRQQD
9Eehgr0FSLcMsLQ8KPnFrlHduuHdp5nX+X/5iZ3I1wfl8kjXtIgvJ2yb3vngOP5R
P3KgRpxltaT/otzQI61sCeFZ5l8EiVwlf1AF/Ru2l5VkR2M3EQ3yzOk0aPEpALVM
j9NRUxehtmqCQHZluCROkKugPYXxoWSVUuG1/sqd0HGsykoYGrjH0ffCWT/PjOXj
miOQsgsM5vk8Noj7E0IyReUdnki/ZVPkh6qhKrM1JpIGr2+PTXC/PRyKnvHlbMmQ
evO0s40saOl2ExZZCHGF+6SooEY8UkukJPSbnzswssAxB1GeXQ4ol7E15ccNcrut
xJv0OwKlysM/oXy9ZmNqV3sAcHmLoBA1XCZ+laCRJYE5h4NMcHQu4oI1DUy9HYoM
g299N4cHi07LnYMLIeGfpTGVv/UvgZ3cyVI7+WCSEtwwN0MUnp1RWavNAGsRoT/s
pg29jrqsPa/AIbpwQs+eXWvGmDenYSmlhuXvHKQARnJtLyd5WOMSpK7yC30cMmC8
W61svXgoCD3nDGMB4Msp/BkNucg1DB1hbLuM50EegYuIGSllW7BN97vaYgZ2KyiN
EjynqoRSjQEt8bZTwpsA0O3Hmwim8+P+SvrMChh/6fbdG3dnhvpXCVzxD/8PAOZF
oaZk1MU8XAlf5BhEELzI3/VR6FAJelsLBhR2r1FF0FsUI2nE0N/2ayHKcnb0BDY4
HuhWGl4gXeoOWJNeGqWccPZ1d3hRZj6d/xkGW0tV6S8dG3IgLPQpkWLGzyk2xTRv
V3nHx6txcXcjteQi93D6pBbW6/qej7Ag9NkZud3Gw9BotxCmK/zT7QttZ9unB/J9
I/5yXiueWDm0pQgqkWMuLmWTmrLXTNmzO7cJaveAC8qnxhGy3YFtxMP0cVYqQx6a
yBZXP8qynDcf+ZTavEAxFgEM9f7GUtMK23VRPZDOW5rWolD+veLN7Tia7U3Ywxqu
x4VNqkUj6VPx8NDvypTmuQyMhwTN6dSd4aQ6lDlKXW2z+fzBO1pI4XTFhcaL4bDx
uPFvNYkdTLCdQ6CcBmbtyTtELShoMxk5GrBe+cYWeGqDgYfXE2h+S6QS36q468+L
q+FvVpAQ17x4Uiz2kfqifKCHNSB/prIOmZjXmQlzTTBHT1CAqeaEGctpwjUtdrhc
T8447xOYAB968vT+s0LFqH6NMA36jqjFGviLxXUzyNhO+gI0e0NqFyjVtu5WVSxQ
mDYUCdyeSCKP+/uOGmQ4Lvuwf27J/ZXsFubLkJ2G3mGZPpzkktoNEWZBhzMwqCbi
2K5E0+gWLUf4b7inzB6Sk3r77O8lZ2L+VoeU7+1Pjix40Cy4FHE5Kz9vvLlF5DDc
82EzPQRx9gm/i2xFWjz7YumYq7yfxDQbwNwnBSfnZ3l+3PigsN6nIxah0c00+Xx3
aLH1GlLKQ6rzgaiBoiBexpoaXDLYrzOB2FJrq3eipcCRaIN6YpFVUMqsJpY7xOzp
uAJURv1SfAmTyQrHvEll4HCbsyvwbVC2BWBs3/bgvLky57N/xMHtRFbVMYYS3qPA
2fpxtXV570PBSAFsgcS3CejgXoXWMrItAUPv1TsrK4B90LyQ443WnZbd1uWW5qFV
jAXlot3VnCOP2ymLDLzascAiXgAGMLB8wMUju1c+NGSZrVYw83mLc/xLeoWU1gzU
/xwBhhhAYGzCRPbl2o9aL5M0pp5Jpm+pruwnUKeWmZDF9KYd125yZD3B55ZFyO77
bCukHeVlB3/G+QhRcVB+9NEoSkDU0L32//qA1zA/kILn6KohnlJBiMO7DEJVXg2m
He9ToaorCY/2nh8XSGD5XQ/2MX5bXEJ82hkyPgfJo7Ai9UoSJXes2Jha+nqtRXRG
CwRYXDmAcLwvTkim/fsC/Q==
`pragma protect end_protected
