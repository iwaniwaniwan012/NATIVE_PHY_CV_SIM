`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Y0ExPjJofhj4M0xuYaAmC7SkPwc8c6BxLltibNzTCwNAgtNWvryAwwFSO7J3UMOv
IGZf/G0fC9Uu/E45EfUVmM9uPnaDWT9g030nUq4OaiphP8mCc8WuIvvxGYMyBtA9
igugUZnMXT8hL0YSli5Rp4dtOuFRbSHxegzhqyCpHXM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5584)
iSfgPJ1xwTEtFWljgf6YQWYvex0HPAk/0F36IABEh4zlC81GyFPzb5rNVkaO0G2c
VzgzNBaTF13uw0fhkDjjJikzHoCPgVd6VoUr6nlorSmUOXZSGRcyOtKwCJiKeNCT
70Ex/MXJ9VF/EM19OgJHqREHx5SdDzTYlzGBcOCMS29hqdSkXd8uvpZPOCvIR/hC
P5KT4yyGOr19GizIpf5nMCS5m5wiQtIY1kCXxuZ9lyvIZhmAUOyESAKz5VBvTjh4
T5ujnkTD7PqMBzsquaD1PFZRz5MUawS8CdrHmtsTodLoNREIriI3cINX5JHlkpDs
YLJ7AT7ExSxCWsNz12yrMkn6b0Zo+Ezq9MBxbnE0ifWdfB+097Wo/TOzY4N2x68i
wg8t1uBf6MK3mEGmG8L6Y/2kPuHI+G5XilKSDGOZ8/Hv8NInAU/+bW2plEUSK6YI
d78KeFBFLEoy+J3knitabQuJFeUK4IB2a5XJvYNFpMllcI1yNnreiDmA/rcGZeqA
Qp25ILMS6cIOMsUJ0zBF9kwkVr9XlZcKPC0vuhUyk5Jm5c+EF8jYvqnLu1cmcQ+I
CbbN+NututFjTK1fhAZpI5auQFz64a7M7IrsiTchFjsYmRXtn6kdmltTqwZ0FhwD
MfBNfBL736giTMTVEFh7+pfJpqkaRT2m4I7pWAcn27R4zC6kUid7wGTxwOaC1ksl
KHcrPnpXAuFs5m5Y/rqTxL8ETaf83osX2tFHobkoeEi7e8r1fBkLxjOJuwtG9rc8
vgyiytgPy8le/scrogZdKjTe16uYZUKn0OWarj40u4cCQu9BvFUXtslhEXfAQmgB
EFmVre2AucT2jR4giC1bbk0kU3GKgV8DEeW9PIIEGDlpvc/ycMs+SwCd3FPJiAFM
ziwLaeQVbNkqMXyPHYYL1lObm9tV9RmJ5NiXw5Xq61yrVz1mnA+I8ThZz5DqDPdd
w7aWRrMAFqy5+37BftFueDefkGc/OYNkyiBes7UCeCBz3V/qftY+zwJQxuNE6PGA
ilnIg3NWDO0VYC+XiYhDuww1paILhLj8sCsfi+1bJH1MW+w+v71TumjU4jpHDtJv
DFg4PsL0TykaN/NBKyCsrei0MH3AbFK0j4kzvZncdYlkJ3E0uNWM89PjLnIwPLi/
UCiYOJazpMrPz9XqjwqKkb0SyborytC6NFdIFMgvKu+RIg5H3BeErQc9c84kn/zR
fJkFy2jm0a90zg2QWFfOT2CrRbUmXHhpt9Wu+MWu2iWxudU2JiCQqwsJs5Zbh62o
cgts1U7CU+lEPaTtCo5tJSur4/i4U563eihs9yhGMkQgu6+h/ErnlG3TOc/2B/GB
6KpIUDNusUHPuf7JMiZfHHHTRu3tKHJwHI+lwXMs5Fl+q/JDupVEm8twHQgHEiCL
NQTPF5IHFjvMGrZSXLYThOh3/WDFp2c0VPMpCeYfDScEDofM5ObFd+5YvD2cTPgo
IGBtj8lRSIJnW0mSfI8AafENyNN33BDpQ44W8TdrNxYJqGaePBdPAyKXiXJYhsAt
Q/jegzSiAc3YI5OY8m24mYCwhvLfxnvlNemLJgqlmhcHTb6QRQBVwCEHL4yGRf0u
7zCmWgP+Uz0o0UsN4XtcaZdvQQ2/v9e6eHvd/ZOwFgiS4HbDp+4K1g6dtaJ5f0QF
TD1zFuMdNLFMO9g2nMDqJjHe7MCywerX72++9ZgfDh4iWFOI1iwZa3cjnmAu5aux
MlsJdVEKRRX0m9ZvPYc1GMZxxPqovHut8GOU9NCpNa6jOBEddwZr/gyuOvGjxmyR
zAdWlweXU95ckhZoiIlJPQoH0fZSnIm2YR5YSbu9kovrOMYMSbbvZ9NrfHL6liNp
t0l2ih8isPv2RnpFpuHmQ1jN9Xxxfbf8t1waWyhBJuF+bRnpIYKcmsGW2eVAPWTW
gIbNCXIyNDAHB0ag87PVx1xmUikab+RbGBfGmt1ZyS7PVtadA7kIKsypIh0LrrjB
0Gikxnt9W8Cyg7Hcnb4hUgOXMBz9t2N/cPnaz3GeoHWDTPuHSNQidDVp3y7/WEiw
jkxigGgRVgMEYC/SR45WRX1ovN03k6Ch84limCUsG1PYq7Tvj3xdmbzpwPnqqJft
fOcxKfSNcTEmLRkAY38zCMMXcIjx/3TRDQUq36ru5Mk+ldTnNcGFeXY/DZOtmJ6b
H+KGGVRIiuW26sb+G2rPHhJKXAs/odBQvf/NL0B328oAEakk5TrxSKYswdmlx7Dx
HIlLRTOJxrCi+ofoSquAk7mhb/QPFdj459W7xpx9Nq7+QfTR3WMDxMZxd3gv1pAE
hBIUxkxfDVghmIgZYZFSCUF1OZxczZYacJ9KzaQNw1XsRlmS0SLLxsi462xqjkoS
4YuacjIAwb/uX+O9TA59RT04PGnFdWgotmaATO3KrwWCOjIsWTNWPo6wIb1gljnF
vdfztBQJSocTqEOMUF09srke5oBnLKURbxBEQU7Dveo1dnFT6A2dS0Mg8HqPhaJT
bhHrnjtvek7nglmwlCTvDBR7NMYpOlxhPSbsN1gjX2TghGmhiM1008xmTXJY42bf
1cWtWm19H5Ag7J+t8ycSEGEiiKI6sg2g9u4UGRouvrStbhL47UgLmLVO7ETdk3at
b32PaOT4ucv9eqsW8vHPKcraWVgVsgCCmchs9JtLk3HPuXsWDJ1+LkXPyODdApKV
WV19vE8UKTESy8UYhbivDDfyHqT62raRywxdlnxe74q2fVl15Y1uzp24pwpl8Od2
hbRgppIbOgd1FODuExR5IcBZaDOS74ZjgecuOPUyrH9gLeun7FxnCmgcg2WUaUxw
x+MgtPnbuQehEZsPpLn8xS8cg0VfocyLDbCHlHs6bkZOVzYS29iHMlbd99Uw8FA3
GHSfxrU+FDoo8uYbEz3QMcFaDkn6L7ARhzNo9PulYQ8IOw1FnT3TogTZGt6TV7Bq
xEPqsZYqaepDNlWOxiD75Je9ERh351tI9MSCipC1hlI28TV6YZ67YlY/eBfW/91k
R8tuhCfoSABhVIrAKdqDa7j9CTPKDBW/Lmu+fYqO5Rj5v4iAMFhRMKbtGDYF5LQ/
1MeB6Uq5AEZYnQNOmS3WChIDCj1L4bDNIP1ZpCJaxb52Awd1aHmoc1igXFhNKn+7
cC193WvU+qExTXGp2rCwjrSVWvzMyx6RXhyqNV/fxK4/um40vsIHTI2Uzc8O/58u
hJpqz3g5ZjctPnq1CiTVF9z2cQQ4xbw8fv9LAbElNmZ1WU6TWnIP3MSVVJc1U9qy
1ZXKabQzy/oQsjxU9fjF8wNWDwGx/uteW4G5kCGdu1wt1Gvh6s3H/YE7DO8PBJf8
MpFyTa2D53OPUzXpggR+tkJnxaYI7vy8ALF8J4Zda4gthywm9Fg08S3DRF2ov5cL
WjFnZ7AQbRT6F9u6TXO1T85JvHCil866VR2V8hBoB589sMi8NA0P9mzKQT91wlKU
xre35xS2ci1q6gM+pBsm8gLzm3OEK/rjeQKsPVkQVgL3d3sIepoVbPW0S3QmR9Dt
U+cauTERYf3bUoOr7LNpbHrmMBD3IQnEkqzLHHghp/i4ddvLf7LTW1g5eUbcwyOM
gxwXEssihGVtzL+TVvaKddWXqBikuqyd6Ji2dycxDj3ZcPFfuleAgmhWOXrkWrir
eVUJH6rxmgcqnIZMA7ObD4Li6DE1niNX07TUVQDki+PAU30UxTfJsASfHd5niq+0
rbb+iPRNAEsddrqUSFy2atOXwECsRxAkV3hC2w/uf3JtPalqroFsr8abk0mQTB7I
5UZ25vzDWlKaKNEsY9Iu/O6gfjbdxsfqTNCQ1obZ1LCqQAASCBRcVp030syP2MFK
zDQtNw9BWLCqFmV5UFHHtro/bXZqwuFl5DXHOByCXHsadD/wKkXgm4nXVlfDezBF
9dXEofX55Hzxr1Zw9bXZ7rkVPzNDix6kuivcXdJgX3S6TNmZL/TswzK+4+8Px3ct
OBXKoZXP6/P0p+lcX16KhIt4vwbH3TH/H2qSyE7YBT50VnSH9bqdZrqPJxv3hnpO
mW62ymu/T3WLcEaTqG0wTcFnefyYjcD37QJWU0SF80RQPtRiktsUaVd/GoSlcIMA
x3EQy+XJ1ZI4olDEQvlrRGPN0dxWj8bfKcnrQUSNlmpQJMJT2zj0LpEgyXBIT0Dx
MuatJU1v6Oj2fVjbr+uBMunTLY26feAFuOQ3JKV7LgwxeS1kDXr3cuBLYEC5CzmJ
HdlBzwp7392aHPpvm/XIMTPfkYfnD/J8acDoearCpCvtSRVVNB+aCyamhk7mpkFj
00aqzG9cR0/vkGC49OIeoRyGTvBPS6mXCZcGlISheYF6xd9+ueT8mdWtjNDtN/ra
g1ypbTgQuKXOCnAYJM7h1kdb9pShn/j7p8/e7qFEwckeI6IRc2fSEwPLYTlyLjkn
kjdSKG0wvQr9NUNdFk9LOxLjse6e/CM4ytBEWLKi7GERgE4brNy+3AWXjKsxFHpi
LUoEl5Ebk4TFeKhjz1nQuXA1dUXh12ZwcbbbeJFjAReiPKikyVt3SFyfZXBmqbiW
Nj92lFtJAAdc8pQ3EWiDSCYh6yfFqy+PycAu7GUzK6obARhSAgHS9eDg0+wjMFxi
wKtNcSzp7rvHVtcXqMYg8XQLeSUfWN5iVSga7MQYmOe6H2XAsAv7LkTYAMNB4dOQ
qF5lPJb1oMk3uYeECHczqJVybuI7JdLH117+4o1mNlvIHJ7cnIgPRUFFrksoUKAy
jykCgd7/JmouZKtrCItTG/7AghRaTR5UZGr6FltteP7+204PLd75VWZn39EB6Nwp
BNDDFGOi0MeSHma01E7UyYXyACLs3PV3hI4Z7+vvcFk3IQKz7usoy0pQiUtLY7j1
kxvevEtBFuGsqUw7CKX5vAVGW+8gSVGqNfwAKSQwYUN4mzFRODHugPxqg30LLgRS
vD56lRmyjaKzqrEiQyt4Db3Se+pgl1VhJYs+NrhDg+Uq3R9iuP1s8Ln2s0mNtgiB
3oBDSUsZB/P91tZTxymHfe7qsAGZhD7R0N/YbYZfOFexB2zLWm8JuAa2TtxzuOEX
6qUbQnwgJIz6okF3hEKlZtAiAQKjbSeXAzX54Vo6E3pQSZeW6SuZmw4PXWhwlq8o
Et4zCL3phwArdxBUSccP5jZD1FpP3ONAJoR1ytRqh4cSVtsqLz2FPvavJ8gcYD6d
s0lVFPEQ5icZRx6nMV6iwMjsRGH38lk5gDBipzWE2dKdD5ZTBfaZus57ebH/TtOi
LPbBw/ilEoGVjZJSHoxJe3R/1l5PV+X3caJoWBLb96d7QkiDW9egQZOew/BO2Hsa
4ukGBud0ULJIVoiJWBvlhKTrCshz/1DEcJLLryEjtEog/tlyR4iNuJ1DvpwqM3Tk
Byc/PYvxj2hHXskNYpMHJJImmjMBz+nJxzFW9sZPX/VC+4UkMhutBViJZmTf95GI
wigZgiKgzoLTlYjohC3LuMPV4vre8DoP2SIeYtgn1/ZtS6NbY2rpJgOtWhONS2T9
rmlaAi0NHUFoi6LeNb4YUZB6qO4+XNyp0E2VZQUpb3jfBzkoQidSm4wgSQLBGJzF
ubv6S0oauSWa0JoofZzM6Pp/J73qz/7fwkIdxEQ5BOeCx5LT8FtYDx6McnW8rRUo
B1bSQ19b8gCQKiHx5okuLJijRCXW8CV+RY3VRTC3PLzY5h0xtkhSPO+xT8CIRWry
bl2z5upXn5xgJHm0ypUp3HnMATakTxiHEh7/tVY+bdf3ToiE2Qk+pmTGM5YA64Ql
Z0qrGW1mS9Be3y6rdlc7e4f5xtVAywsRKRuRb3EmwntufK1ERRk+qA9sDWiurRmz
Ndr5A+HdmCDGHIMgwn/u0fZv/i3qqkJWK/VE6/YpQdy/PJxy7Ft9ZPou9wicehkN
lZjmwGjV9eIUHIuTF/aUaGojpk0bcRWnR1HdrOa0QJSEX3TZJz8B8tT0kLDZdtyW
L/4B5erHzNUCmgzTOW4JdqsuLFF6aAwI2wcnLiIhQjByiopRGRYjiL4a7kr1K9s5
PclY/MIqlBwgk3DwkcCODVJk0oSyr9Rsue/vz5kB5/fB+qzCqM42wdVM3XEP5yrQ
x5s19cCVLu9SXk9V5zy3ODp0F+HuGQFiUIKt6QDOauWECHODZCV+crsaQUsHiD/n
tLm6YWP9VWgfQvtmdtrJtCNs5audqKYMS90mGmgRbvIBDH7T6sN++KjGIdZNnvu/
/pyzHPE0ZYRYk5qXwsUZ/fkg5rM/UOc1UN9MECiN4XqylqXCt2Hjng7Epz0opm5q
wITecfrvxiiOc1fsTQpfsL7tvgwRT/HPFrtc/LOUyfWOIz2xQBBDIMHditNXeEMy
ooSQccQi3VV/KRXeJc/TUBXN1bE8d/BiLY8RAjCY1n8JXX1rqYGBqHnBlPgTsF2e
tYewRB3+INX6Ih7insTdGctqKZrUW8BKFwNekB5Zddl3cYu9x7yIFRC7HEVE9r6Y
mArW2F6wB/x7BBtGum6NwZDBvgnEwQckQDFvJepbkWF78nlLWAdO9lamw5DAZF0M
xqvHOf90pbMKPgY5qTNtXiGvgqgxtWHylm9lc3V6WVbxOHzEGcFRhyp7lgTUsGnv
Kn3BaYZ3xg8GI3e/oPPnkPOXdd0GB4GWP45638UwedO+LdZHlpZufbGjmyHax3kM
/ocf2Ratms+J7xk3LYbkRr61KrhCsmCoHMVMMAiL6fi1ODvJwEoDoXeoHimVky8w
r/5JeypEMpdBiAaWi/KFsL8sjgsZvamCYaqY5GLLoOeyehl4A/W7N1ozbc2QCvy8
YTGxQG5NnmTjMZc945EV+2YC99/4k4mroKt6dE92UGwAuvPoghN4mEb4hO9PM6ov
C9SGmlnXyf72tISaGTLjDakhlXFtQQReIS29sWJCyr1oe29gqUd7DHy6jSWql6AO
Pa1NI9lgEPXHypwNcI+vCMk/drCq25aj9BwABTBDrGvOETiKjpFdCZtwf9GRHaYZ
aZtO73WO2dOiPb/51hOxnv74mh5TEZ9xij/vRy7IMvigT+1wKI03nQF/NhEVThfm
C+E+aFWgJafix1kaPYDVVsPNL7Nb9inFQnoZPWZdNUzIUxAAl3FRYdEq7Jc+gqI4
ROyvz4Q7vHs/t3DLeJXEI9AuwVLugo5hqYma7I2UKrycCOTbrMR9ZE35D8ReLJCP
4JZ0Yr9D+PELgvq2W3cj7CibluCV15J7knF0yGJ6YDPcwlQkdqXy8aOshM3gS67C
UVw+VoUnB5JgyY9NsWzaQyyj8ChPlaWgfGa6L9itraH76rJf/E8J0itZvZidjaeY
Bd/1BCa0vhB2BjsW5hU63lWsm5B2c3Z0WRjbVmkqYuA/0zv+sSa3WgN1SO8nK29f
B1fv0czStkdP6eR0YyauyziPOls+ovi+X2czT+SSybmHfKYHmuaRSlPZvrsYHCC5
5YrRblPA/v3SO6ZUlgBepw==
`pragma protect end_protected
