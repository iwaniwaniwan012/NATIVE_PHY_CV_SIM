`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
R4d8Nsjk4jzbn4O+HqfLMybRwzTqArRwbAfX0pVjVCrpELJhzFpEugITSSiN6sd5
VxGW5F9CShjaaeDDJoroZtUE74qOuC7x+JNWIgZzP7Hg/iIj+qUuEmgHVpnt6TS9
2jres3sBmjPct7YC5VdIUSfhqEOcaMFybPdhwOp+H3o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 34464)
C7wEFs7vrcu1pU0xh8NNsh7XF8WbwTQQJz9Pa2VUBoCSqZnRHlrlwMzhkU/mNh2d
YVqAoBhy+EQA91Lxw5tPydOXdRloptfajRHIEQJRcoE1hJnljqY36w7Vsbz7DECT
aeG4jc4Pgnt5vumbEST+jx5Xgr+stkGEQQwD4kWcq+RUprMjVqJCesqZKBdItyCR
gxxwLK/6wgnVUnLmQirWgKS89SIbmxUXW1AstylOR+rIY4pTG2T93swSXhFQ16oi
D/1QVaz4+71hGogxMtI88wE/Le7nHsFpVx4VZwTZeonq5Fd0gnzlCJdAftkEkQFM
GglEOVEGBA9KM8V5vWUv3eTF5Gjm92T3ETQ0TNGX3H85SoECyJgeXc6vWFLOv6dO
tUZwZkvSaQtQuj9WyUDl84OihAjvoULf11on3RH9FDswyYTMsTzkW8aDJBn/ygH0
/iXcLaWfegxZ1YzeR1TbtDOdWVFpmaFijND/Yn4d5V3D4vzjdj+O6b0Nvi2RLA/y
Vivuv6mDINjQU1RwS0ddMkTX5Xeqkzv2IfyJKhrcrlF5SeNkidCKCLQP+ZmkPc3W
Zpz6XnvKVCVmRRFw7mKKSM2Y3A9HVHW0FgdriJKn4KbNLoPkF6cEuRKaulbqjBw8
hgX1u6lbGCl9aAEWLHvzc5JjLPa2OH0e7HrpE72bzTzRGHUrj+0kxBr0X1tzrtus
62JkXUyP788CDEDinb9ArESg4k64tMGNC2XkfpwkgwwF0ITM81yuym+DQeGLQnu9
yyvWU7d4CwLl+/lfnxsgrBxhsrlHQN0eqr2ZjQ3P67JmJPLS9Z/D9pZel7JKrF8c
0RpcUrAP2QPQZsss51Q4iRfILH3Mh9UX6/FnIdeRLxZJdD1MPjpLheEB+95xzB5p
/JXa9+aMco81t+mLY16AtKWsg65Av6sdUL9bLN7AA/n+zFR1Xv0DHvNREMIihexa
uNs/Yo7jBLys8oSUe6SgfKTW+uhhbD6cbfbuxY+KMxwynu/0yg4plpwS4dMfck/v
9uW1Bfe1Hk9G3tAdQ3xXjcyWH/8Vc3IaTH3199nku7nbdnbdsaXywL909LbYuvR5
FAUBIZ0Xs66sUuiJPskjg70rK92tjwcwvDCA1e2wBw4gPh/TFGVehjQQNP2E7PrO
j/V7Wvo9G+yj3dFQ9JPu8qRX6/4kDxR0z/MCpng0JfOwnuaOSMUR+X8EssY63LCS
UGrkzswXaf72uj1L4dIWyE6M/MdV14a7oeRvqaoBt/rbtKE1GIN2P86lWr948uhv
45N45HzDlV+VL06j1ZzwAPkyrpLUJMRNYg0ysbQJdrEcP3fDOG+Wd8rJPAhEtUks
4ecFw2h1QpRiMdPojYKVXNO3zfXda4UvBrG3P5R5aeKxSmKGfexnnBKKvbvBx0iS
ezosAvbj2yuk+0CxPCeoJ1BSB4JnMD/VZkdauMCqT8zie2Gii6uQzeph3fNme9uB
n+QqCh4lvQRD8RYbobb568ZWg3Io+tS4QsFwtPNDBW4X4Q21BvUrf6S/sf97Pvq3
mxlL0KsFQPDyxOoVqlKPJt+30Drl6hrY53EmVgHez1ZADIJk93JDSK7lg7mBb2z5
v76Uh4sGlGFgLqJfNioiuM4prLEeC8HkXTcbAqxT70t5qPsmjqBbXkAtMlpHefg4
1uOR9e1m275pxCg++qwjlcWT6yxh1ba4l99tIGxI/LsKyQw0l/THxJ0yMqqRFGAO
C8yGndaIVWPSuERph/aKfA5LADzctgYybP7JuGo16rU0hgPxA96XGvgeVSJhipsu
0OtKJOkDBP+MCUPK/YvTyPLW/d2Dns49JAsm1DIGqJYgOWHYlnKIhVTc0Sn5jKZn
3YKmjHKBWieDKeBu4AgmFhLLO1b1KCpwDKgrA7eoTOfq2KzMi2afBgOLVUrpazEK
1ic6ehI4IhC24KFYbPWNmi1GfQEEVhUjtWHXRlSnoW64Tb0B70pmzH7m3kaYSFiw
6MZD7Xxz4Lz5Pbgo3BAH2YfhqA/yWHDwq3JKQiexwZlJ2xAqoxbQ0XxtCkkVPe6/
96YXBa/GD630SHHQ+kpAKsiSH4jhYYSl3LflsZh4LXP14z3BLRtFupQBb8ue5/3w
0vFGHVPdy2mx6DeA1UId6EMRAG+o59xFiJCDU1T4flSf6dHv828GpPcXYtVy2Eny
ir36mELbjFpV63ixI3IebwMJhmI9yhu8TTdteJVHSstmpdtLzqM2RnGNEU8EA3F8
7+TNt0VROChdK7fkL1rfeFyT8olXmxfzjQIlVbjHD4IeHrvnQSUgcZe0GlmaqeFw
RWff1fm5RLQIE4kIYhxMcq1YIjuLxpFeq8CuJbAQr8Ls5ewYuayXctH3KXZt1YsN
lHiIOMKD7yEgaLucIAyN38HbhQPFKI9zFXyI2IxQaG0vxIsUYyn806mQVD8wxX2Z
qcF5HWKpRYccnZdD4qh47OvytmyZp6oj/Ly1bNpPzj3FI4uQfX1LZ+ASjsjaKlho
q/g0FZnsGkDa+SCfbfOmq+dxCoCdDUYJ9k3DXlu0gCIYxIecG5FKfZCxOtdJCWlC
CPr7KKBIenGhSRUS8uo28T1ASmooE5e2NBQ5FIoagaYOUcBuBe60I3zyhVDD/soq
jY+gNTcRBu7arLAljTNQ3NSUlUesBsU/9ikf6g6kZYFCkE0puZP5AFwaEMyjdczN
0W50Ae9OO6a/lbXRS6GgvjBztAAA29mM01yOFAK52BYVJt0b8oan6nKmCH/dsvT+
P2HQFY+RhInIC3GaQQkjPnkRugkRQ5aGRttTDjk0cJGo2TeVEEbrx/0UYTLwSPdL
v7zp6oMgFP/mmmZMSRKc93dURzvZeSvVJ0wJBWEGoLvbKhuv6zIyc6OUhIaYUkP/
xZ2Jmw4I0NUmLB0y1J2OJFOK2ZDpHk3q0avF4mYAzR9zl5R9kK0DEgbYJOTuWHbh
4p7kaBP0jZnj22U0zIiBzVeb0HGYJEp6wuqRMbkMJ0MMbZOLo7uq+yM2NKxJ6EG/
VGPSYQ58iotoAjFnA1S3Qn7aHkHKdvh4pitD+L/vhXAwQGvkcBzcvScYqAqcMads
b+HkGpflepQSC5mr+uXnh5vTxIcxziJ7UZL84VIin04VSJpQX3Ka5/1uVoIIeBRe
MULBC/MH2MdInz7i+CcKZDk2p07Wy6fPgnCOakCZsYc3onfxnKniuovyzgEvM6KB
J4BF3do36ujRIUs0ZRfRsz3d7qMdQZTo9XAayD2lbNX+aC2pbLucE1RFBdxD+joe
Wusxng1g5Z1qJd7Kr9SN6LARAXAhgvtSBWM6KqKmtFsiRUbQVIT8V0gecDImkWMC
wc5wR8nSmhlBBr95OzOc/XeuF3T+CZTsyhiXOWa1qF8M4u2s30pVMmqBMGWX5F6D
qe+7nzresiL/UYrcTJFoa8gv+oS+60YiUDwM7/WlJxNLaQihBDYqKeCJD1kx0wc6
3TtFHy0J1XrfFrC3ZYzX7ON2kfrOgBWTjW7R9l7AjHmwmUMko8nKYRenKEYo6t4G
e+ir0wON2wDs5SKUCFeiJ6Qh8piPfdgm5tUBLRnivPcz92uLgEJnbvaemBWdYalE
A8CDSKUTP0MoYRdS65ipfxT5XGjN/8v32S/AZEEjCdRms6AlQ/7vitUFwnlt9KeR
+qQrCIfGhn+0YvTTehRVgp1zKwYW+iWlnrPxiC/+KbuFWL+O8G34p4KfhqvWgO/k
thSmWt7rGrjCmv1yU4E/BvtrRfUFnp5t568qZW0aRCAntCCNRePi0Muya3fdLLVV
YEmpRM8ypx7WGocFJ+5i3rncCZTgXMyHnMqqC12Hhjne6EO4e/G1VLmhAAMjPcub
mIeLZ7TOZ30XKP8tsW1e3Vhu0q1JGq1a2BZY3ZOzLWl8uieY+WWl7TJVmZOCGozr
Nox+7OIF2lSgDJ6zeB+JSfbZ+T+IGTi7TTSLveL4XhAF70gkZEXcabfB8+iCvN2v
gyNQYgQnfc2kgm/SzqCzch3xyiCuhjEfvR5yTtUOwiIKwtVn3qZdMM+9LDM7zWYW
pY5dvxzD/+ce058m0evpJlYY590rNTC8Up5BzK0hhhhvv5Gw54+O4tbDtNr69uEt
hgZerFXEsok5EFAx7VWcdggQfmbhzOgYGp679sXv0klJZlWeqOSdemMjY6dB2W8G
X5ZcTD2mEfyFPJLNBwPOh+q4x+dyKQDNCspIDDGkG/geTduQQ2nCxkIAbMpZ8IxE
VuYJBwQdxIHu3ig70+aZkOkeQocH5JEiU/whGodfk1eZDYZ1Re/Ia9wWOP6MsIDW
tM+6DZXOz+TWfsHM12zQKc5V1XIDyDyLELiOK4Sp0vZtpKL2qizf3QZpymnUM/di
JQ/jnC3fL3ksw4eYcRzAleTiZsUm5xpx0Oa2+w2MfxuIX1PPJ7OTCyqNT7yF4OFL
TJ2OmFdF0KLMEYcVw32Sol+4NYG2+Idct2l4Wx4IvEJInc7+PADCTtMKXupTYL2S
vx/t2BCnssnkY/R9NC/MO4PMCsogZrwuwebT0sxXc/cf5QmSHhNiSU5b1+SZhIut
0XipdTeSY0vsqZJbp5xBv1DggE7jVajHhgpeeTuChnC96iKft76qAnPM8PczPXxw
rc7NIbvNqJ79+Ozd8zVgOz1GfwmdDvo0Nc3wfN05fiDnwofNf3EGwTVpcbB5Mrvt
eoZh7f/UkkC0bpbV4R4+rJaP6aXe4jHQOHd0Z8B5I/H57CzSRlcz3bSHvCudGdFh
1eCB3FNkII5K0lmbvVwtXe0QdKePV/+2I3Bqvkes6a6c9veyXM1uUc8BUoyxDR4I
p7MGTEo/qxh8NgmRRLtCCAWjoh1a/VunoGlSV0qskQEg//lu3rwu2TmjsYBTVftZ
XNVaQk2K9j0pfiUl8diDZw6vcDBNRmae8/W4VXgCEqp4bf4Sm6G1o/2MmLyM4wrI
3M+K5XRH/OYlhOUOmzu5MjQLLy7LwvcMr0lrP4oPnDRg9wvFQrBVgJT1pcMLUIA/
0eGVOufvvrYtjeApB2qVOCqm24tAKMVVCW9Qxg224zBVzIHnTN+N+91X83725lNc
sDuaMn9jgYzuEaSra9xuDuBekKOK6V6DFVof6ArsNGEKaHB5rBQtYDpnBANiBoxq
9b2XaWhLR2zaU8hR5VdeKoqV4EBJayIUPRT7MEPC1N4jswEM+Kbc08ibl1iHR3u+
8WMjfcJvnoopQAE2tXOUdVjYqGMt34zo/3K8Fkeo7EBTpChMlN7g8K4gly9lAJGd
1xTerbC7X4cDjBlidRXFbOyilMUYjmU4Kez8cvyZkZ2jkyhT3AulO7kOw5kTz9bR
s3LSCXYJ79LRzjMefe7tIuBRjs79uZBJkZGfucQafmbmtoYUnK/xTeJUS2vI2wfo
TYRfmaflOSS5PAcVPhKfoc9NosuxsIFqqPptpRdZxsgKxsJXMvxEJOs+OAHIZ4vo
6Ag+hkVqpxRY7n5c7YdSQ84ZNcShRoTG7jYpvO+NCmOiMr8aOhSs1PMBvzS1lIQ+
D3PJ3Ztq64qdCtpjY1O+YWnZvoCu/m3Wm6WYAK44abYoukxitG0ChTnTfqW1IWlk
0RQ2Wq8+HSm4Ss4BChAed1q3K7ATk3W0ZvZGG2T0a5uUuOywc4HFqIXXoUnvbN1W
9bzaU9WGqd/sJKydFVNCN0M2jNJ9M3JCfNNCyn4AVpnFVBXm5LIu9/xOsCaRAbOW
OZgobbQbbO30OEXNejUxomdnhsvqx6/3cxffDoRnGSQ/CHc7VffaxzqIDAcxxLPG
W2semLMameAzEf5QOasC/gIi9mNdNiX2J2oOOiQfZRSDMRx8dvDn6aVyjMnot6SO
E9TGdRPIzhK0Z2T1kullf1VJjr+VbbRK7XOKTispwItWofMzdU+iL1Jn0L8IDRzT
GWSD98iXa4pyVEZnZeyfHFwpnfGLfGYFJv35glgBe0kaGNIzabPpxrEY/rm9HCsy
SgDh+74rn5oqNqaZTrL4M+C/6cVqcNAPFJaBjBfMqb0y8XgysnoCXMxtvsBmCUg+
GZMeuspzyC5+cIRVLRdVAV2/4I4K+ulpFurIB/5jxePEXaHs6dNtV7T6UpXqMlyH
KNzs17BQy3yIItaPpXKpw2HE5O5c1XEER3UaxaK2/AfuAURQdLXBnze9uB45ZwEu
Fzd1/9mNyeIdDBIMxb2ErqT4cTLFT7kcbfS8D9IzyZdb01EH14NBZEvJJOw5aRK0
OQ1k5RofRr0+xsu8yFnCm9+BNfbzmnDoZua81Ewc4Ot1lCIy/ZyG4gha9ydDtXTU
Jao3Sqf8vrghmban9zDtInSRttLhShvWEHHm51d3418T5418FXr2ZW/2Lv0ityYH
gc8V017Y/3BGljhOtfmnWL+nRL77a4aixWyYjC0wzQlO3cigYAkQgnZx3kYn+txY
6xBVWxwV0Z88jq02/yNKtzvrAK7r7FPIwSHFu3+HWC2ETNY/LAPiu1FqpCxEBMKG
xa3OkE6vyOBSWCdUDYkzw0eaV6lYMhnKYOYw5P0bohaOW1vnysVPA1yvBxv+7o75
8WsXH9XmyEWE2FexdaYeKYJDMlIm+v9ltL7Cl9DbtbEQmDnMzKD1qBJYj2YrxoEq
Hs1FB4N3RqATmMUAfNEPgEQMTBQkrsYTaQv7g0RI7Nscz6NAXqsNy2A8OjHOOxGM
/fl7fSQgAfgZMZpn2gVlSanroj3QYUDR9/HqrnqPi4dLTGQpk0PaA57Yq2J2CpJl
9SyQk6v9vgPLiE4xCBMO1Hdd2XIFtdvkNz4PF+26MkR+o+cn8+2pJITDVyw5K6sz
jzi4wGmu9CLWtfwwk4dEIaQz4IhA0QqIXj96SsKE/uzm8H0zrx6i2eEo1IOvu+I0
fiJ7tHdFYqrk43dDZAs9d7JvL+xCEhoFzhy50nbF01u/qddruQdqeycxbFdxYNC+
6Oc77ueIdaK8SZ4sskbugpkvARScIEsF7fuUBZb0Zr95OPgU0SkRWfdslf2sWxiH
aEsn6hy+eJEjtgO/QkjYuo3fEjGy717veJftRIItToizaDBZTDtlLKNMkpQbAYIe
golcP9tOELiARAUMMckKX69anjwj7GNSePu0doakUF2ans0pbgZtKWPnS8c+eMQF
Nq+bOzrDu9VRoK6nFzAMoYywN48JDMG12b+gHr8k6IuCZP+06Bj27jh12Zek+BaN
/zNKyD1dNKgIuGIwn+khWVlLVw516osL6f9jXsowMYghcb7RrRMinpZTtpxQSuG3
DhdYZo421HhUi9rjZjdu4dQlS+v3ZXXe4t1Z13K/mYn2maTJYvcFfJJ77k0wgY9f
Tc1zNU/MTqnZMAB594GKw9Wx+xh2ypK131RK2lk2d18hrd0NsG905/JBPvLaSx3s
l0mWfjY6Vp1ykmrt2z1MSjJ22wCP76askCDzVXmOZpeU17TqAl/F4y0gch+BAk+Y
TdhV1ZOi9oThRgWWE7bIpORGOWZggCyDjFDzyuGZWjDH1Yl/d+6I7nM76g3rfMZ7
TVw6AZSQxrUs3J6Ww7ztyl7rjmOc7EGtDg3e9RKNIOijU4XPQp9Cq2o2q7thCPzh
bm62fBZiJHX7et0bbbxfdQXCokwPBLoI8yn7KkTLWCXN72QmWWExOs5W6ZEPnpMI
Y8X9E1fA1Y6tmYgQxTgayhdzDPF1eIsEJdyyoqI+3w3H13b1qc5dLISFVEhanhG+
ihrX2MWIYBvwAwHI31xQXc6Ez+MI4u4n63t5ZNJ5KpqtZ1idGpwddra/kHxIniBs
bEZFSTarvsgn2d60Yvz/Ix9OfTZw1jstKetLTF52AB39mcRId9RtrswjJY4xyB2+
kr23gMCc2k6NDG2d7Jlw3t3KCBY5a9hVxxqJzOq42tQsNKcCDfujcUSB9hxnr02Z
SjLtnbRKm1Ry/ZV0ByOUPFOGMoprcisK2kmk5BmK76i1vFgmnU8rSPjYj37+DZXG
ypT1AJ2/yAgU1uBZOg2t5XbDNH63IdP8xRpR82opHnA1YA36fifu4rMw51esUaNU
u4MeP0yD0pPMK8reuv8zT3PdsYN2+Q5Fo4ylmZkNHkZmuWLeV66xillBmZMFlZAM
R6rF8ZNbAwtr5O8GRbqvT1dW4OTjxAokoJsI5RSBzXNT+KXo+CoL/0mhNpmnO4Xy
5rDT7f18mhHrpq4q7SGXZibNyQnFk7+MHGr778Tpvy3nVdvfDWKt/DWDDd37WXVm
HHlfbThMs8tyx8k5WfBgrdQYlN/4Yl/Uo8Kke8aJeyOWznm1z9zbGxJodw+P05Kn
BfaGLX7JcrX0ZcdMeRiSYftVg6a9wEl6fZSWoac/t5lLAzMNMXqXawNld1fhFlI8
lP+QvoAzMzSXj4C8GiR11BrZi8+6+VZQAfnFQq1eSFdRD5wJpPvuL2xGlK5GGN4r
KsyfSGoyn+KmjTH7FISy5+cHhAKBQQ/s/1te3xM9dI+EaWgUjQtuIuHakA9u1Cpj
Vqp9KYFuEYty69fgIZhdnYUOXgDbWpw8f8LQgMgPcCTl5pJr4IMrrYV7DT19tfSa
R3WVJbqCxHFqYKtjDwO0KfI2YBn0WJ7tMGChiNxDazQKo+U2vmjgY4GOPBISFidI
ghcP/txbt/tGJdE3BuE3JExCBVWBTBzuw1BgJP8sgLVAHC9HFfsyvIEg/sbWxFVr
/NW1TsdfgfIi+ixtAvkLrvfEUiYtAZMgOYg1mDbUDgZO35cKiz3MIrmOkTpRhzr7
BZ0ril+3O8FwrejSxhtDtOGzNY0e3W3TuV2ABiMrzHMcmQkhHIDxPajN1rr4BDSq
yUjPninzONtjJFUan8CEQknuhNJzLZrNM6FnpnXA9j/jrl5gd0m5ES9wnx2nmjuP
a6lkTNwkNE6jzW2E7XJx7/e4QvAhIbN81Ymx7fPhGaZXv/AfsxE/DUQAHQ8OKzpt
wjsfJ062ZKXThfQYT5Y5UYblTIrfvoQBi19aPMTiouCf/YEoV2aDcgmR6AGlW1fN
re00jhAlWJ6XqdYbZjGAM9OM+xsmuYk0+nUxH3s3uOM8gvQOo4LNG2XYuwcPR0eA
K60gDsX4sK7nR2jMapS2SE0H1Uyj+zr/pugOP6snx8Dkqu5DrIBhu/IY6ahzJ+MQ
1QPhO1nKUs3tvzw2sVnfKayLJMYKPukb3EcDccbU3PHX1vfCWVyw8cUEIMwWRNmg
GFlrnkNOR19Pp4I+0JYFWMpDFr+XKKdeRrG/TkItc/DPU+yH0tujPC9GvuQ7qKwZ
RL/c3Xm3blprPl02hIA8ujRrV8BL06VfBvtpI/4j9U1mmKyXXOL7mPY9J3CoHmvb
M7ZH8vZuAR7Y9Il9puepoRB/Djiqhqns4D2kNmEw6JdeT0Ow2dCZh6B/qbpQH+cT
AUNIt8NCcOrq4lwPVr+7iayqyggm3BfSp0ILslH5EFeYR6KObtuRU7sHkBWTphZi
XlMGfCzMGYY2pZpfP/tI2FNPJkbc9pXlnzPYKww2i5KQ7F0R3qulZ6Tvsbaq7EXC
veu9+3o87/npZJqHnfO/UCB3BfIg+CHtW0/ydT0nmaqzv2fvxXqZyNDyorF9jlda
EOK/bYrsoiqsi0n02bxWUSw+7dJgqz+WAwxluDj7qzbIpXl+Z5BaKiRruzPUeW36
4TR7aqbBRqvgW2Emo5XevQaYW8/GYBIJGl6+kPdy1z2yzm7ymktPZdeLUy6B2ybN
Ok/DifkxOysKWsoct6S7ToZEomU+9GmC7JW3FfkdQY10v6tT+lnziCkkd6yf/iQ+
YDmfSpM3tJ7UrO4K8SrFm7JVLKtLYPjtgq1aj/5+CbmbDp9DBMtxIZpRPW4tntXf
jPnls+vDdvAA1XLwdcKlvIwR6OFTKZpcO6bVeSBBQ5vk4q8Kn9Fk/ebP7YxjY+N6
G/8UbDkFg/M5fUU54PSj2aKEOuq8KEsga/12Y652mQg09hf93GQ4ZmPQzyoW9KXC
qye0kwcbLh2adf3W3E6UznaJvfTRRvD9Ky4+r0poQHrkAxepycQ+Kqdxekh33V5I
tQI7B0xvAgMZwBv6ZhhbCZsIqRNqAa11vABg2hbZSGPc+ZGtg2O1EaEt2Nupsb/a
AycdIYTCyRioAqJhod6uBBko0hrmjxImb3tXN7lc8vvtdqKGBJMIBlAP7g8Ke9cs
JULPZu75a4HBqab2zqHVM/OgtNJj0fRilkZNnod+L3swKbPEuHY+YKatTnFvPixN
V8Wv7hCOEoIPCk8vSgZ7u5gLwleQaX3+YlfsJzrSloazYPeF+P4gBmqsUuuIde9a
wQ/iLqBS0N4N4g9GmzAGFzYUCLosd+6U/sWVn2P0FCo1xE9GDnv6YY7KceqDOweo
qQadM4kw7lo0YbhkOgof9m29aDx88Dtlewpb9G3ydyBZKNOvGeqgyzl3x5e8Q0/A
TcH7nUZCM3YQPT7/foPbzu9KfDkuaE3Lu7AuDTU3cloUdVEV2MvSKiZtsWdXxWjk
u+Kp2E5BO4SKCePWfrUrZSXquaeWoznTuhVjlyhX5/1qfXn8EdxUXcsLBIYnmrt3
UfSWwJTMyKR/K+bGKOXLTFjJOHAEs2IuplYHMd8/rbXCMGcJgYnOaSNdHwQPbJDD
MxijiWWup8wttN2qD964868MqchFdlwOTmvNsp5pl4IjaQLFjBcsI3YQtAJlHpgh
978VhDNUIe/Yzfdp67/REC/J+oeuvwx0+iBpaBk5PVZGG5IhzMay0LuBh5YTYPPf
0CpGFgbzngkZVFpYTKNUN+xY/GpwJu5+wbdWZOLxkw44Qo5olOmAJ14bdPf5YIsX
Y8GcdZB0dcDVBjh+rCHBS0a1lF7sm/eCFeykHVMW6yI30fSZ5AbWMwxqEUbLvE+5
a7CHlRSj8rbNujQp6HlJIyWU0GM8Ef3o1HddZwHsqiEyKVC4QaKxhXfrDX93We4e
flGcFo+uZdNvnV38z3ULrmJYCxvr/wDbQH8pbNNkIKQPkEfgDoTBsq5SZ+YOABmH
DeURA2qMB3oZAG7dXxm/duCjp3hMk8qjmoEOahAdgIux8RSdQd0D82gNoish717c
v9FX2eYKL2NfaZ1yvewOUVLrsKF4ae/VHTTdT59qJ8TL9/tgxJkj060v/KJjsQWP
0gbUuGu/sv/l/oPYOi1sRCrzpxmH3ZcFZgF/BGdhJaf2sA2zVEWxNlIUv6+2U6fu
jcy0ExEN2RDih7wZK/o2mmr7JgwQgwVKHcGgUtoYMqJcjLjM7P9E4NZetHuXVs/R
Ivtp/VsJ3CXiXU5XO8NJN1NJolrzWN4Vji9hbg8RpibwD1PfQZNQCcD3Q2o4iM62
N03BCW9u3cwZQO1lcjO1UTfYjznmSGskGbXbwFD2xljHwzNjlA+nH33DfZHFKSvj
wetlaGJCKyaXvCBvnunIvjiQd8uSVuU7SJB8PTxETcIE7REyOLrcKEQ6nkiSSbDb
GA4sbxiDydFEk2AAdmkkz/ac0W5o6ZUCufOmThZWzhB2q4OKAfxQ8kpy8ok3Ax82
K5VxR+ewHoki6rRzCcBg3Z7zqNNo6og0QPoroa7BVjvbTuc8czF3qzy/W2Jak3Hs
i+CHey9GWJ7WDaXUW8Y0SL+Bm/9YzJPNpqh7Y/AjgfYU/td2xJ3npMOQ3nRzYEek
yN8wGyzTbd/mz7U6oQ5ws5cJ/4ZUHcXUn5MiIke1BK5fTU+2d6egs8zFObv4n8kK
13ifalhLccBxnjjDiq0XAIzlpMr+nrJB/fANrzaboVXnPI5LxvEAFXRRrR78NBkX
+KuJLqtaFilUXbQ5Yl+kBk2UOHhDL/DPAX4BsLPN6dxyb8PvXu/6/CCDAqygF6mj
WBcX6BpcKEEqzXSAEyXAwEltV6LbAFwuqMT6vfZkGYrfxec59MTb+F4iCw2iyQtd
EEqrnGjpgOL0EIwbBaXQ/G/e8p2tvXmmaUH/SzfpSYqV02vVEqXIndAX6sMWQuKa
HEgQQl75WlkDSF9almbtj5ZP25OY+5Dhb/WY4Zen6rqUOPx2Dcj5cpX5KQFJotLK
zVpnZDzzA9jEbEIyON5W7QAkRw0u6fqPCqAQ2eczn3R8lnZ5xBe5C92LaYDs5iFw
UYenqTpvYZ0aW9qo/Go/nQsGUEiiN2Ahthe7CjBUyuvSOO6mQIZCx7jq/376uUe8
sjiYMbcSZzk2HOjFAyUrF3EV5IRmX0TcxSddJR2jxrmDO1hWo689noIRGNwYL3+i
mQ9Sl+3r+Y+RBlcRDS4FWwKFKmUBtbakTeFXkJ6jTsBcSAWIvLe/rNl1zhlybKx6
3vTG8rCPGXp0U26hTQODde/TcDsYC0oA7t1AADxuH+0gGw5FzZlGz+wOJhj2MSxS
Dl5+TuBjrWaYbgk4xlJvibYGDctdvLviEctgkcVcK7gx8/fm/ZkNZSrkU0/ZaCCv
Y2BoCB0FNuPnvHEwzqtfsEi8b5+FQdnG3moTuHsr265df4qD3awxn3pAtIZKLWr5
4Ovi4cI0+wssmHPZLptR+mRZy64NqM1wM0gvn7BBCD6ytSs+gecbRx17UExynfDM
n7pDD+b7Onr/fClYaH0cazLpDGnRbV5NhI6tgoSk6I8j4okN0j6nLfTAWJBNdZ+u
Ijaa7F4iSuvZH78vGJ40YwxcrxOyZam/3rja8VFfYuetde9wE9eNKwqt3a3b3Tub
qgy3o25e55P60VClOlCa1DOqZPd+3zt1bQO1mWcikYdRxKx9tdx4/6U/aCx8s3ZT
LroJVi4Mx+y0Lb/7Yu1k86Pf3x9WpbbPL0R3r89MXmKZAjXwe0ZQlzYapcwBdU/l
GELqFjmZf1SKPbUfjljGGrfJDarE7WCwXIOFEVlwAtyFpnDcJmyuXO6dcIW+rbaw
BRmPOx44chA867MWpPNZGF4qCz4u5cPI1B14rHIh8R30tHo/q9TJZLPCSp63KmwK
xdzfTEvnMIto7u9p7oECHq7o+pFuS+BwkSPtHx9yibGrXN6YO8sGk+Cg2sVRhimg
0zx5q2PRlyJyGBQnzXXXgnxxnG/c1WPj2w0d8Y3HMJSVq1ClrLVX387UdLqT/gqC
d2KKSpG/QFS1RcsfoibsbpW2Q0JaQtT8hO+PGn2Zat8YlvsLZOVhAbtuQAKYifUW
EhuxptbF7Qs+MnDXtetNd+fsle4Xl5k9t6mebb9ilGbW151drJEx6HP1RfMF0eMQ
+54eO7cXvHG7dWUPwGLIuWU4tE4al9lj59itJYbxaXoyYtYtrT+PBezTjjsFuIvc
0vBW3y+tpy6k+Hiz+auwNFdLuSknWFwJnzmGcKGdXlVG4oN/UoCVIDvEr4jq6pcb
+fU4ABzSFF5QaA7DqHxU4AgTFmtg0eYGtc//ggPmcU4eY6Lu7DvCel9DEWH2UnmC
m147lZVnootJO8DCXj9ovHKu0g+QE8PWrDSU+Y46x/lcs1M2nY/DDe5Sekulu51S
k0uD1hW4pCU5vtsrHtLDhfsMED4JFZEhtHCMjscBUcjRuV1NQCcP1siZp6g5ca8l
1+Q6TnSl23dnsDNWSnbWx6lMnQFWO2tHkOR5dUfVUNYUnjwyp7iLRLlYFfGyu308
cLwys2hZZeQW6x4Q4xdQkN4EPFThodhtCm2kVqr1vlmlNwBm0yBqWLOWG6vwPDcW
JsMvq7wKzBhZPuNLHTjIE1fZRas2hMxo1b4W8gf8pIFGGF0nNW/cRJaCLLcmfuwX
VFttaXaAgz5OLyrmSYvxOjPoCnv4x+pzHLWbwu746XRzgRVzGnsO1Op1v1fYQUlt
E//7iRrPlKYy2qjE08rBvRVDgY85O4losINFnGXy677xCz+uHHAIyfLb9RlfzG/x
FpcB7EGIRAZ0kipstEzpO7VICd1tJ7TbvBYRok8+08J99IG+PPfl5IUslq4EDW5v
NiV8MpNwhN8t7OAD/C2sYFvANthcraMykTx00CuxzZd5kcqbR5OL359uXc/5VSPd
j7BfzHrLQ06qC22lW7stLfCJcvZe3hpHnn9YKYXMI/uMq6189/QHeZ/l4H5DSTAp
aVhv7bfgYCnkmRxvnn9L+IivsrKFOt2vbDpAj3oCfTl2UuCvfLuRPooIh8gPjpne
ABymru82oWXvvXyqni4XeTuYXaAX662bTDl4+KLFG5veqA19aRsGXuw9HoWV8e+t
jmk66oCMio/Z9yHm3l7UYUXwuEwVeE2Xbk/wyOWonNKD5pgfWZPbRz4OXroOoJA7
YajrJQ09pu4Ki1W1kmepZfLgn5lyWHZPfYNL+W2y+rssGv8DrEFDieybfvVwehB/
DiJD2o8CIktOP9FOifFoGCwZ5QBF18NpTr5Y1CAm3+4S86vk8M1zV+Izo4g24wT9
qqOO1HoZHNVRHIsK/x05HTLRUq69++mzWQrMoZHZno9mMSikn45/TdDDvUBRZsFN
NBu7KuVUBsxx/b61FGSMFeaj6v4qIN5BYKIz0DLEwus5b3f4ktpsO6M7I+moBnnw
uttacqp1BxjT3+nZs7YFhPBcZkpCNtezA6JP3MZK9epnGmEfKhScQW2uaGn/Zp5h
WL2h5MB06LV4uempBuaH6VLTlBmwise+2Vu5sr41OyQvzi12fdIkXwWXz7n8jO0K
vubWlkxURzHLU1+XQh9W99cQqceeGkKRvq7WnuoxUkPM42TQMvAQseDj9NyU3km6
Udo5piWd6ijoEQTrlCmK+m+lxS728gpKf4N761RrA61u4L+kdnB7UTnlT6VMBLSr
nBfAjOW2Vaxfy1oPmA2bst6pqs1Gwh50z/F8jJby0jpNuIjlpg7R4u7TeZqKWsEv
N2buJx6R8Gs6SCEWVS/5EkCYuCqhgPDxk32pj7+JKV3AI+y+wAnHpquGK2xuucOR
8l4+oDdxUjnZ0GUBuv/1lBkmHyPwq4zw+sd8BN7wlMGVLelG3idBAlyp36zxx7Z0
aAOnKUB7TwgACGrXNvvDHxADNqb0p6Hnsvd3tMy+MvYs56Z0hqQXtJ5FMRm8rqZC
+uvJuqtdTDAcghJ+TRMP+cWLtTZjxJSlyC0m9BQHHZFi9e2vhOAbQJut59dHAPDM
CQudiW/AbkOyEoXrnAbSWeRJLl+7LG7zRZM7/DpnK6a62OTNqmrYqTx9LNFPFfja
AEPX4yr0VXmrtrTn81+7YUqgpg496+8T3nXkqinVkVWL2FYl0Sfdp1ETwHniQePT
X3sW9i9dEdyXbWeaDrS1kf8f0Dfgm8bMC7iH5B0khd9tdmVcZut9CDTXdCBEe7LN
w8rvPgdpZc1FHnlazDQKljll4DTB5CZj1A3IE1vGYuWEw/S98DmTNusOI3lXsNdd
G4V69bb/bd8ez3qvxNug3MxswjS2gckoaKl5KVrI1stbsBrCU7qehU/ryX1goMFU
UghX7pCD6FNZZ/tzXTIdUtsyHQ7AemITdHinn4mPkxhG9AZDbKGgn/r0XP7reDE4
Acqcbow0gIRjgDVWW8UJIpWRiMbWcr/v/fok3o2rjtIXPeSjc16W3Gc2tJhAoM2q
hcpkrVmWt4SOVnAnQ5gp5j5dgqOcQSc5GCcV2SR931Fv5Etu7gM2JiB9Zo3yu5+q
UUxynk731UHogM2WBzb2cA7L3i0Mk+d55l9yYRnaLCoMpVs6jFgtr+kjzogvhgGw
vVnYPGF6jZ8iyAiijSicOQeFmP+N33HgZOPxVThjqJQX/6LCVAu7SJYWSHp7pRyQ
Ilj+IjrIbnbaa+/8E6o1g5R7+MQieAm2WMpmJ3OeyNGAEg+OmzvrN0U9UzVf93r7
xsN4Aw87YZj1PuA7HThzfrQDnkbWYbEQmFrIPmVLkUKHd8WFhkLi0/5N1mVB0ewh
vKRH3bUz6wOABdNI/AbK3x0+5xC7xQcK26FVaGHBk6fzFgxJYUgtk0ThGVit6hHU
WWuByRlVYmIX+VgjJoEm4cWmMopDlTw5gdrTBY10yKtGB5bRagdPcPUdNiL0WECN
eAbaPnzCMNJy2o4pv9KfROylwkOcw3gEEwF+MkM4Dw4/7iHz/7NKDe/z0afuFymr
dCeuDT55suZ3vhpAMK2TMHOwORmDbaQXnfLFctvrLv+P2EmzJLp3O7dEct5c4q32
qJ3Nzh0lGMCFW+vVWQ9Z7mDc7+mDFlw0VGBFlBCW2gNtn1KCMB3ETB0Lbj0Sju8D
K+WcuO29SFHIi21EQDgWMCLdULNzY3Affo+xWl0In3T6PGJUjgENC0hj4XlqjjEY
9oYDJf8mOeUbAchUARSYVUAwwUXagRqNSA7P73ubPCNs+klTdyoed9AmfT2Zr2My
rfuya4beQlwv8sStc7iPEwHheA86R90Pmrg2l+7GW+Nml10p8cop136LMjr/LJc3
tiTV6WrVHesh8CUa0XwAIbqI/9sTlBSETJsMahZqL34/SIDAQJfNxE0ftNT5FGhg
DtMgoG+ajDhV3igT5ayS7H9lrwfxMDiHLsgQNDLU0vK8xwS7xZv0aJg2E3crakbF
0v4ruMjrYs7z0c7lFBlS+sdagplKU9kNLWxlSk8+vkCdDgdQJoAKnZQxcI5LDxSP
2PHJ0sRzW8fj+uINJEv/qDZNlxnW8VkIS/7OiuzVhGH6XOb+CubuyTp0YPadBrgc
PKmukgK5NthXyeiLwRQ+JChK03PC1eJjF6LjNKC7HTEw8qAYEErGeuls+6msZP3v
iqdiDBCcZhqM29rYfol3Rda4PbOlWzOynuKvGQ9eJNkzT7qrZhCF+Eh0Ygz6UDhX
zDL0vnRX0NLw08DGkQmbuPBIWwb8Y7AucmCxEK9P52YSr7mHkI7d7C6zW7YVb1cP
Mmcb2kN/600FGUtcENA6fEL/B02lZL0AEfmipImnpGwr/Nb+/q87soVBn789q8kV
sBeFYIoai5tRpqFLfV/EAlLgPDLBn/SXoIWI8sI7877aLRYD+qEuTntpII4K7Nxi
EuQzuhKdkEzRZNmbSMyvIDHXhkAXpFOKnLw8UiaWMLlg8PG6hPIF8gJx1dGpqRjr
0bKl0sgycFFNvMQ0xcEv+1Y9RO6rblDWl0Z/wnacXq5EioZnphignn/IgTQJlEJc
U3lUoT55f+uqdb6BLWTCuWRidKwW/hOLZkWxwuTYSVQ72qMErjlHvki4Usg8P3w3
T3bUP4GLjJF6FXBSacr7r8wQ/N7mCqEAy6Gv07TmeQxkQJLpQZCLxDjgKokan9Qs
JV51TUWS8PrShOAgUZqzjAPL0WqmthLdxwQRNAtbyMLcAZOktE5fSTvx4dEoyK95
IXDkAOommvKAWjYA13vZSf1Az2PNFzooPLII1VlYyVUTqzD0j1xkNV11xIhDFGdy
inLG+w7pXqWWn7vDZd1+H+iSTP0UX61eLxr82Ud58idDJkmHVgsLl/7LVY/HaA4o
BoETkAeXIfuyCE3wrbo0o8UcZLvjmsSQHX95Y4FeV6u81Mlqazai73DFAUd8OI2o
OuiMbgqBYVj5K4C9BnD8wTWQDym9n61qxfyji0uYR5I8pvs9lSvza6PMNRAfyqnT
nX8K5zO1IdTliPBOc9p0OdFiNs6+BWaMeRUpan5U4mHnpbSVQk3A8ZRccIhGHamQ
RKM1k5f/fo2ZKOvG+Joj7H9eD0S6M6oMwUcOIzi8OnH4F9bLWa6UNZDB0JEzoRMU
OYuNlEhQWZIowV1P/7LWyswvluA2+RZg3lfbUUNHb2NyBQmRDB2sr1hgOQLlsAGs
QJubjrfQoFRcTsdlge47LRbYutYW7gqiMBk6hZF8MkNoe5WOdQTI1vwoSIoQKLVg
R7QCzIbSSRMOhxZUXaGp68DHFyx7hSEzZVFq0Ymt5ffYqLWerJnw8hB6YH4P0ML5
vdhUaeZA1zTBkF31LuUvoMpRAkWlCUOOGEfXpl9zS9As9FTwcmkzzrzFON7eQ28f
dY5xvN+ITY+OTkhYmSW6Io98idcFG5ezunlLw9mOLS1ofDr0qhXHXEebruAxZ1/U
1DWtMl/WpIEvDxcFWLnL0KajJ/OtNNeAFg7NpwmAhHnOIIGm4/GF337LFgofjRWn
vlW01MW9ddCEF2FV6FrAC1FXIvTpa7VEl5s6YmMTn6PnZIGafh9vjH8jhvQ8WLwz
4ZVgsnw2LQuuRTcfItXE+KI2Gt2tHRr4scaIOBfXF0exd/3gTcuHqU1mN8v3NRRE
ajGQrAavGnwXunHKypVli/yQgiMP8kG7y+qEifUVwe5E2u/Z5Jn7+lVBcobToK8Q
2mbyxhMn+qAWQAk8wtPTVWeaWOP0Ij1IKvqU+b3tH4z27ziobnznrUGUD6ki+4+x
4Z6u+zDfsXnkQ0X2dt5gvv/ayuY17kMj9HMKjx6raaOgVEABeQfqV8+BVTBRFRlT
S88XEMg6A5em3ZHp/XWHaLXk7JqBOPdgLVklRG5J/6V6MfrMVHYyS4YaYMnsCYFE
h8KEIzEmi2X0Vmp5xV9R10GD6fovcl/avedo7Nnai25zudpORM4SBeabgw0CA4ol
PEZUeTJ3/1lqj41F2JG/uNZKjkkBosWcUDCsxBGGmdlT+nChwFHXin26IIqEdSmh
vffR8hI+25eiofBH4AGISoTHK3wi+SW2pwgI7rqdkQTxTQsI0wlLRNbMyc6AXwKR
jVtDt4jcE4aZFxBycK3zLl60zOZyblcpdL0/5Cb1UJhNIwHVlyruLZ235Ga/fA7L
GPoPUeASTAq3M7Ci/eSe+jL227w4shceWuI0GSge3HC2zPS4VoBB5JWWKuNRJnjC
7bDtwB+3MygB/7tk5YKoV33i4YBIAABAINVI9P/EwTbRoGxKhQgkHpVkCri6ZrMU
rTMgVhUYNwc8iuEtwdZh635fzqQCB2sQxzRcNueWU9yS2zRq4+YME6nnTmLxpumB
fnvK2VLqlf5zHUsV0diYGxXX2dmEQX1yO4v33mAlP4NrxjVCr2VyptPrp5QKpco/
tE3VNpuaD+roCSvZNI20P/Sir6sTHHaj1uAiD9okm11QTfW7QD7ZuWXQh2tVn72a
oAclaXlXQp/ZpvIo35El9Px6joTpnE6vTbcTgRHGpW+IqfuiL95dUFXYCwWSZt75
DIQq2n8R3LFicaj94qI80Ubmm58VSXywLBIAUgzuQXWY3I4NNSHB7B3QTLqXZYDm
jUp/RWyFdrXNLUQrNvlo8bT8lTfKA27O/gzcP32qGXZcWuzO0/jueOZQI+IwxV0T
KmaYKbhkuQL4oLWnyIpSq5nlp+Quay5j2XxbzZkrW8wE37HuWjBAX9nXK7gv+R7p
rPMJKjikNBzpuQCQ8Hi6N3bBi1NJLqk2Wei7ccNwgXbdmwM9A+kQ71D7TU53QfJK
ASJsu19w4EkqZodYHXxMAYkQN2z9fF8X+r+50CNfsRp3IlZ8Yl4hICoJyZAidKZk
o/0Eq6Hl20zhshHhyq3s1sCSYEuGNnLxYQ7TMx9rykmrYKGAlB3ZLU2fHAkZDfQN
GthqxSzWi0RfiNhgHW0jGVObpWzN+41KlDEjVhToaiMWm23JVm5P1ingsgSfS1oS
LVDbaX/g/ldIi6kul5Wx5mycOMOV8OzhxKnF2GP2QHlofHEjiE0p3fhZ1VeDzMHs
GibUjbTWmy4BziyEAKsuH9YwA1LSJhB1pvWN98RvxUEUKJ+GUWahOoTSlcPP4fPA
ehNWkRHfGHXzxCCyvOQ2dVy7v9scWZ/32A3CZEDBVzbhXo+YAC1Og6es8NPTGFkr
UN7y5a0a4hR0BxxmpA9oQIiCr/4sQ4q9wAICnCQR/kNCCWLUKCJVtZcJnee6aJ5P
FdZplU1Pwh/HH1UbzyF+2Ale01S+mrytUad4nAjdabCGuQnOyLRPoAyuVfqvBPjh
zAidsPT7QkN/FIaqivrpywxgET9aAzw3BTIdFZ9QQntEpTozk+OLeBc3D9QsonbG
3asqL3qM6F6HkEhtc5TZieNVCydsq9hvfHEaoZWMx6PyO/6GTsQiZYvpmi4eQmBf
UMuNZnZHANiq59kTpj7lNkHnkCFCw1r9BNU4mzGMdU52qv3jKdvMj4od6iDjAuvY
j49AbTfNedeFZOxGzT9sY6TmSFeqAzTef2aQ5der1DLb269vm4NLhtAewhVfgX7X
LWMzEZd2dHBjd6WUKJELuTWkjl7F4ngUkI+XcIoxgUKc67uTpNchDf6DgYwNONdW
/jk/1zBRhzSiCv+PwWApOhl4DreVs+hrFiuzhfk/gqeOEyNNUTvWMJgYRdobYxqI
LQ9U/s6EXjooi9jWBj4O+b5lcg7l3vjcVuFCGidX8WeHrZirfx3BjbdPwQcR85Jp
PG71cw9GVXfws4VoLOb035FZcmpVBmJbpkLEqlTaDgwN7ciKkh/Aat/ZfMgKQYjj
U7l6ICsGCfEb6c2C5wIGxJ3qnbY+MVXbl9OT6axJ+BI5CcqMJCYRIpY7q7Q7Q/0o
CPu/U1G54vryFVw6EnfGL5Qw+NnMcQOaOkX0A3MHmj8CsRt4fqI+pJkF4PTD+0mK
Qv2F88qXhF+X0Lnu/4dWhtz9I83Sfztw2IZKpDZy26FRsw1loj2Q2qTUW6fckWap
UwcF4p0ejUvwseoLtW+wudARdAUMNaxTYxElG+a4fT/0VLr7nDiDetHScEBUiVOC
gMae7oJR0HTfFG8zqxgN50/60Ju4yvwpf6hl8OWTiE3oNmFSi39+QthhWXohol6Y
++Tz856JmPMCYgd/hCSnQERU3M3K9I72e00a0kbvsZUXDloYEtyBf+OiEQsDK5ce
JiiR9IAuwKW2teDYlicDLkawVJCLhlSF+ZrTtwHe72KCu9TYXihnqJPrbgvE/BuR
6rU3Q09K8jPufyvGvQejPRGAE+1uIsSP730X/bTvCyYEQ5EAqwgc+dfjwX16JrZC
ZE5AM/EEgx3XWKXiEmw0g0YZ05YWVIIy1+2CpLV5T0IZ+MqYbZuydKqKhTyLE8vF
5mhNrdGRGmp9lpX1AA5b/fctp5oskiUgNy11XKbq8r8RXp24TetaRwgiohZzBG6s
bofhs3J9xXlSx20US6gZWU4zFPyrzwbQYvLZfzLp+Sxc9grVa5LQPotqqrNWEB5p
4tR7fh89ZanXPxVDl7QSuFiltNxjqIorm2bBAoB4cc4S4uwAxQVwnzNaJ22zM8tZ
kJw2vUG6wKDJlcVxlPqvJnxKKwJb3aVtEFeCrGoszLvdk/HI5Ckqbz9TbPNr9+y0
/J+X+i6mTJX0K4ts/G7ys2lBP99ptXYEuOQf8Oe6l2F3bALMmBUyJffn/y+4yhuK
VKsYaP9ZWFjP+TtTkDaEnPp3ERJEsXb8exyXcNPFcuEwzxNTNxvGGSiiBio9g7B9
FBYJy3NDSycVLo33dyf07eGTzRij8qcJH3cLD+srXdneferDj/Lh+HmOUyw7rhYy
xsp2/bX4y6i4bNJzR35j/u6jxDgcYN+qfSmAqy0nzPyJ/obxf672HoNK/bLpEF75
i2fOfzTT4golR6MktBtMhSPPqWM8BiXQuUbB6g/fsWEvvBVbN5iwxTsp7PP1hrJ8
H4T8oZUm3CS7Gdq7ruDAsghH5uuU/4bcKbtjleLLg5sogHKal9WI8CRVrcSvxpkU
6Y39X2+jKMA2JDV9ujaYGVCE9j9DRtFKe1NHtWhvYw2Dsi/KDcB3a87Ue/HFBdvE
Hum+ukBNNLt2ItzqgH+2paFIDQJTsEq0v14Sk17P/d6zKjXk9WfjrTdwJgUC1wGw
AzhAKhAsU8f8B4iPhkrwBHA6nE37joIs/evq8F6zH1hsz8J0QGSi3K351w6WB3xQ
WRA4RQqkxcJZOeVf9SlWfYw+TBQi4tr7XMupJZ/MCDUMGq9ANoKQ/hJUAaUm9xBG
n9gy6RYcH3+42m464euylnJ+VvbDC8uOWhCOyKwqITd5hxur3cdzE1YDOkeFILqY
q/w8aTVaORRtgYON6CGt4twj8Rv3bvg/r//7E7gVZzIr3fbeKhZ4Gycs0fYQ876E
Bkruy3Q594TAG3zcW1eNWvju3g2UkIvJZ5hWb7aXHJScIrvCDqS0m54QQXXrzUDG
hXUlaxSUKezxnSK2ZE2J1d8H47mIO6JcO8B5Iel+F8DuF6f1XU4sPiOZ2qJsyYEr
rqv0MBXqVvQ5MuCwB97x4Dnjgy80pC06sGmnnprt2vsbk+PSvQbVgDc308nVvhKS
vPsmKOM4EfH9J4Hpngm4TfyY9uv870FZuBd7UgjJTLByD/N8s8OpL6up7HNOmysX
kufxuMmxchpddT+RB/zKe/3FCyKL69wlaXnN53JD1wflVoYfRgRrX4tFKPtBQwFX
RzpkOmutj5lgths5h8TveEosR9hy3ROotUCQDFyJQbTv6Vqe+mnNV1VYAWYr1xUn
nNOXwzKEJWO/Kkhu+MpRfAKemuHEGouBxOFSVrEsqI9oPfSWSEKI/vGOFoe+rvR8
DxUGqSRKo6t8pHHR+52ZLHmVCIo2veV0SywmQl3BJfjUAAEHYrLDFkB0Q6fCQrKG
fE9Y5OnpWpdLNAq3c7Faexveyc8D5Zcxtt4zWMmXA8fGE4gt0l1tOYtvwJlnMfaR
GtSqPRLnB/dA8ZWBJrCYY1+gilzd1Ws5adJhGBY4SmiKj8J/aAPP4ZeeSBjBicI4
gyyM6BDhX0StcaU8YxqYVtyTr5N0iA0HHhoEPryrVl/gxwO05UG1xLjhjGBS4a7/
ks9LMXOP/lqZbzwbBjYvGKRPBiI+0C4iuKgqSaMJ3fuyGRTXSya//+D8s55eMR35
Gda6gI5gzujq0htxZZ/fET6InF2E2ZanfeZlgEFf3qz2C/69kAZhFcnleJT1GZYz
yNg6MMMhacTfL0Xr+Ys+0lenk8i5MmW31yZiEnj0xjy3YZlEcLctOqrUr3ABtO3r
fNGXb7w4nIzIpSILZySru81ZbVt2vd1wiuobEYtaJ0qNOvsMIEPOHxEi57bVVX/C
81KA6S/yubBDpp9MmjX/VLksvEBrLRqft4cmSZEbUalpRqPc/wPFQpX8KgXCFTkJ
SF2uAmvN4Usy9lrKoSgJ0itL3moI52Diys5YqqIfy0+fRu7F5idQEwbdq/HEDoHW
vV0Q+VixDCUWj1Qks4r66LM4N7HV93V4HA6q0+itGgEiCixfOFlrAN1imXIOgFlq
UUJWn5H0FbOaZC7WO11kFAFZP0BgViYm5VzmS4oCej30E7ehxjExLrQ8yzppBS12
T1wcYFzNpQb6L1EEfhZGQvgMnhmPgLUjG1/kchAH+LTrVGsjW+qtfl7tLoML3318
bldN+0wwCy2LrFeD+o+jK9Khc2+0jpC+LsVKrxESvLmN+KwmtkB0WTcuCcLsvopx
oJe9lWzdefHkDeDCnbnAJGbxzcvaWoxgWg0X8sYvQN83oHNlmsVs95j7g3FQW6gh
PomEmk5IFMlUYv1VqA7Pjb5uWU0DU1GOvl4q+oRFhXLUoPpsiZ7bkFn8Zw4Hdlo7
MJ7jhIZuSR+sDezjuxVbAAHlTzjZFOtdQPGRKl3Zzch8KN7X13H6+81HTl5F8OqQ
6XIzgt6RjJQwo8Uh33cOPvhf+MQEiknBshtoy0gS7zTD6fFaeG8+VrxalIvf2VUy
FmlxB66zr5uk0hbpvZnIo7h3v1evZsB3bSO6mrrQtzfVg7BSe1LGc5jMlejGnzHS
j4tl0csiRN6sIr5FsG6YgSypmCPx7EQts/m8PKq16EmzZsrrImuLGJTGwgZDYLBS
6I2lcW9Hc1Ob4RpVFIbi8nUsHrG/9EQnY+ib6AhudN+xTY2BnX9t5dWSE0nPxZK2
w08hPeYPHGW3twSbznYfLeu/fsyGqsnZPY6eWi6bOvzR2LzsLeMNBq4zr2O/WadS
+qBAGmkRFWRnItgbSDJhFO9IE4SCPbx3UdLcn9mF72yWEPJ4LRz9E0qSsX0jNAia
AWsW40wHKfUUFxUrTYRvDqpFVbUp3trhR8z9NQnKFjLEVQD6/U24WUa064FtROO7
wUtoGjKm4Kl8gf/D7LmuyckDDhOaDta0MXuhSOvOooaV8vQoXCRggs/JGwPcyqdt
8SiosHx7UD4G+pjagi/HDPSzvyBRTuQr/3DV24Ix4rPSAty/y0Vs8f5Jfw6x0mCV
VR/VYkDNRkE5NJmcEKFr2yVQU593C+6o4p3w/eqbnPxjpTe3jOJdhjK1UPbGM9R8
AZgXrA4gFkncnxGSaMt6Wo7jA//CrLESuw9nIsSz/lX1g8R7/6Qm5tb4iZz0lYaD
U5RKGSEWNAul8v0OPkjPSR/jixuJWDCe8oZn0u+FRjEj9dHfOpuqJOY6W+E6MjmE
rd2hLUvm2XLxtFkUjLaFGZKpHwz8dJCNJbrQ7b5KQULs1ZKOU7w4g41Gs0MKWK12
LXVftA1B2/q4Vd70SNm63GVXp5svMLjF/I/rnx+WDQtQP9UcN05jLYwsqlVe1AaK
fhbd3iGRH4lp42pBu5xpR0JyfDjPZQ88Xm9pqneEaVK16AdNPNZzLb2e8rXVgaBm
680OHitT8OjIXBQPky2jyYF5LGQdtCxuQw8tN1VHfUqnt4/nmdsRjiHt1pKKYxmU
x+zbuJOCj3P5Q0xYuHueEGZhD2cbVxGKGubJ5Tq6G1HhItgWKmzeQN2LQ5Ia2yAg
Gle/2B1gIbePpSaYgHgby2hhkoOHkg2S0k4I3WvvCKjpCjF6Od4cW37g/mbQ9/L4
W9aqlmBvWMs5LoIV0l2slWBBg0Z94flxpoSPj7sZn55XisM8JXLsUJnBIGhYWdPw
8rKjRVnqlkDD/Dg2Emgx7lGDxhZLdMLE12hgbMBKUSiQa40NHUsrmEAFnWdILg4f
rh6EmG6dVPIxawgH0VqHBF3DOIDtwZfR4SHFXBZ9Sp5PIEm35g9jisIJ9pDCAjWc
eucgcV9gIe2pVyOBQvOr6g+cBDARBvVa1QXRy8Q+WX/mZ7JtRz6FELwak8JqaINJ
wFjdVBjQ70P4EmEUgEzaoLdoqdfLqowK0UuIi0+woiHrfWpGdKoQ2md1VBJ8vmY/
MF0brxo7lDBegCNE5RoYVhrPkfAVY7S5ehB33tnMcgv9HOqTvTG9sc1C+cKcelLA
NuM2Od5vKqkmF33pHfrYZToMcTWEL+WkqGcdIjwM6LMU/BHKanKlmYU/y4mi2Q1I
lr3tLrdXeUqVEQwHhmxmDa/YAAOZ8MTvtn+QwGRc57+OpfFcLnanSqbCEHIIk3v2
2SDwMtNUoFR/caWmrOUbGY8vMYJjlmK1eVrlXhTqZLqBL2hB/RbS1W2odmK5P4jO
Pe+ZQ/PmquBLDFSna5IgNJpyxy6qX5dRAqy7QSJirAnCMpkw0Wp8K8mCGIc1Lb4N
6oIRk2ajc272fNnec1+Do0FezZScchbabLp5gIf7HLqF1K5ctJJy5yMUTIeIEeSO
y72VNRIn/WBOOSSANNKX5IpI59CAKD3Kp+MA2cp+ExK4gRxa3OinMvZ698jaHUDO
9uIXZPCUIak9b2dGdVLJb66I3RZfat5+GcyvmdgHprDbF1sI6XOtLbYofCPsqdsM
FrSagtlkwjRmkiR6f0e1zyoS9MOJlVnNaRtQOtQv08KkO2bBKD/Amb/OCvFsRBNP
6vqU58OyvUVy20nS+/3ka61z7W6J0Px0ntFc4Vk7UiRpmJloV97ZeteljtyHRXmI
BS0r0kb+YQ45PrfloP2+7UFruG6I5NTIhUOWsRMeIEb+U8AoOPKGssXztMqoQ1tu
4i6OqYnwpCxmgfsjO/wj417j5KSXqpZTrz8ADMKRFohzG2DziiqNE/Aj20jsXFjf
bkrc/OBqAKrnu16VZIeZ8pU06JCnjEg5C7otNXewAQfPtHZ5tCYvm3nGf08njXCF
MwP3cunATS/i/X3k9iI9H9wH5yZ/XgsRUuIzw38Zsxe23E+utt2Q6oANei1lxtES
b4OBxNOtucbZs5BCf0fWjRSRh7sBXTXRpIWWlTpbKfWDwTzifLN9RH4J0XnaBqYi
Eg5CK0qFpvy5y/N//8W7rFE1fVW4AMdrWrtRoaLO/cpZ73Zv2Gz3I7LpuDKlXL+V
LMOBzJnRs9VeS50sGUSo+FrmcX6hUwcyqsnehgCih+ZYz9PXJevR34NdCKumc6q5
vrYrOEAGtbKbVHkEcwYFjP8UtNUSdA91nNPcLyLQKv8F2jdopdZ3O4thveIGZVp9
EtBGQbK20h2HtUhRAYJvm2joe7G03EznNik91WDo4X5bhe3drFD3H3vI2HFxj7HK
vwtRctVYowCifbFozBjyuwFa1HeZt/qO75VQENKcehR/ecFmmogXoJGj00nJJxCx
qY6/gEPv12ulRweutoFo2/Lp6gYk+GAKi94NEpLTnaKzYa+C9EAIyGefuTrfusQO
wrP8ydJZyEIcTf9qMgbEfSSzt6dI1jtVbFQ+3/jI0hF3NMrRtLsjetQijRKC6UI3
6NreuYTiMCxmQdroepFwQe3Bn1Ixf9erG2n+j7yNeEYW1FvySw/0jb+TuVoMOz3T
EhO3rOBzSg/CQtQXe+EvtNgrrWLhm7/bY6/2KpfASTvjrzzv6+NF8hpQDzgzcxQK
IZYnj/Dgx5izf/rBwDmP0hNua2ZNbgGKcTDnJaWihJThc9B0WSgElL1IiZPH1Zy2
H7smLUdKtvKutAuVdaW9JUxUxqxjm4/wiZRytLmrVET9jjpJU0sYF8TxeKtX2msp
1sRv/WdFuAa8/ljZh7yYN1cQd1VzvhajvsiZArdYSkaLh7MSTA3dYNtsyzYPZWZi
zIM0oTH7d34ME0b2OTt4LKPPKTwA5JzhZLGrDLlaqZc9YAwhSI1PweRiN6WwGbCe
5xvWzcd8c9FG51ZenPrkIAMCTXA28zfvPIdQ3vY21lpCUy8GznDgCR3EYN1ik6B1
pN5P9j8DM5mGdcxTNntRyanTQx190/r3MCADkZrx6vzQ/tDwvk6VkotpCcB3nf13
UM8MoeTtY2mOJYmcsoZry3YR43IxqlKChN64K6ojo9yl4vA3CfMZriaRt0SJnIt7
UdbnV3WwPQDtuAtdrRcMgZgNknMjFGnBOM2oO8Fhbd+2JjiWuSXr0qrxh+lFz/lU
QnXRUoG7TMmupzK/+OeINgbVZRsNLXVU+7oxfiQHqc3J21JCE6UOb9vSnnfj1k9e
dfu7kwyxEj9t4aBd9pc+P+dtym+5KoU8tgKcUl1sfj7G2TmWBBneWf3QUfsV5Xd0
3kFLiqIUP5e5HWVdj4Qfkrk9Nnqfji8cB8V9dYGvquZf9YX2jgqCY45JI95dTm8j
kPdOgTYVb96zrz6AXodKSrCE41s/AspF2QBXGhndwChksuwpgtW4m6D4bLb/vvf8
NHLoyU4+ihsCX3z4N551uIPzQajDgYDUHFErKez0eZLf1lXXtvTqn+JKKKZRD2la
YsArvVWLmZwrY7uqO6BFDFqk/nk+7rdHcwjpS8PtGZzqx1G8SFPOhZJHSXp6uF3Y
MAuDyfKziiN+YXpOtaf3uHxoHbD1XFaeZJlO9NLpuAuc2z6OIKorzM2NJSKIuWer
Kj33f8jIhdT1/z13Q6oAMFfZu+D4VCOQEbASU3qXN9zDXjqjo4Lkn/spstu1G0rJ
v7+dRF8E9DzhGXJgr1Ory+4QzQbUeCtvVOjQ/BrxLwoidPysTKxk3JCzrbIkEJsd
Da4D4/Zm1dMIjE92OmJn/RAauK7WY1QUh3Q4Qa9xpW9/Q8woN30AVcDNwzrdXvpX
5Rc9qln0MQ+fX7AArGych6npLlqe3FnM4Qyh9ShW6gffuLktupbmBVskUhx2x37U
G4MWKYSAj0pOn85CRUzplfBfDSw4BfAKa+0Vvl9xN0CDJxk49+F5o88L/01vcD1q
p7j5Ic4JvLEa/sYtIzBoTG+S93k++mXwbst7jtw08OetaRc7zo5T5Aqe8iepGKKp
7vXW8xT+uG0TtKuw038Cknt6OXemdNew3ZzucBC/5CcdyN43WkgEViEpmYyWSbpG
uloILcNDAw5xxygPxDIcUNSA6WxDzQcAnFDzo8kO8IrpgGMPMDteG2igZQM+nSEO
d69CqmbWRJKvX4eIJRAL1Cr1NuB3WH+Flf5SGKuqNJRczVlynPNir/FGa3H1/gNZ
B/O2XGRMIOLr4ng0gueHkXbc2Fq1wZ8NMlRaW+wCLLqSi5vrVPrihIeCZWVb2Jom
jEiLe0KscRurB9+E5wY0qL3eJ94aVviDO7ghcF5GoQ2fACAgdQHqQfPys4JmPGuD
lSTg4OdT5hWg3a05So/Bh7nkufMhtUocv+r3r9L7IAW1n4AkmpHR365dULa253cI
AqDxDa1aj3aWA4iHS3ibCN2CETBZ8Qd6ZEePmJcvpblAno0MX0wS0IfU7qePNSrq
TPRJSM5qsIfgO0GzuYu73Z6OPWEBPe7QAdn1Ap3uFNI8zssBKlmkkfcyq1rKA5ij
h4FEmGkXSq9JjkfqP32ODCNMVBLDb/dSW9o5tB58keGpeuvEfg4e20yRmz298Krz
w2rg0DV1qE8Pk1oz/bmFqLwGoHaQwEZWY7dHMbYsFNgcRQN+reXn6XXHJ4zXZFs3
JL3PHUHnTyzDvsqSy1+GprbZ+eC8sD5x9dFST18iQSgTRTIZHg6eXpT1YGFRkR6s
7e2Jx+JboE0T9Zr8V0YMQ7VhVbazphFNC4MP/YBJLBDRYR9hkJm3ZUZFVE99Kw+/
jpBfqO22J3IFDASCd++jNmbYyYi6ANpGP8nokyAaMnqKGduPNL0Qb8Td8yp6Q5h9
Dz9crdR3ECzvpIFPdn+wXizMwfHZWK82KF6b97k8hCounGQn1g7MUAIsqppOpayW
JwTEvM9v5zxDBUnN+T9yzT4ux2eFUVb+QCaXdsxqZeuDwyuiKuc3rc9k1eCZoyXq
G5QuhJhM1QZFMVQuwyL+JkPNw1bIEgWSIrqRVPAIehO7esWIxWvDTaltUAuyFlCI
1/jyEDwrdJ24IknpX2oJam1qSByfIPnzYznHSvbKpVQjL/4i9GWjOBXeh+Wh9xKe
x3B5ATab8MOl7/pg/in74V4BfdpkbLbvlbK/Rw6LmB0Z8iMoMtd50VekkfYnwA7X
ioYni9oYMv/kKA+H1XY5fkRRFbc9qVpvK4bl4UxscEbSHsIaURQRZ88Yh59bfdcM
mmwE9wQ4wXBjbMk5YXoiSTq7G0BzvGllinQ1ZNrkk1//QgvSerHt40pvCE+LzmXX
qY486TU5+7+yjN/eBnPDd/LwV04jWr2HW0hYMoM5rhQvH1ywk/6k7Lh0fAnkK4VE
uyS5TTZTCnHPpq5TTKdAD5na05JvpQEciw7oXyQThI4a5w4O6XMmRwjh3Bmi4/9r
PEo/5OnA4ixI6WqhwBByimy+1oXvR/RqBRvg5REU/uF8rYonC6iZVnN0Pbzu6lXL
KoztWfHug9167WeSlVsipKYCnVcrzb2zz4LWC5qQFNl8fPf71vHjsIwlUGTy5yqW
l8GgXQbQDvrxpqd7siGmm3aIPKhKIgEhhFn/YfRRnEm5a1V/kJDOqUwT/03SX8qH
R1dm2JkaEe8vuLWtZEy20Plf/KuuEIP1Jhd8o3K2fAUcIuaio0+BiaRFJbhVKWp3
6VrAPDxRXaeeJv+IRlZr89OpIwZJOT9ZXZAdw8NwoGbI1KUBlsptqQyIq7xrP+ih
ktETlTk0eC9/LkDY10z5Kfs9xfnfFR6ce5/wY+iA9oi/WM39gYMw4KLfg0GNIZeT
jlow6DE7xzMDmP3ScklfLBRIU8StPqWufDcUG0XG2VuY5vXeIQnn3z1qN/zrNrPn
8o4tAFIZ/3CTZxAA+E3eRUyrDQT2qBvuXK3BpsFpOIAJZBOiA5zhVoRdvCOjxgDE
3BK4wBUIUnMrvD3EgNzFwK12yWRCmUWjr5n9Ut2Lc14jHiidnC2XC5fLPHAaO3nO
W5oIlvVbQuDDTxfwgA/MhITh8zZ0DobB2B5f3W7Shs3iw1d5va0DWjXQ0PuYuKPY
zfcRvq285mgrxDRqpg31YbXiJOc61+LzWWwGlW5wKpt6OtvHGuq7HXUjfW3pQT6k
DSkfp0q1gHWZOvhzyRGK3NU38xFe6rORRkgfZR5KHiXiwH7F0NIDD1gWKa83E6ik
857typvXDyxY9jN5HCwigOo8O2u5WdxArz8kDmMR1NDhPQAXQoPv3VjAQ9dMsrgM
Z6+1uPzqaDKSe1f5Wvpz75BISL251nSAwBq+jUJu4L1piJe4iJISE95jpA0GkOgY
EeMp7KZL9rehxlLU7LHcfGPiu+g7jUHtWtBeBwOzYVGmLdWWzFr6H7Vnr/I4GEuK
IQRTTRILADSVxOthIHulUNekmNnMZO9DJ4Kqb/MBQC+Kf6GajdbmfmdpnKLI70xp
fiXtGsuBKJlspB/bTRHelrkWOReiV5sOVoQKT1y+SONcD1Y/Kx1FvSS5T5uSpCs/
JIs11uj9mZDFDJHhSPcw+w/ZRRQYQs/5akXc6NVgRQpHTKqU44Sb2gDfd/7r497E
5NrrsvtbBTUaCIRMzRhyX+iAfLXlkP683QY29UVqnNaYuEvnwmvUnzFgxojV7M5r
by98S3AHj6TXpDCjmspdBXGm9S2ye/b5r1/o6nlX2YgC/jAIPAGPHrrHb9lIqnbD
GjdzKuZtGcxlooaH6pKGkLHsQ0ZhXrn+2zVWtdG15mruBF18Ibe5D0WqjdnOn+Jb
+8Sw12makqE693z89zRDnXLzo3NBaWd274zmYkg1C0fJnUGu8oL+Ojd6yaVOB8Nt
VaQbewqoYg8+ZRzM4BD60G6hF4hsCegi3unjiAaGR3JSE7WqfWQ11VPLJG5Wly1v
3BbegTfsVSW/Ly0POMP4kgMLHW67KT+z8ZMKIP9uUsjsy+oGMj+ceoOLmubvXL3X
Ud/CnB1Z+pWmgkNVUwOeBeY4B0B+gfw8gqSJdbNTNoNAD925S/fvajnej+VRM9pi
o1Ex9+LQzGPzU/wkRW5nqGBeei4RRAGcqD/FUIML1ml487zjvggJexRmEspA6mUg
xTuEXKOh6UTDWcKFsb5KBL1WECWbghf6J4muAMZJHWWFPo9jiHRYMh9bxINHLS1T
F6tdrhRaIXUTEEwO4hXPgY+z75t2UVHH97TMlj5kQpOz3gmpPl2U1eSKGFMIHY1O
ijerfZOsLhAqkGAVIYvMXbiLYOJGz6hRjJn4ll/nmPwI+6QCeQ7RMUVX25VZ9qDk
vjvuUPBxLaeU6hNLvgnK5sYIArHWxXw3cijUxObXogQqqlb4gCJ3ai29+ewbRpxS
KYM5USvrEXfXrZKpWYXSqgcXMyEB/SwoUgCSsgS65DFAOc4dZrifhiaTlqHQgqEQ
LoyCeAdAV9wWdo3acteGpNdtyaGgkejS4wj4NmTyvIT55aVlZLDhBIs1b6a/rULv
O1rjEAMv6mOWEzpO3C9cfMXVwFVU2EVEKzf+9NUW6aFLqvCYJyQrhpWJmG4cgwKc
3NdI5Jpew1pcdAUPmbU4II9u3y7qT3VZtna+atRE74MD2aa4aIzo/CHtF/89H/f/
FrEC19YbCBz2whrX4GBWE3wu07irGAtD2qJnE63FW0HBJ+ariWqBqx5jTdseDAvk
M0xrZJNiLvm98opk7AhNXoHUACwueSyFwqocCW92HVmN1Bn0FjneNXcKADNfwy3t
Vus+qSYihlkEEePoZTv4c7fF+RAjVjLDKaDbxOgK+3MNbPiS/cRIreyaU7N27EBB
61L+W+P+7Gg+P4kkTQscnZjfKZ/KyXLv7AaOd3xDjX89tMx+vPfa3sl4ExYZxWay
ZxR1v2ewX559ce7HlWjgsGoK10nU/0LpYo9nqxnaXo//Spqgd23wcHRNdzizhCYO
upXkmhmFsmM/1e6BiufhzITWzeEmzyze664YQDgaM/bcrdGQfcA8KLNW03ocQ0MH
MQzKANCBIMFzYkR6qactei6E9NsOgolSZDuL/NOHLw9D0hnZwT8ZrWmHeW3k4Lr2
/qDI3cyfstrFk62Qznoqprk5cL1ysWnVnYtWyIXjbTOJ1unKGMWuqG/BSf6MNMml
C+7x+/wM40JY9BVFgzN9tA/XQxkqk60cfLcKafhOKIEcA74vo0LD82DkzzKHydBe
z2zuGRa077ApDP0HsqJTWZc8V7wSAVvjQ2a4hUROZDpzaJtbPeeL1YZim/bPbgZc
vJwvcW2vdXsPIroAjXeC3drHU53X+xVho9Wt/s2OhthNfni/b77/qQ6RJEl09pdO
w78cjWZ3uwwIKdswkNp+tpNt3JyZVzrXND8Pz0FaDZPXMYtOISp1JLiJkmqChbev
FDh3wnn1uXrg2is9f6BHOAIzzI12sDDkfXNVDdSLa68w2gBop5QoKnu+StPbMCud
Tbtt/llBMJOdIGfp1ArU8LG8FDfb+MsHDqLPjR+w9dn9ryWhczoxaf3b9jnXwJ6Z
cTYY5C0BsjgiWdl2XYRn+o0FDp20SeWXylMKlHWZpOhXRw1bFAmdX71Hvb8NAWFp
MMxEwtDbBoRYee+iQiHx7Jbm7KjN9LvZ8uYK3noVH4p/o69usZiST89KukqbivHW
577uNZ+zdK4tS8TwWrytm36ZPnDyyeuEcepJVoiIx1QRtWp09SpPJ1bRPqsrRfcd
kuRnDsUb06lw+Hn24I2eWx8ExcbgejHHdMBGussmBqLsAxXRAC8cLaycsMWTj7Zb
YYAm+OkcLF26iD7jG2orZuUyMbg8tK1BzyGg1Gp7+koJvqR1wmSS6htgcVGo0b+A
/msf5xeLTkKryW+mtt5ptBldqcGyKfYfENt8+1RfGo5n/GkCuXh7KHNcwZ/miWcM
2noGQGTz5z9pfFyPc28Di0TeoTljbPDZ29DT5eFi4vQWKKw7KTmG8A4YhCwd+yy0
fEyIbE+FRkQhs4fYVoZbQnl3X9bs0SNsgbhO09F/sBuwv8UQKviXpJBW+S4jShJf
QfJCuKVEh8sNkYEZ2Xzygmq1xH0XJGwykdrSGuL39jdCLznimjVpnndwzvE+Sdkk
PI1BRyuLnOMm2UQR63duqzDOjgVC/pS+QGFvMKykDjkW6V8JqjzomRMalT8smyt+
SW9uSti1BvbxHY9n7VGQd1aOQIe9Z4re04ybDZzpFkRHFRVOJKexc/Mg4204LlQH
XH5tJj7PCbIhcyYA8Uuz/Dt7w2VIOftaluguW6GDUv9jiQ6p6zNwPbCfKg1Wxj8/
9Q/CPJQWIl2Fzj3n2h1NpYBsgOMR1YcgsesZqRzwyxuoq5AT+biONS1IymDfrbRv
dhqWZLwYd1JWpd1Xg+VELFsTJPSdkzuo2sxJG2f8tvyd8+hxLStkdK+Ygy8i3u+M
uYnu3cuqEGPh6MprmyPQnY9Sw9dJ5wWUT0/ia4W3kg3u4hpWBS6zIMHomR2MsUkp
nrLrDchtBXYOq1uMWIxx4zORekywPFgGNQm7RpihP1pYpOw4OQB5Ibhthr2JFwxt
OMCD5Em5j2u7XoxHWtG7IWJnQ89KjCtnSF71R5QhP/hvzrXitFoCg92O7fPuFzwJ
T497T8LevGspUMbHZhMWLzYkxkb6JN7/Qf0j5Owpq+yLSNWGnyYGS2nY4i7G69RQ
tMb57EFnspPwshATESjEOP+5Y8kmj/HhI6KljBskt7qnL2GQ9X4Z5UwQaSgSG+cH
Y3QIhJBB+k6n56LeScYr5xgrOKmB2/qOMl1+JZHb8M5p0Xpwt9v1F+RukQAoiRnT
/0LH5Q3oEABMe1QQCNO7GjSa1kug4In54u09Hiapg8hgNHOJugPtG6E++QHValvb
iZBkM2+feakg9WWm81HMc4KqEPA5XVBbxEzZg6hr3PGDXSzFgR5boz1L4SWnRMdc
6ohVivXpW/sBGbqerFpaUW0OVh16C0F6c/aCkRjuT6ig1o7O6ge8DvAX1rpev5KR
7KzkM8uXXr1hB6Tgu4hDneglrH9hx8cjqdocEAtRppvwDg7knWkHKdbaqapZxKhu
Xy3yqVfXjoMBiBTEuzyxMEH/IlgudjYutIhHKcNtfN4CcLMAB4WyHv4Z+KlZJjKJ
0JgrCcJyPMpw5C6N7GkJ7T60v6qNS2/CQcUWlNkvya0vADefsrRqYKnxfL03Cafq
8+ms9buHv5X8f0M7RWEXAuhOgZQ7y6LKhqqw3mfyASgFeOobNwAZjSYTJsqTeBMn
lJ8mpf6Th9MDtvGJABZOvGENcZaRevKdZ48MBcrBTfUQcaFSS+zuyn+hhbc1MPUa
Ki39En2evYd3BWV8DvpzIh1o0Xg/lpj7NNr2kGymdAhheuqDGG7rMYFh7k3J1VrL
tt4QPEHcPc8zbWapcjo06CN1jZzIf6lpEYQa8cI6fxX6tR0oxWRwfDkjcVlp9VQe
YeusRbPvAu3K502F/9uR8158qLJEaRN0bCTo26Xa7gc1Yf5b4660hjnbblY/z3B2
Hke+7KTQSo9haZJxDBXaYGNCIOt802FiXnoQK5IKQmX5N2OyratDalWR0vPY8PIL
QzjNXxtlRfCImWAIko8jv/Wnx/p6k8AsBNSRjdURfRoKGanFhwD8lY0J3IZk5rQ2
qft9F5D+4gACU5qdMmYc/anHTAQ0e9VEQYfN0CMytFm7IbC413zpW6ZiDhhBx3+l
zsBcIveD8hBp35ToTnLNgjXDyFsFkV0j11MN2E0VGMNmbCoP4DxUj+tfhgBtF9dQ
C4hb0XXnMCYAXcbgO1tvAdr3IVVK8Cwc+oeUqcAofeOzTDERFxO+KvmF69Hnc/V9
mkrMUPfcJ4K/reGcdWrh9J20Q7BqQLCnaiGVlKVPi1pIvYrIwO71cjWRLNhb3/TY
XJ91g3+dgCdBpyzAg8RQ6IDjkMdO33jRVDUKSZJoigg+wyLcZjOB9lSDaZNiNdgH
+sC7O4h7IyFCvkFXXGlV9WKJ4PZrq2wRZPPhgZAa6nEzlYBhXVqwM3MV9n8sDpsc
qZUdADYrntGdwjMUx3XHS44Vp/IqzJFlXmTcBBsYzQQjpSUJqK9xjNNzCGguz6CG
SVsCKWQ3mIL9Tmggm49CyYZa1h/4JDSpsHXHVdKvUWD78+qD+bhnJIDYGkJct7Gz
k7SLSkJShe8wGwSTraPF7j5WdVlVKEWa194cNMn7SKzln3cUC+pvM7g5C337IjuB
3XVtHT8Q6h8KenGTi7tSEq11IGiOOVQOVCJnnhyWQJoTFj8kzelXedQ1d5HMzPRV
ORJybOmSzHYZ6fLI/FFzIkvLEMI/K/WrOd+T1yc0L3CoipF1z5RFVETRC1xuaN9j
Cl4clWd7P9HC0p3M3RjGjPeq0dWFZDuDs0AIN1lHgAUI9WEk/h3qdu85crx+oXjH
fEOc/Sm+nv5ZzKDHccNRuOmkf8wMuttBjtJr4ac72O/6kITGTJM6zpK17ExF9kI+
QVa+Y5jkr6/nj41evtAIk8085XqcErQSlDfJ8ikfY2h1BME7rCTKU7RY8Ljf0xT5
/wkIUkjl60xjrh+0hM6wv5z4Yi/rM5wwMRLmuXTfthRK35pz/OthpkvX5ERKR5xm
XYCQYh/8/laSOJCoVlFOdQg5mOYJhm0ZOP0jP9NYjJeTlwBTrTrwuAHhJnHTl/3D
BFQVcFsWieEAVWZas1E2YT0blaM1R5EJ+6P7AjBiJDL3dusTH3ZFKU0prtaAQnpk
HP34B8Lhescs7paTSFrxoZJ7KsgLetiFfP2HHr8WS3BTz3yaHqi4f4dqui599Cwd
jqj4Zoj3UE8bHewMjuacXukKrHBfn/KpuRNFdu4UMoy5zx5bHY84b+2J4kfw+HRV
WWZrO+B96+WJY5/rymq4Q9AKJ/2KuFa1V3WssCASscuytOrC1EhTjGZG7MmSv0wv
t9sVb6J2gWLUrtoq0rba9YUTBtdw7F3OCRuhV/UK8wQeseJkGNwrH6026AWpVCl0
1Te392InsImMXec7MC6ayLYm7+9MmaeztvZmL0mXe5ren8SWW5tWeSZTPTkD7Jtl
B8Gm/B4MKEt+R9dFuMnXSl4V+/+r5m+cex6O0qVsXNsSI3UEQT5yuvR83ty4Dfq+
e2A/MAFgDMe9Bc91wNQ6phrKeXrbUD4OYie657UG3NOj8guPWhI3baXp/ZwQCAEM
HXeQTEO82NwG11oxYZ+qI1MVv7+/7rTIz/CcQAh5RvlBKbSLJb8HqDo+b6ISzY7m
lmANA5PiuyyqvXPQAv9+XpX8xnXd3eDJQFt1SU80lLndCTLnXLGkBaoSUsvqqDHq
Uu9mP060yVpnvnCJv9BHjBiK1DHgC6Y6ZzuKqISuIPc5MaDRu0jCUuI68aCIqF0a
nXXlVYdETDf/y8ewGuaJFlDuFhaNaTJe2T92yRO+DYXFMpNupUbUjeI56B6k3F6g
RHgDlrh8bjbymjzZGmLBbvnkss0xoFwvqBBkBYEmIjQ+qvFfiLnTXCpoo4s59FL6
NPt2Gy0SIYTHcebXjBqM/Edou1ccEOXvx/Ix3AHwHBs0T8qcrLCDpzXcop1xqxq5
WF+WR43ZF2LwwKd0gEklEy+BsfQzsVHex+81Bvn0XyoUV0/YocIpCJAz1GZAEBer
enEOnZM6KdO3io+6QGbgErubhHNruGejXdjsVER2on0Efzb0puY1tepqmP2YauZF
uidWiEWZcyE5CInlOr3zAPvIAP5bG7OvuUF/d92cVhp6XNRwXGx8GQdCmmP/H79Y
wfKUsEIERN3Hl/Y8bGx3lpu4B8n1CDT/+HjtOyUKpHTSwuhhP9bkH3rDocEiBnPa
LlMbR20/WJQdRrlRzEmkuTPfZYe0MURzN1CORY4FviAVJa7rlaQC9o/nCHJYy5vh
2lSy2JusVi9YCy28/lFlecwrs2bQlL9zSCcv1MeFyXreAkGvbn+g9ei/cDBmP8N/
Zrzf+89EkO76jtxohR3ZG0GzP4qqVwItjxqGW1wJUmUogXUk1ubwPrRCCyRD0wYs
KrmN1wA498WjQEVo1Q9tc8x6m5NM3ENswtcesC0KWcZq0mXR/grTQv0wPya6JhIr
K5qdyoQtsfDR3gzK2UGnufGUrqEcVmVHTNNH1EzbyguRjmy+sp75AVWu+gV1Nzgw
fJ9TtvKwzFODJJ+1meHm2QcEtVsfGVc/mWQ/7O8VNVSbg24G71M7RyeyNJEzqsmp
HxLDJ/LYiTVUthj+Tzpj7BGfL37AqJoI755PTAsu6xQhBDDchQcZKaGHNF2hIWP9
PixAhgDkSLoS7OJ/Yqg9yjBkICW4d/nwpqNbzSEjlWjFijS5XVVIwQPyESpGAfkS
bv9qY0ehWfAdIrVVhDVxrTrhPF/vbpXYiqi+zUWcQQVbfD9l9j5F7WmORE4+ZNcb
1EBIYiPSp64fzB6QRATxM3P8IBZsfuoB32iys0NDq6+N/C+TRQajnGe3pmOJAS6z
+GI69utpwnY2beQJBjyuu0oaw112Ynervtx0/6H+OoxTDc5t3QvGvxewZgHkXvjc
jEcZRRrXW4maTAPBdzeuBoHS5oiMH+3EXUXVs198/08wN+OhbUs1UbkSOxcYRsU/
qMQ5BLCHXg1lJAqgsZrekCw6ItaxmRMcgZ3WIRCP0qYsolElalpTaGzlo5l6ypHo
l94Xd86/KyQf6YwLup2bC84NOA6vdh9DSoOz3oFSY/vULqk6fYbGl1mPTIU7Vf/J
E/EegFJQo4Ap5ppRFCmAtBaIKtINgNaGi1uafluvJHB3lDtl1+yNkUwCP6AIQEGd
ZNAcZJxSUHMfIdt6kULL573ivf5LlSTHsuKsqvOoeyV39eAHmMILcA7XCK5YnyJj
kZlXDtYrQIl2tSQZt3LwaWnWxotJCLSq6n1lKyFOV+XQPlSnPxzjzgmGjUhUl5bj
qINaLcgftsE/6mUnwpCFoNzZ9E9ihd7CiOYPLNsBaCjFXmDhshsegPzvgYfj/URR
Uh8sjXCcq76DHKljcF4lMRj3TFZg6IQhma9YVJX/B9sW7cfBav+7bb5fY53Cq7MW
Nd1TkglBlmfNGHJY5+za217g2q7kNYVKlpHUweXM7jt/IEvCzrp3tV4FMWMFSf1+
kEAD2NnJCrL365Bnv3CZAbyEazDsUnFpg33w9bGtacMt8I0P6wGGvqnStRWySSuy
0u5eBVY/TnXSbe4C69AsPemJ+15SAsDYyGcIGzkUMxYbddVpzGy2Oly46TFO7m3w
X52gsvvZCVR4TdX2Ka9HeKAgAQdce+EtjHxrPOP+uEVj7MHRMyuciBjHyPwRd5CS
6UDeqQSvTpl5+AAbOomXVlXkW6PGrpqlirBfZElvCBgtSr89CVRWLBtonqGaT8vN
ePv8q/ZyjViyFJbtFEqXVgspm8OHoVCDkyRYWUKs7u5uzdkvw0Kt18OtYKSnwBeR
fTi0YwSBb6/TOPX1jzNaDus+2/G2mJ2sDd2WA0uIUCad3eK/THdvsMtVD5N9xxjC
SJeGtrKSZyuthSN1YGlG3ZL6hyY3RHSc7t7p9/OpRWJ0toq5VWEILfMhSiA1YfLr
9zpSoucTraEy7Z8l5sMSX07THpVF0sNDrkD5CqR0uaxLmfRtEBRZjio6mJcTDrBT
vRo7vyuyU/Z8fnbXScLvT72S4Ym7T5Dh1XhgUhENk+R2Ib0gkueNeWtBVNI2ukl+
ZWBEdYtVMHXDVR1zz9TQDQXO2tIShLkOBV4Nn8S3zrXYROfAa1zl2eVD6kGSZfcz
/UM7sjGEB8jGopatp91TLOgxL4eTNaAacNc0EjKekMVmWNx0Z3inGSWIydNoeDnV
jY7LZYpszU2DR70KEe6cVri2rTL+ETPNHLDwEV2pJfGo86RoshDf/RmVDaezVtx4
lFJcrR2lAU+Y5bmEa/XJxGIzlA5b99FYM0tS0heWbM3YZ4DEx5+RbCTDlIxMoTu9
xWFfhrZM0ZPWAlKsZVS+CJQZLXAJB3I1DU4pUlv8twAZohp92UseeoW2NG8wCAgt
jZWIS/e8ijlEtepHvZpCTXZVyv8OsQ6RFx3ZOiKFoVOyrq/kut+m6f+jzM1A10xn
S1DORR/Fbki97qHa+Mf9nlgKR0tUk/AjE4Vu8e4ZLT535ANedPkZdOMRRtyrBu4u
EiSSA1qOfzYRhUWDnPLkjPnRPpIhOdnC2ZOVHeDkX/esGh9ivlhPkJbKFumvvXHl
ZOrtLB52C2fkcJG8oaQZ0js2ED5/Pp1ZEiOc2uCB4y4wC/9b3kYPK8SGE+9uYx6x
GzIMdjRpp5f+GR4jlWlyGTJeihFsx2rF3SrDm3Tvhz7O5qq/bP61ce2C/DsIMcS9
GIJow2mS3dr8EkUgw88v+WDrOYdyEJPI90D15KH5DBTmw89vSEMlzr4tsNtuhnY9
x4J8svRLUV9z28YxJFRIcOD9B9NJ/5AGYqEqDdLsg2QljXam6FJB36CuWzZ70NfU
7I/8LWXrjXvRyQYufCZVbqk5enUqCw4eWbKApSG/P0kQ3AHEV1Xp6qDGd9FRf56Y
C+cmWqTV1al3AV/ltfzd5k/V2nfazZlZa2xpjmjzEnAI+DVjRdFv3DokY6MiHkr8
Zg9ef166Kp5Zcj9Xvg4v8prviiAARjCy6yKqfpkQ9rpfy+KM9bSUy8+JKXnJgcyW
ETmXLRSggK++H0/460AoDF+3/frFwXrTTkTByCSmMbErNSskM45AcWx1odXIli2p
g8AhWdH4kCNvL6jGHPBUpzmqyc2p/5/mTWgqvkC/54d7jIhCeF6xZ2RY/wBcsz8+
QiOcg2zOWoNiwjwPKPUn0l3u6l7YCFvJlhTsNEMposHrK9XHqtJDhMBQXeK8L7eQ
2HghFGuZa5BbEqLacUjJAYh4/WEInRCV1O5g1ibihJtDMplt1NCZ8/XqbBcstkhM
EbBNqSS48rPs+pYzQFoYXMdG1MsbSCyxztmlVIdJQVTHUjC9xcNLICq8ZqipEvXl
B6patyOYNVl+9CVS7q28pmGhelUYCf42C6XBFr18iAKkl2YvD+cKq2NlImjmW6oV
i9QBsmHPILtWrvh97gcW6Ang3c/1++dwmdpxBSscPglXJGJ0J11C892Geunx6WZ7
W3dDti9gcs1Zk+grhPdicZaTGGJLyQNjlH9x75l3TPVH3bflK6AOgDctO9WK79nw
2drbdwfUOU91PYYMny93sHuvXLH9Hxvu/WM4wDqcLRSNZPWXXO4hXYZSsFk3rIyQ
xmqwMfJHAFJfEF9AlgLcrTgGaUN81aF6yUxFp1Li1eu+hSa+nsfUs7+1/vqneI3C
264Nkm2BsrebwxFpr4gA9yXJp6jKkyG6GDyUq5Gl/2U+7E089Hvun9SAOvlFC8qy
vSTgL8rz8greK6ZHEhyZqIINK9IzG97P/6VNHvvGnY3ipvXjNEmnddzPi/RUu1xa
a/0Tdd1GAP4CzE5yMtVMqIGH/Zyyq/JwMRC9Y/pYY5jJEIcEEcg5P04d/qmFxI3Y
5n2JMoNpYzR6ZE71M8exaElqldW0brwv0ykiw6/PfiarSg54yfaV9tWiaPA8D+bn
zNPsVKEvRW9xkv5u/u5imLoWtS8bi00+hURfzKfs84PnY1J90FEWtXArMjgDrHf/
u4FxtNDj8p0dmcO/WrTk2MA1so4hY3zQRs3GGPnGHt31ehIEJOzEWEGArywQEPJR
6vEKNkumlJu1L5DtMzl+KREYfTf33vwfPDq1Rb8xbZI5OGkist/WM6JPCxynd2S9
4/AGlPWBqsCOiZD+nM/y4J7V/CmyP4FGNkgtH2XubuN8EZuWeJWud5QmOS7PNzsE
w6bnV4A2FcfpdazmnovHtHfegcnhXuP2EBra/s8Z5S1NtkCt873ui8d5VUSgfdDe
JaXTWqWAvbunQS5VsuLEdIcMFh5G1N3wEwjJWips+RqGKwTeTQXGEeR7YiuLUdKd
ZcEgCFocVmxVp1J01vhLi7DWkMCDrMAgWZ/BY8EMBXcDsheCGztp6MsHr35i1qjg
t/Zd2CSRlTug6S2PcdmMtPdVZsq0KKytXORhe6n6M737TYrdnslel1nms5DcqHOI
BDIodjDKmkNSeaJVticvnc1IS0YAV09rMhhxDkRsP/aRFyBiWULiuYtCRL+OwkXn
v6Ka0HVsyRp6fZi4LzgomKF7AU+8h9TBK1WplkVl5N+wXwK53SV/6PEpQAVcfrBU
gW3iCY7tDdR/+iWZOJaoOsReGnAkDDqU250xDpj+lYmTLi/r9yY3ar/trbXKnu8c
8Ik1W2KFGspkQrUKch/hnBIzORxFWBVQhAUkp+whUEXa2F6wlgGILJKZu1prQ7ap
JiytVfCtkYvkh7tKQFZWmn+pvlkQUQeKxWkFmsIAnlDscStykEdS68RPRL0XVgLc
EWK6SFz/EMv3b+7s7B3aHKqBKXCbpQy0tUuLESU/FwRCC+WrJy5DtpiE2I8w52Bs
H5MWaodJZFBjKQUOCDocqFdHNtZ42hUHEf6trbteeoVp4tCnGmuBXfqXQGe8LoeW
TqkMtPJjJ0fAV2MAxEeVMsQEdzSJilK9hOzLVdzkVJOMIg2Ol45BfZa8JfIrELFl
3wj7o+FWOHUjVfQ767kqvKYWa/sXobraPPvfdG2sdI935eUAP3nTv0OAiLHeGwOa
S3X1D0z7j5WZvJ16IBC8mh9Z4pV4R/AC+r5ARUzaLzAMXwokCtttBp9mnnHz+s4Q
ogEJb8aKejUfC0PL9U+/XjOv6dxQEAUbHmVuapi91FpLtCdaw9JAnVn4YNEC9ocT
MluOwDK1JoAZxeCxFOXUQS/JusDNDmx58H8bLJCqjNFqZDKHpjyR9cFGHAv1nSbm
t85gjfJ+XNLeBb4TWo5YcgLGYwo/sVTe+hbc8re6Hlws/CE0oXoz28wktAqrc4BD
5IHRQex0Sv83Z/x8ge42Cz9yKFUc9jRvveonAKyHcpypXzJ3Jh8QcZweSiTDO471
hRJV9N2cthIat240qBoHqbzgK8qsIkOSblHS6imqLGf/uUpxLdm6cDI6RgGP2+K9
luy/Q54UmrAtxFyrPG0XPWksVjugPo8iaHxvXoFBM2EJ5RKFnYG5AP9jC17bYysj
d3az7BbJTqKt+7ItDdOe7aFf2Stu5apkjJEm54TlTiBkrCtDC+PRxCylfCi/7Whn
SxHfecUVJRi2xDjBV2Fjh7/HIyo8pPeZKYfET5qUSyXyhtB0g4XOG66+Ls4Q4S9X
X/vKNNaKLMCAbIN8wGcvCGt2iSfZo1iIEG2CY9ZkkQE9lImeeoh2e3fuZAepr+31
9/qzOpmVrmM+Q7ET8T0PFhCTRVdM1smS5f8YuLozP1ylnBHwJVxZUoGjedai79B4
atyhwRbd0BS+ay6z6WwzOSdTduxF7mZtxZ+bEm2/nu7K0vY9pwc0ZIYzd0sJrOf/
il+B4KHjPgm2WsdV6JsJRErzcE64xdjiM2qyjE8VtWCADjCTD7rurR3RFRhc+ym0
jiYiJewur55+wYhBAsamv1aDGnB6a7108Sg3Q/HpFBIO3Hrb/eEsGR1LytgA6l4z
hZgmLTQnEDWNuzUUkbuvlLRsGBGLGJlniHsoTG/WMHrQqIQsfK4KEJWd36GI6DYF
+yGYqLWTUho70mKrq5i/rF72Jk8oa1t1+xQYVDnYwqfouPQwcOUOJ1l17tNYTMZv
y/bTBrRPNd30L47Qq+QKOQ5rPZkuGsNOLbtCEJimEaXZpn+0wRBmSds9f24nK8h4
0bckgYWxLV2bzrI2Fgml8gpj+OvMZk1IAT4pIVSqjYPXBZ2qZB5HoADbdRFFa1BX
KpxgwJUIfMwqUHdJep9Wd5xCsKQqC8leolIJqoGbCdcu3azYFVGWqFYpfX0OXg5M
lUkFGxkz3ExzP81CaMPd8OllEHOQXs0d2deMcSxqsxlQ2Wszh5kJE4vAmon7BWrZ
C51mcCT9Q1gSEipA6awjzCsmfVxJnbmSxP6+EDjJg8OzJX6OtIRRqH60zuEbV7pb
2B7OHNlPUxDIqycI89OJ0LkG6WcwqYnVFRYgEe/7LN+rDtgOvQSsJLFv9JNc05Lg
oKLwhfMkqINgCEzLZ9mjDWjyAOVJriz+QaFPFNpOzxMF4G+3Di41FmDZmxDf0NXq
6WAtpi9MasxlQr3AS6jf1QOOVWqpyJonpHBIWzEaz8VWQkbywb30Q6RCh9Usf8BA
1z2Jfjmk+3g9fueFZN/tVJ593imexZYBovFPhAK9LiBtLX6K8N3cHTjP3gzR1QlO
oDLkw/JeyWPyTi4mXJn32ekUpGLxtLOSIXdDkqrORP2l653egVp0wbdUCktIG297
Pz89oYjTIiiYfocJj1jEs8I5WOfbWpICULaRmbq4/eLFeEmn83ZDxwD7HbXdZUa+
Pi9Cls6CduDIUeFVPOCjtUyzcxVxg51EOeRtEbSEJ4CjOL/bz2l1N8Yge95bn+Hx
+cDJs5WeXF9xUPbGj74NmXR6INFZOMB62uM4mD92xKSUI4x1xuTYQP1rHqZLLEkG
r2ic6RJF6w4B5XN+wv8bCQUvSurME0yJ4NKzZHwBtBLP+Gm6wCK0cxDo26hrcXj3
WJJTGwuZsSrVlIYyMAUaeNZugpGrGIgHnyPoCBoWDc2tIqtjWe118NzRQQOmpvv1
LdtOUm67DFcggZeks0U1n5qwFEqYeLcjbZzAN3dOsoohFcc+jt0Bu6hw95bl9XMn
nA0KG47VD3f/ytCbV9gAEC8Vmrblxh5dp1K11+1sT4zjmt/Vlp3gFPE2NsZZfujD
kqvifCl5tjbiQthEDX4lqVodvOkUcqeYrSp42Eyz7Pcr7vhyO8uEVB+qZRBhFE+Z
FRee4KhlA9nLkEaQc1odB9BEqBsoOtPpiZGX3Gm0SsMq0OcOktxY0Fj1ljB/tsbu
ucJbhLbLLeDEopIq3HLHGhF0O63ey0zBXkBFnRgOkTX8P/Kty4EiyfjCeaWl+C80
nCbwHzi8qq2FDjdljsPGHP9ctgHc49QUzQm5waR5+kp0ujYuNk8UsTysqsznLHwg
/bMMPI0oMRSNk9uaOqJ36gLcGggKv/Jjik2rb/rn6K2xmxXwNQF3dREfHY0PqROl
bo1FmVXKMoDhFqUhpww5Ez3hIcpt7Og7URQ3Wol6B2sBahhgUG2j2qFMPzdh1h6s
ZEYyt4Qw3vr9RkTNjE2reXpQlu/6CLO1wQb+sviduLkZ4JTIxBhHUeDEP6pFlkNH
UXWJI+oyzVwJBlmES4TtYhDFo8c17uHSkUF+WDoPmn9C9ApVHL6xD6uZUf9BsP63
WCu3Y8TBuTCUKOYbqO+Ka1MMerTPHGdlWnPC27YIIyVOfRYESGNmIJqwWiljR72a
2qgqChvNKYju1WzYMagoftgu8hGotgMMrnBghdsIDQM1DEMJgNC76zLVpAmIR1Dg
hEkyNqu02INN4l1Z1d3nZQenX9g1Wy1rb3QUIUAzd34BZ88b51y8tEK3RQlU368I
ZPfg4m+fihIjn21gedVABBxaPm+Vl2VEiflZsgUSV7mqWY+Q1kvmr0PbYd35ABrL
JqtMqP38I2GCcj7Q0LJBUkWDldt64gtbvJV3lUOYkyel4DXmnmvRX3CP+x7Am5zz
zHT1XzyFi2+IexFNYyOGtkoPy0elvNbTTn8+Mn/OgpgenUkwwuuwH33yIDZViPFj
krLDGt5iKrPVkhxJCkqGo06GiLVhKx/OY/qfDJ3JVPWmmGxtD/wPvIclcjm9opeH
EXuupMznzweWxt26MibvaVOLVz2CiAxP3zOP6+g4JHOZpEg2LeTG5EUTE07A1D4a
xQ3ccHUGwYAd6aXAb5YLHrdEWcVh5XINmDnnNHjY8pzKi+uJzNUKDDUR2BSQ77kW
tx9bmVwj9cKNWDxYhI7G7aroxWdVDZDDVQ7+TrHCO9ElgdYt73AsLRvZI7hYPzjD
EinL0qqd0nfOvIieEWRXWHQaNHjZNuSo2hBko3UX8hbEYvSRysn/byXrNJs4VE6R
RUWQmKQlazZBv8Bq2bdhq5Bt+BTUBAX8OfPffoxiY47+qWg5LYc3sutaOWgs8LTa
a7oj4fDBhsDeddaG/+c8cIKRaycRA5X8idWAhZsrtCkWKyKnPJI83Mws2YbdpVqh
T2GVPiWyztgsJOp4YQF+YSJ7STJeIRBHq7Dv+GZsYccPobZ0sN+yPFKUNjmxSmMM
zV6Qpqp4CwnaGPj7xoQ6E30zZFLVU0EbnvMuyJqpZ+ZD2ny4R3vDe2p+yqjdZBg3
ypWw+JDObYVhm9hWBrGLMujSh7Mdkcsy4/Qbez9UW1yPbo1zuEfRMwZ1PukIvVhO
bOWbx371ZDPQoVBupKotsArhuf5MmtcMzpPgpbU/dQ9wzuF/5IIFeCEdVHBLsPg0
veKDAaMS6Xqnzv4/X0r6TeOVdo3oOiYVMwYLbDaX1FJd1SzbgzxnZC17D+/bXgtK
+4d3H0KdfrW/gFlORt1ilIJnEeHdZia9cStdbcM3L5TZ7+Z7PaOvS3NHRB5O4hT0
G3mfFF2+naYlB/zfMDZMvrV2X/dai8PxdF3nzI+XHQyQiRWqdT+CxvysTN3xsTRD
7CsPtqdPkMZguAtTzq9KVT1SAhGQFVrYNz7HCxD8q6O4jkcjapJm3OSnwy7U3pwt
CMAMdOyc8HgdC+h3lceOGhlHYkfG4MbQ7k2GNKLKXscGcgoVEbKmaMM/34hZU5ec
AxJExuXXGfZwCFMBcXEP0sk5k6nUVGk++/gwZ6/js40HRv2LZ2VOJ54pRdAoIApf
h2CthH/30i0OR9NEQVVAoEY5U74QAA0IeVvj69eZbvKMNQOKSIyFYZ3v4crmEsL5
RG4wrGwRtg2Js42brbgoLsz+akLZbl4ezDJiwqSQx8xq78+HHCRQKJNm0sYCuOsc
I5y/ILeQFyb+uqkrzPgQS5R1x2LqCZiffDB7HdtKYI2iS3dkrslkCSdGizGvdC/r
AhIW9XvrC0v6dQDZFghceFrTbAzPHF3AxnOZ0lWO0XCAmC5A1Iyvn2zvSR8qpXtw
TEiykXJjv18qcNRDBCXNcbMCAK9AOTiMin+y/aVw0uBIuT7P4HaSBziPPbKBHF8b
EKU7ovp+i0tVmafoHIQuTBXaamC44FTE4XeFlAvg7C5C/mLYgrJM19kLqcFRf8wv
ecM1BTyACnGYEmo9h5bW3FNlseI6kD5Ja9+Gf6rmL+wC1Mj3Q2XVfKuYxdWKfQl7
LFfRaU8mKtmmtowlWonvRNEViwhuVq6qz1EBfXm9abP1izS4wZTz6mWBRBimcaep
S6hILE5znQ9wjOdkBbn54WZavjM1Wxbq+2vURNvm8CJPzN3tNNKUg2AJHJlcLswd
`pragma protect end_protected
