`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
clZsKU+xOztq/MzK7gujhGspevguNxlujm6uoGcuJXdJuwkcTgUfkYN6IGBSLb4J
j1iM6SKjaCQUNbJPGVMHbbLwWaoJY2/g14ZHr6p6DwGfAuOwLo3CIke00Glqqvkr
vqQ9xB/YjrZhAEA718Bs4IkUD7gIQAIuAk4SRnJwBj4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5072)
+QyTICdfy1qa9CCK6y79TRtEe8NhXMjRjYnytabrguMjbm+iGRqYdYx70dFZzf3J
q4FkahP8O2aqDsW2OCr/RH/38AWcKs7h3Di0c8iPkq8OsItMi/jegJiVEaEEP2po
JppvzUGu08RdNmy65kWMvV6QKVJmeHvC/lqshYlr1HSK7ZDfdAdCUZ0toVnHqj54
r92HVWD4ZP52dz2gdsUexl7M8Iz40qD4QmSy/wDUJqttZzm8y3QlACU4/4M4uIEl
coNFcVG+atX024HlYavWlj1Nmk3uI9N42K3FZrzrJkM4q7tCWswV6jA14jH/xQgo
myAQUrJyWZwZ40F55a/3TSW24FapoqC7dK1DTExwfPbyrEiVIRdwB3ewcLCfvSJP
stRp2g5RMOvex/70/JFPPwOdP6Mf3aL4y3y54kMtHHLXJbTBldSvbklI1Lk/7M0h
jBuTNxh2pXScdb/55kV/mg3NbhXibjYXxjCEZcpeY1CX2ytV9p8XJ83+anjtrWe1
gleL2XaXVsBs3liY8ydNvgHp4KYN2w9Wd7iTbAOegsGiLkOaoCAlMEfp/hj96QfP
GgR08yClqcJ2K76xMnbjw+KRXTiLXjGS31v8KuKKIGRjE0mmTjRhPcBqX0LT8Ru4
aeGOQ2+4oXUiRoxjTWDBN20aUa9dGL0OUPwKQJh3gjS9uVekpVV9s3tf2VfueS/+
JCjJOz4Cv0hqBsolUr5ixL6DfaGV8W6oWB8jFUOCjqJ4WBuGRIayfgBeD10GAQUz
9xLA78ye18TgopVT87BRe9KW5gnaEphvlMyPHjmuAnZErLmcblzLcCaF2c+G8XBY
ct2DhbJn1iGLq/+Mb3QeqJa1Sr4KOxNVV1Les6VXuxC35hlmYWke3rmV8EdhURD5
+vTx2i/2v/8U6IOvcRbAlXi8QzVlUoqu/XAGMsK2X6GAhM6rVxHgy1/WB0GAw+rn
ENqgBud0Y1V1TLP9slVND7rJX9440KO6FSGnR+nwX4k2csMCh2VT366o1foS+jgy
zkRGdeolfBcQNcUk87uKn1MLNlwy88Av8PbwU4ZihZIMTA58SSKU/fqS3+wWDu8k
I5GMaUK7j1WnKc3qaPGHNR4gwex8113CjVq0TNH422S1uBc603N2XLN343ZZRswq
TbmDgAc/P/6lYNfUk7kFV9Cjt4vC+/rBErv4cSwc7XrECJDVt0IFzU4GaZbWmOZ9
OebLeI0AU0M8lj9NYyJthWUez2CQ02n/wZ83PZ//5bXmGsgpTiabeZnPTDEYs5tV
Py/zg/ltP/kKTnmkLv4/uhk/EfzC9bCIo4kBr5GpobzsbwsSihRU135Lgdlq72dS
nxPQP4exhU5NaH9z4N7mYeBEqmCNJLnWS67jRvV8WGskUzfnW5GkogGQuRBN+4VB
AlMWEBP2KGKa2JdNeDfR+KJVT7mL+thR9/97FHr1sprtWKRBJY25B8lH85FZUL3r
cmWaoeGfBS/iGmgyaypj5Xz0efpS9Z6GxPlVm7k0f3yQvqd7Pc+6f4EulTMSmm9X
KhbWRB6hoalwzBlCUva2N1NsnWyMXrkp2qr0KMMAOSrBQ8rLZND5RpopxoZ57GZ4
X3DVQMPwCCLBDT11qDcufJCSwWjis/zCpCpaqJZuJ5f7op7PMWLzOJXA/fxTl2hW
iIPdeYfx48w1B1b4JgOaKWny+mHwzUKjVS4Ob1d/9gsibnne9m0GrHTDK/q6EF8p
Pv7OFpbqmXrSFAnVOknMBqiWruxt9a4ryRqM2PJrWecgX+HLbvlU99eqM/XyZKDB
PcC85rbA3NbdQu5nbBsqXutfqFykqf2B/k6CiohqIpHxYm54fvwtJlu0xDW8CeGH
mLZSsR1J1P27h6ocyfPSyMj7E5ZDNtcYggkRt7EROj+9TKq9SoOoBze6rbX31Ibf
bcz+vB/pUUOJDWYsfj+u8HsV3am9GCCgR/ZPGDWMzPKW97ITl6pNop9zdBrelOt8
zHB1CiP8CVfEVGL0Qd2+eR+Gq3/Wc/6tYu0G2Dnlqgh7ynShO1z5MMhiwsuOJoo7
gUTYbNdndfq1UM6gxZ/z6XQDEPWpp+kqGFov0QS+4kg+Ydpk0jdPudyQHAMlR3IE
qsptMdcEIJBU6LAq0qsJyKpwR4pbCLqgjHmsgbYyBbQBopOXHlPox1j0ymcNWUa9
OIO9X6H5mBte2eXdbjhDSWZMagUn6uYuYTUw1SAa9fZGDEtztMGYXkYIV040oKc+
UxXcyk64VCmxfk58Z9lKFfYYd9MHKkPmNZ6kP+wM4ZxhD9jJZl2AbgPCjupuL5oH
Ih5lBc4oywIQzpmak+R9yG0vAqa0QhmnVlU+xSil7KBohQwQJ0YMhBDpLIb9M+Ew
cSentwieR0w4nafr6t/9Eyrdh6tHmBTEJAWo97Gv05ovzr+S+muI9YPKQuxkv17p
BoYql/jfna157tNRfGRrzA2EFmpIrRWWdqyDa0ggnCsaUmyoAVijv3bpZjRffa63
FFeSP3/40Ggl+OsPCZT+Hllvtl9Nv///uPm75ntGkRRJeEgsPWtQ78iNPi3n9DM2
uwYKKtYK9gzvsdmTLHnWB/vP4RNvewOG6j/hrHSzRLi9AoEz0/Az4LnFH6//9Zhk
zNlrKNtH3hKSzuh8R1Wy/il9xI2O79nF5pd4N29kQBpsEWbx2WBmd/P747IPklD4
ZqChXHpMPbpT/yRGpsvs6yVQdEvGShkkPFSiT70chwzjE3rL5sOniKiI1wBlKzBU
eGjk0V8hcZ4UGzMjt0CKp7NUynkruhtMwkZL3P44im+6vEC8kGkXBwMGeic5Vhvy
9BLe/vqr82F4uYSKnXOuy5zqSy2+Nj1DWEMmrBw6uvsADtQmyoG00ml27k4dwAij
pdXP3uq658DE+nZFMjB0ZoCaACwZDUsmmxxsFbwFVT2msx23TvQzU56XTIJFwP7i
iET9CcSRTUA+cqgNItf7rVhEhcvD38vRnVUeittz+QNa501RejMUGap5dRCmeQ/p
OyJRK93r6UT10bZtJawXGgtRvuY/3qNobkoYyfcxJHyRYz82SqFTMxlm4WtEWeF0
tOwNZmmCWquoomJPZx9tzCx0LKIYSkDu0BW0m8zVS/kz3GqYY/B44c5TyxGfj57H
LrhdQG+3cua8KpTY0pJgj0IBa67JbyQxFKyEm4Wr6JL/cymJ20v2+kh9/wGthzo1
5bld5om6ZIGvVlONnPMgd94gnCZZEH7thKRycr0ueOrQ90CNByfw4lqiu7e4BkLv
9mP87hzcS7t1pHFbXOxyu+5YbTcMApj26QzLrztbUxW6cPq7WJMFZuQBMQZehqW5
M9KGYLb5ladryRNpQWctUg9Ii572jnsRGjbiNAtXQlwowVDhrMk+c0L72j51Dmfv
kMYB9NLmHX6UJfTQxO1u4RVgrP0ppiUwjODYxTd5A3h1pVjFvH81l3U19KrBF6hE
c6TZmCAkcQL8YqOUKXv0bgoCxpOZghKtv6fTKrAZW+7W/Gky+b5jaO9+eSpqlJCp
7RsYiOesZNPPq2PLVwDEceVb0rwyNr3Xy8acp7Ai7t8QC20tQuZuKbmeJUIGbmaq
NxSES1jNFxtqT1viaD7t0qc7bDkuRi5H6J/tnXsnfOp6hUlu+LGUpRYB3lvS7beB
iX1E2NUaOuFziQEPYSwqNr8bxR21vqzKxsZ7eRc2M9DJfEkJiH/krgrOrBz5ilz6
zk0FB4g47mapN7IIk+wCx8A11VpbWyH5axGMGOo7TXlngzR7M52HpvhltYYCr9ke
AMgv70Y9uUUIQNkdokgvgxL400CzWeVjbgoW+eucMnAhkNiB6dUlg+Oj9TsYXR2g
3W9S8opAI+mgAbIvBDna5aniEXsZYyqSJmkiOuSW635m1LpgrT/awXaYWlokBI/R
+P2A/eRrZQTwfmajG6Bdv3M47yc6A+lkIIsksMAsYGYGEAVZDj2+kvnXKZthWQHg
I6RmevGCS4nUOTioli+SonHTLvz3VmSulc6d1ix4wvb03RTTp8vbH8XYfU4I7iw/
F9wJON9fBYOixxUwF3mFtrY2Kd/tDbNgUaKiewnxuxh9osk6BowwuvJ01ZY5OVkR
lHJknLAYVQJG+Vi9nUZQJJvfeRjS8UGF7fv8RPHCVwFmO9LkXrE6pWJGMMsNRGy4
vktgNQoYEVYM7zly8yf+KjP44b9b2/Ty8Gs6dglKcyksnHnTU4LRIqZY5lE4SjU1
K5bVSQIrjp27F5EJVVgODweFuq7Bxz7lZlvBd23+DAim48/F/GLwbwyshj825ILZ
71wR+H2AkPiI0ciI2vhdxFA4T/dqaeu+oS65p/MwcMSfwMKL1MZ7Xj016EWozvXm
/coaqmHRFaQOsKA54lM9zhfBPF4R2RjO2FnNzbLCrgjnP3Bxs5bERrO/KzilpgFt
I4IWeLlzUDGo9tFApcl9zwvqypn6gBhGOaz5sd9uqYtEsiA6zeFPcbsufK4bJuaJ
vWkV7shO7W+q+jS9Bn6uMqKYJl/zr3Qsb/DJoF6OdNPAcSI6sNZ4wcJ6c6bJg/b9
4IThxXGiqamiiX9RYYZLyC0Vm9lNjXebAXQmU9k93HgbM4wg7tlaEAGTtF8+xtDb
JfHj7jWMlqkNc+Y3dPMqrCBZu97wp2n8LwV0PXst/0/mjicjwweD7UacUMGmP2wv
CpigvDFl1BfbI/zObKkiWEBWxG+rEA89xBSbiFbzJIqf3vMXLMT4cfimubCN7pqz
ohk88bxMJcLZBYiL5BpW/nPotQhxCXh8jE9+FiyOG+nsSXtpPs6hiZ1eNUTcUZfu
cRyP5h/EBrZnAsHQ5ARTYscU+SkC2gUkTbbn15h3yC2/L9PVYvQNKwYDl8E4WWPi
LmD/iIQJM/un11fxK25Wu5fi0RYNNRJ5IDTE0y098YW6MzlzagbhN22Nl2jYJY3x
Q+4oWhREhJmMV/ZpMbOsmmBYlRORuMP0lheKOzzi5+LfGkOUaWWwpf+9M81BI1RE
80RgMrT/jXM1FCrBeVhyvTsW0oXKHIr/RI3ipH91mBqE4L8CtBjZBokbVGjEkF8u
uEn5gh3KuIekZ7DLPYoP9yoI4OAfzL0xS8tXEx9no/6YADmIJrPQcGeUbq3rxUDR
9WQqzRYWtvl7b5U3hDMposYjnYnFuFUjp2c3WVuUHvUzIq4ccyJ7rGOEJHmZsWsn
5jwZGgqU4oBmKXURgH1yoz+MPBzi2wDgQqhx5a8zoZroWUrDnL3swbe7+f9AP9MK
IRMW0xl/7Sm4aQyKp6arneXQR4T3yVY3GcdwlXhrYJYEviWZw9fOAI2eqJu266Uj
Yp20MDpuWzfuRxbg6o8JWasSHJBDrovHSaeiaGPcZvUECLxe9vsLOPdkDpbNrxTD
jz+B7IJFEzMRDKtSYwgbmAM16dwSJv7IN7szcUQTINqaFoLtJ5i1l5YAHMjVvehs
/4Niv0wIUbh961preLg+UG/NoOyzcVQMHxFODgUdnmV7KghX4Cl4CMTxXsR1j9SD
Qd3IbKIHKexroe3LllP3yPUPeq/fBCFzd7zU0ysRSoorvhLHXhK+UgeCDcj7aQ/q
8JMKWtujdFysgy+INowqRxz+0OAv7lZ3nBE4Umz9yn29iEWg4vKGP5QMXerit8fw
8hm6tNrnip+lhAiAdomJOGmG19qv9RARqVgpEav3OeH0MmW8IPiJcSIXmh6TWe6a
GZVDawPMTsF09/pijt5N/6eoGXPssHfa0oeEg2NwbmJH9Uhl1PtpDe6aOgLNPsla
4qeyc3AQ7E82yBPb9HUujE3Zxx6MvUTLuFUQKVg4ineDIB/GpA49+xqx1wzEmBVD
J8w+EY9IpSAjHAhGGUczS4x/0ktO6dSsSWPnPOTCpdNwyS7UeMXfPD3Mmj+gNl1w
dVR9qku6uOSzclWXnfGOjtuI2r6fshMY9MkHh6nSg4u1eVrDC5UqUaxVj7jmIVhd
9ZgmLJLaJq8jlUOQ4KxMLbKeJn2vFf0730UhQAp32BgqRVRj2qHV3Wk9jCYRwHNM
4RJcnIKz5qwHZDHL9KEHaEW9UCsyL9m3RjlVqBimbumGj9N+gsQSFIYKDekXWSl0
ycbZ2BLac7Rr9MQSKUE/zd9wovz8D/Hxc4QWy3IwfbsX/5l5859VbroO1AQUhu2I
FwX+Vz/jf+RmjdYgsK/pQ1DC9tDMjyk+6m9mfDNjOddFF4BN4zTxbcdceXflgIEn
h3Y+ihraFXbweNfgzZQIg2nrP3Y22Hxt5keAy4Jct7SW843lK5mOgjBnW0gEeOwq
YvEzh/ITsA74ETy1R/+mOJsPGgL8jPJYP1e5v9wklzisSV7pnueMh0+Ek8NXHHR4
vFQDjrZcAOvJrQ55Stbuau/AQLkGDQheJ/nGIRvZImTIqZs+7z66rtXHiYxRTf8D
A0fKU4KJQPdXuY1kuo9CdKvHnnDLuT7O+skL6JFCyLTBzTj4WZFKTyrBxUfIICiK
TpuJZ23VtPoLYDN0WWjB17y74w+YdN6nkSylDpDtSbzYBKy9u1KZPVpIns5IBj0F
XEuLyK18STLeSGYxwMyWTVVJmiVrqitlZ6SzJpQ/qhJp95xIwc1EvVRUfprT1nyc
l/bIeXRm0MeAYWBhNl5Pc2L8wO5ZtPpvjo+suSCShaSDNUs5ZQYY/aN0edc5TmBL
CsloR5TRArp+TdCWSdH2rNZwcefTmSZ9XcuC8Pap4+VIJ8WecF2nE1AHUaHxUPFz
ZqRYDMkLw8EFSPjmKwXjAJcPOKoaUA2tgANYSsAPB1g=
`pragma protect end_protected
