`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AkyaxrdsJqq7F4QC1lorAt+gue35qJK1AlG2POJnMH63eIs09lLXQ/eAHg7xG+wc
bYrMM+qGGB1w9tu4FTAfULNT3cLkJvnI+7Vg8AzDlfOpySNdl6Q//9spdRdWYZc0
+bVLOxd9e4kMS5WCl6c8agGV0Jj6xr6Oxk0+BEvRoJk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11072)
9+ppUBsrJiF3ZPs0QOr6wPKR8AmIAyNbhQCaIcR2Thn7No1Aw20Y2yo77PFhnZIQ
mYk2D6lYBMA85nWjuqm3isbN+G2lBQvlDfAsg3Y5VQkz/7CYONWj4J73OIeEOKw7
tp2V92AWZKZkVqsvk2J+X3Ja78WNii/DlObiESRPsMxKF6zkhcPgDL5ve1IrztXe
S8PNL9/iJRcQZsKuMZecYaw6H0DIWsrzV8vCA9L0aoeTx3isGIg63yIxo+tDJuPB
OQbMkgT3SchEKosAhHYuPQwr22gV4/7nodLrMRrhDXCg7QZGj98aOdrn+1EANeUB
RtYRPMLUPs/P73H0CheyKqew2t4znoURpRnPaNZT5SBv0DVwXQ0hs9TzaF66gmnK
dZubRYTDkzI8RHF+jkZ+y2eExTRwa65yYXj5MclKznIDigWQIafNcDL9UXMb+/u+
S5j3+t9ah/mD/2xw5WA+VmSac4S5cXYZrhF/efj2WlL0pz1dJXwR+6dZlAsjbCb6
7RezRZrJyB05LC7pXOgwpdhOj111hefKH2alQtHGzcZl5NCK4pGKubLgt6AL3VwL
rWM5htm2a7uWOBxl7p989xGQGgpwl/Pv9NrQLaVK6Q8B4PygiwMupCs+md/2NwNO
bjE/0CktwJ6weBlJ3QL5tYYqsZKlhEloWkN5wuokrG0bBzD1g2QD2k8a4YX96lOP
hozPD3FNp0TkI7uLLUhEgWZo5et/K5SlVYpO/FEkkliuXn9fLiIzi4s9FIcqzRG+
MEmHX75yd+rKG3GKwWYND7lxcy2omIDrfVtO5noqrd55P/5dr8ojQIxF0RtyCCIQ
ziu6aenQ2FKcGfVXZwvw/bhiWDtohG6cCe4XGdSgoJWre1Y4Untc84JS01Ck3Y4w
OeEph/Ib73PS6rRN6sR0JKiXzErYCZqrpvVVu+kXQIx/kVWVFjVmKRY3959dkyIv
7bUB5eBQh/UZOekoClIISHkL8ZUObudYZPM3ENPRW8WBkNXYe+yj3GAaqohMYMRE
/tE5+CrCpx5MI5ZzPHh0r+ijezqUKeFzYvfievs7YFZ7UvwhlIb8QF+r7+GsKqxN
S+LoKsXFsjVQQMZ7cSZE1UB5dM5OHYFWRDVyrU4uyd4lW1QIVmD3t3f014oi+LIs
wG/kc+eIHTfzdTCWj9SKHP7VpkBWc5XQOGqsc8aeeo/P/rQYCyh47wv4qsoKDa4C
/CPqseI4kpYWXvoU764cjm/q+JTyyvVi3nYjACGe6/WefsFir5I3FTlhrSMAzmyo
gNm5RxEAiPFqirEg/Yp2qVCG9En0X9tXSNVr/AuL8m5RKMv+gIS1iIVEYMxZXUOS
sgXAhlbgtje5NjN6IEd1UgY1VbNRGxyJ+CdzTzvu5KAhKDICB09E5O4141h6yE5K
7bx7WavSKJ1X3zp2vV745/gb4DkKhPc5RJYsZQupsUw8lAHSNXbF+dQx/E1vrAXp
603W4NOv31KBDfWUiJnGLUzpVlcXoFUzYejQPNE1KgSzRMEtmLsm3KYXhqEqgPhe
tpjvYuLYNQCW4qqdkzmRN4lmNrXbgnTdHslxrOyeEuBvt96dEq7yirhbUVb+NsZj
mE8su8qtTEl6ExeoJQVEeSqgkQyfOQWr8xfw2kJEXpAqurEfCsvmOe41NS0bkcz/
TB2OhROEDpin8ZObRlx0dpy6gOoh0Dvi3Cmwg0230JvjpBPUED4mxndc0c+3Gr9V
76nXLl1NUGWZ/pgAb7fwZpC+sj22teOrBoCsI8gk/yRVcGMxZD7J0KgY0YjAoKUq
+XbtZuKdfUzb6P1xdxZRToRvlcFug6uGMzth5oDL0a1Gr6QuHtKFpeEjS8HBoMHM
7f0XbfqH9roU5HcP6bmRBpiQ2KuTaf+s2zO1CQKKGxqQ9m4mD7ttq4DIf0RZZCe6
5f/QmRAEzzZaOqDFqCUvAcIo9qbV2AVScZcLxCx7k3JLFyWojEzJmUR1limJBI3e
4ekPZtav9TEOGASAbO0slfos+nyEzr13DN6gyrisv8JTeRgBEPvMHc6+WoyyzCOY
IK38YrcKNqWFzmumLiVsF1ydp+45v5N0VMLcsyATfCz31VwscFGS6aCDqbSNXqEp
kHqXAysqSk+Uk8+bnbZI0RESYEW5S1A2Px0fIhZcDutq7lAU6OQuGkB3LqHsaLop
LVx7BCZMdpKCYwi8BK0pZYzormmh7AxN2+2mbz0MFcLG2MSqkBlYllv8UGrSkguG
Is1vda6HRv9BxlF/6LDBg8vepX/N86/dUsqg2bPz+LarElJ3iRXLWA+Vz7I7IPfw
4IqftV9mIUJ5gHS0AKM1I7ZmfnZHsPUd2bQdgX7acWD04F1oYwmLPvKUYzaERnJd
+u3M/Lj1GEgW9rHeHxy5WmlOU5rCj+L5pQtdJ7MwgRzn5J+qIC8snu30GZFVP0zl
yCbX5a7mxWzRQ+BDxA/5eIRgcLWfVtaOgseVLhxacBqdmugc24Fzo5Z2u5fywMtS
6xcYorlyWZfnBBt/Re5052apZR9wljAFqbnfJZjuz5WGg6096EmnHlOKeixgycXs
mTiq3F9eQllfLdb2fbeoYMKQDAbHcELpKcplxIVJwv/ctwyaj7zxGqDUkFZITf3z
SLtE0qJjMnNMDPEBPBZNAvibh9lFDFxvV7WNK0fxUdil+aSruyO0trmwGX2coGH2
9dhoMbz/psD3oTOG0iVtDcL3AdV9RduMCSHPB4IeajGAKpDmTIFEjCXGuNHB/Q0C
hFNMUH/GdyUBWc6qTJz3A6RItYDaGsh1snaRBlLvdhUcOzE05XXamxAiQzoYrGL9
kyIT6qMevvxIWLcforvQGMRvSGurpZo9DwcI2FtOKe7DhjSYZyemb70gvuVpQsxu
XO+vjPtxcISikrldiP47l7YwZyEX08gIGIFwzXbCxxm78Ijp9y6710t/vjjdUl2D
exvilC1H3NJbO6tzScoOfnjAeSuPXvBfXcC9jP+Vp1RDOUnCpM6YqmdTK29SFprL
hs+GLW+81N+iWd25OghFH3f3PMqu05XRf0yzj/ESWNJf6iHySxd+f9te/v8mgG1/
Csg2kZA8dsiVtOrG0PuvbTHpyBryULr26TsSU9tx1KqSL8vMuPalzGJeGbQld2XT
ijiYFXT3RacdRp3oUb4+dMkMGxGqAhIZlm4cV/rsOGi69XvmSuKUf6Id9bs2aL+e
ehOH2H2zp5yVvLX8bHzh7H67KgTY3yxfI7vUs3XuS29srMZS4JxB8WHufA6SSjU9
1fRSQ0bONybP+DoI4qSQB8dJCsN3PeVOCHGagpfwVeWt+iQcIVco6RkSyaeI/1Nz
9ejyB9WJ9WlhybXcREIUaGfq3Nwa46I+kBYzZJsQcS7xVfF/YleM77aXt1ZG21Kq
ZAgqFmLWisWMtw+7oFCJLoQYxCqFEULLc1uDmRbg/vGZ3eX/at4Z5flRov8IPy+E
l67gQ6gJp3EVKtQrtX0erHLcl2sew9C/aZpP3ftRtJoYow5inD4d2jLoMM2QZi0b
1C+CIjauOREhN0KudpBrklTafP/smw1svhOY1aoE2T1aAVTh/8Kbzfy559f/eo3S
yCyjtYugHGIVStEjQADyk1Cs2sJlc47UV6jLkgHt4GK0qZ5FiU6MU6Ud7qSjho8o
gYfd6O/ZJZOd/jFyC8ilqkkkmZNrYQGPEWg8Zvr/mgxwZfEbar6ynHMBsC4LY1dC
2ZK3O5qkI+T289G9mmYFDzSFfBXz5GVRZyPIaH1vhKU0Ow207hY31rnEEqBtqSTj
wuP6lsUDlUTPhpo8peTzuPpmsP6dR+i8mcv6Fc+RY18CRyeG1IS3oXLyjbUr46nz
gMoKYfAZNCvxKGH18SjAhPsMVJTm62Y+dg1aWRgcVyBKRKvWv18aB9YsUi9474ut
Mk0fCjZwBI2ROWtAHVyFJvkvbH1KK0+oK3b9FwjMCNz4FQFyBJKq2eoe2ZkdQGdg
cPcMWZ6/cbODCNottjUHsyeYwb7qKJFk3P83mtH0mTOq9OhNFOdF7t3rUINpXBgQ
b/gycPwAP5agwM73GoowucX8u8UbVfdJh94weWZYWfe3B9hKTQzr1adWyJgxBlsJ
xHYCLPxHuzEM5xdIMAoVvrZpXF66W2NqMgQU4fIHJHdFf8Keo4tTWUDdl1sQ7jBZ
UYSm7dwYDjbCtZbc/i79XVw83R/Tih0VZTkp8mj6jg+ZxJ0d8z6j0FkxUVOH6Y9y
ZHKpez/K1y8iSBPdlDJurOM/NxSzLScCpPcNm1NJHdNwBqPPK7WHyQWysoapneKI
k1kj6c5pDS2zQ0otLYn8b6tifao3XW3cGCO1cr7wazc4sf3daOFtaA+qFZDVfwmP
KQtxZqO7IDZlHiwLiIitCqphPJEkZ7OjqtkdZLCA+UrNgtbHUHAdQcYHevxueZYs
MkjD+ObXPudvVir+K80BeYnJlYKoHxpY4wI+hi5p04AYqY/tNAa+D7cGrSlyARI+
Tl/v9p1BwpN47MEp5BHWKT+ggsvV+Akx+pGNjrf7V5sHcVNTOhpftMzdZ61jvyHZ
sZFvuKWW7uZXYms8PACdQgJhR9mODOjgNxB5YarhDLMNL/ulxBeD+QfRqIAsb9dY
U1ohEZQu6MvGyGHKPhY6fM9zMWKFSn1yLyeK3h/hrqII1RnG4WVa1sqesjnGJE5o
0l+31D10DWHBE+ikHg3ATepKx+P52gJW3aFWtufO6rJ0S1GJevJ+ZraK2sCGFnRT
d9/sTH/hIzZuu/UKpVLyk2rSg8vg/nM25wVeVxi0vLRQ2r/KP6JPwOIfCsXispfG
g8dMpFDVwP9TOOdYAgksw/YZyrtCKVOJ7yvnSM+Odosg9EdiV9G0zi+BgfX9XY9J
130jN0C2Rzfj7vtBZSq0UP4zsZ3+q0g521WjuUlMGiNebICp+R04RoSqh9VAkoRC
GCf5vocPQs3kRPriD3CaFZqfSZPBKyWY7MeYtsIpgzM4sEdmcUnRVOvPYRWBxEqf
gWPDJ1k+CufwVM81F7oI8QxWRezMo2Qmz/FJ46dPn0PDMPRRYpg5YJ+Jo2QqLPW6
IV8wQ3FLDs7TLgLrNXSjB5DElp+jkFO6+Y5r/dMVPGUkR2sOq7qx+wFG+X6dnBCK
khsd188/0j5Bd9trK6Yif3NO4FiUMu5Syn45mC74Bw49q5DqlDgJZb7x4Vuuh9Ia
tovGnAjTLNbybfnAQxgYpmRSRMwgG0yjshUHp0E3ct3WekubARWJRCTsb5l9wgP4
7hrhSe5tZ1wTDe1q+xGacQ/gD/GSFCET0WPQPHeQmJ1AJUz3CD40dIqGG8h611K5
Bn2SKT78UFwdQ3kO4eFKBO29J9B+2IW7vDGxRIIfeEq3xmIiqACUFcl8G5luglcm
ZhTXsxl3gN7gORyGzfwrO7ofdN2u7vLuySxvihbHmqu61M6GFA2+BH3M0Rvk7Fig
cJS/SDnzKAoILfNFPNzNo3+Q0ZIpGQ+DSURocnHoot1Djemj79ZcN/8bRcHF1ivP
kxj7mY7Ty2vRxvZTWlO0JtQcSbPXwh+BAQ6/nL0mm3U2gpAxyCEd5HH7QwT62hQW
jxM7XprTOSLnohjmNyGzW6lmslJwPgStDbd3vW8xN2oIDpNNT4wXts3g1/aRrDi1
fkvZzNlJAur/LszbrYcN/l7PHu0ciftDv94BNj4XCf627L3UYYGTTWK03rDtDv7f
RA1vJ6b8BsGIMHjO9+SED3omM022p09CxmXERqD/cOKCvPg0NO3V9bZcGNC46THc
W0cnuJDAPs5nFY0Bs1U2bnmBGy3LEXiwenqoTFAzrBZs65tIDqHZ0mXCPrmNUNX/
Sqp9O+GGF849PC6nqULkOYFqvon03g3rCWb+t2kYEscdHzlUXEdabTGr65/tgNDt
1qmjHIfloBMLd1ipKRzzmljsgN1X+bZAI3H/G5CKlS/tPv4AJvl5nDGy+dMObTSo
cpap3vQFcCuHQUzuY+s5EZPpHfjwaNJNGvQf6SZBfk7gQbza07Tsgu5iEZ7U3XRg
KqxAxwfcTuRsexkgztGj90nK9TZXKP/YAMHQ1d0Ikjru3zSkz4XuIoQbiBsK8Z2k
dHVKWshy74dGc+npyV/cXXSQbFLXU9EEcMRK9iw515rpZtLhuL6QiZSI9Kguq/Yk
F+nxANEf46v71499znU6xBpdKTPtjSzexgRI1j3bpZw3TmlJH/nb6p7TN4NMSC03
yqSN2Z8mM88OAf3qrQ0P39/DhwyAQcOqzpYZsBuDk6SVdS3HGDO60wtNKY9RgXfi
d/dYpYxs5P7dgCtrQ6e0HmD6BRL40q6pUSjbzPqsN93F7Ni9vQqZD9+0RZGJ3AEP
f9+kLqSIizCpLESkvlAbDZBS1ezAsMd0jYeA0z3WovbIAlWl8aAk8MReyvQMHn5L
q6305x5aUruFT4m4CeZpd6g41mdtWSjteZ4UkY+b9tO48gZQfta4NL6vl9c05gpX
KQrWFrE0cdyvYCc7/AHkH4ee9kjZasn1CqbDyvNl3kbE6FpzNEovpEgNJrWIwug0
G+kP29tMOhnEAJ7B/uMHkJg+m7j0kyPe21qSRm29X+2XI/fyoXduKpC6vRHsuaHp
BNUNhHXWUfg3dCRyslp5WnjrtqPrB5VY7YfFqWH8wmErqCeqal63g7wwVmpSu5ya
6cjp+biOOfW7wjntDw4E7D2TjL85WOl/k4XPA54kpLHHb5ftab9A6zGvaAdCpSS6
tMqgTfV7/ssFJvEVCwhCPVy4R0MMB/hVf7f8jizc81BjiTIEkJ/6AYoebewkXVhQ
izwc3a7VyY0Lmn9ljyGjN+QGJzoJoTQDNZ8SGjDVDT/effwb/t+37HCPc5EN1g/P
QjbVswjvCeN+LXCAm6M1lCxsjyf8B+hk6Lmg0AOTmvMevFgSe9OWvkPjaXQ8jxzl
V7hq5Ha3MVqL14TgRLzZWo3vArS5Fs76u4umapG3jaeGbTEkHibSfxrRFHHbaf/M
l0gFVACIgqlnrBnaD1GzavjFxQHjjCLHY+AOT7os2AEbEHbMw5TCsNQvyTk99RfQ
MKvwG2rrPXMxO/2l9um3eJ+f6xHf3VTRZTWAZYKgn3TGxpd4G/fEXarJ4hUTtJwG
RfTACB1M1lk6dejRGB9vgUqbTISgG95e9CgWCXMuqJvaFzEk3SCr54H8w6mrwndK
Cl85RFGvLoyUOXEvZAq8KR/VAhevSMugq3albicdJKn/1ZXbI0RkcwYfnTfihkU8
fuqPZqlxuXF4vbbLtT6IIK+VL4IF7fvZIJzC8XReO7e2gkfK1yNHgIj3VaZ8O2jM
f27kW+z/tOWd1pQHtokj8AuXJCcMbU5m8Ldg/Jk3QupyahmQS2OdPdJOu6rMaM+J
MTkvSH6VgP9HCh7pf0Lj6ZK0BmhJ2KhkZzRTd0xiVUTaD4ULCCI63Kqx4oYKhUvt
n4321BrERNBBJ8eknKXvzZgLNQ3IPZPRUVsusaRi/aO+GAVg4SXt1A+4GejtQVk6
9Ap4SlUDcMpkfNdv2Y6KoXMMaES9lVZ2N9ZLppA+sHQBWqJ5wwK7Vf0UAMVbSnNZ
mknzQ1QYGFbKbVcEho2jA4S5AYqp30xm2STT7SGQAqBvmzjAMouOdIAF/pWhbwF7
HTnJ9JtuCQyxR74aZuA4jDxU8T8he3/PLZsR3W/D2sYWsV9Hm8btXSqFvDyJCGXE
d2AtLepT3r9wDMNDmihNt3laUS/JQ6wyvQBhzGb98VM0srNam1tXOvWqUkRMUEOX
xH6VmThigbe1ne67uRHZR8t76xnNco+0/4EdwYtaboBmIAc2pEgXUICBMB242iD/
/ZEzS0koWvSehnxKdwy3/SmX2jk81uxMJav8qTywEpAQrxdTiohX2vClbEuXz61Y
WheGcMzzedwfZRjgmlrwmwcaAjZsgk53oK13aFvPsR6SeBLuD564Q/cIMk7Rx3Xk
PShgcAiD14TfZFqHdsRpDJrpe40lDd9hRccnEFlEb8lnQm0vcnfly8oINRctnx4f
ACfLEbJBDleEM1ofgGIzELcsZ8/G3nsYBxW2Ms9LsrWFS13H0UND47H7zIyDmSh+
bOmIb+hlRAgaWjUkA5/i9p0Xe7d5Ec/9IIejBIf/YHI86M1vSY9Y2CoVlOy9Ooee
C/Wdpmhq+tGiwAQg9aLIyFJJrGqmynBxLusuH+BUBIgoOeGtOxx1x6+aYuRiHgoI
RJffuUQKba/DFdNnlTPkr8DYt5DLktJTRQI7tPisjag6aOBQ7HpBj4d9rz9qYy2w
0BaL0oSrx51QGkUnwH5lGffqj2s7Zd/+nWF/5TrWY9tPB7m+fJSyOMmg57kEgGoG
nMN+pARGAENIe1tqQav2RvkeoD6kf/+G9mHTYW1GijJ0mNA1vmUQp7fh6hKWvCbQ
nEDjrfJnkX2qOkkBestDyKpNll4z423v/sV908GUzgg000MeE5ee90YteA0gGXzp
XwQT0SAqwWhJpy/V2s2xq0bcekw/oXGMh4NiiN67xNTEe5PruCYEl0qNaXnPkGCG
NR3GlZH/VwFuyD/NNYEtfmOYCGATsB3SkGzk1jF4XSSx6F/VniH/Yu5Et3ijbpcO
1Jxast11ZRMkIM86rsgCZe21kxM0Tj7UYAEfJduv+HduP3I6oDdn8YbmBWL9f31k
fx2guQe79JeWX151oCdPjexjaGR7aoTNm5PI5M0HVynQoRGBGS+i4r2CxAFz0gIr
OumGJ/T+/UVDfP+f2nVSsHVeucY5vMMKGDuJek757pQ0X2KkaxI5gdfCoGfAuvLf
xplST7arPGoxoxPGpHc8IuzLYiYCLjXIdzEvd/UnCVPuyNLUJs8yFaGQpSrZL8U7
AS78KaXPss7BiXnfhrNn5dqOXLiIdA1cvujrLil/+DBguZHgiPtrjMjg3mhKrVE/
v8mh9Pk56gJ/10QO3JiNgsPK7qp8vmLvZOl9Fw8/BjVaxMACzmOftI2ipCO4FM/M
JeQzuO8A5EGDg/XqQg4Z/KKK/tYFpzy7XhrOrpVZ2W4zEfztzmIpd/paHybOcNUy
ztY7nCq/VpnEa5pODxvI092Kun6HZ3VZS3Sq1M4GxvwbYwC/qOAeqD8pEuSbBjzi
47r/Ob9SE87X+8tt1gOqY8qUYbvRnw46vncO45PHtw8j/2kzkEBvYJ3j0pRLsYJ4
KsIKwH+iEHHaILQv6yfNp1VkkgVNjsYtesqUH6h7H2+XhOOByNAJwPaoeOB2kesV
QKfqmxh6m66Y3+huexXkPuE3OmVQL1HU9PeD51Aes1+zYAKoV3OrhAcC58NfDetA
Jt+g6Uw+kpF0k10EUVmPr9F/ymLC/vRpakARx0b2JsVFW1H1j6W/hINwv7/g74pt
UEC8e2QsKnqlaviGg1XY8/J48GKZws3+bOeLIqIPezB5KquujtvpNbJe2wPm7Vgh
rh7P3P6qn5NHmurSSoYND29mOQ3dkLTbtLfkfdrodO6BebdSdffVov21LnPqe+aT
dnf9+PsPBtYcp4YWjLOl7ZvMCxt9icBdIo9r/8rxhCObiYLF2rAmPJac3S00agNK
97pwD6pbYObQ4aqrQ+00/mZKak+Mo2ilQ1vawFwOapcFATOcR7txVd87Bab/DcNN
BYsIPYZxHh7aIip0AknxFh0Gm8TMHxJU8lAORkC76N6wg4faU6HrmA/39iHRWpMF
oeg0F7bx7OWLbs+sK8Gctw8cJKCbTuqGdPRzFEBgQf5LwtFVLWfuwb5rQNj4sRAf
Lldd77SlkyShWD/UJj/055c3gjuj02t/W53nLztcz5OupTbKClazU0OsnbEDM0Ap
wDo5mtaNr4x/Kw8nNSIDhPqq77BvzMvepPcDQiE1JDGWLFOIp++X7l5q4E87So7z
tFVCGCxKUjMCuFuv4Ze7SLwIo7Oen9ULbeXBvloo2FMnpzK/E0SkzgcQ8IeoXmp1
NgoQHduye5TdjwNFnHpH646LUg6wzfjg2Jyt+bg/YynTVQ92kKw0I6i9jmKfezsS
mgIYXTiDdm/KQe8FcCIEBr+xAXcXFCY28+HctQczvGc42I6s612tHxk6DtLnH9N+
OEm2k64TJ5A8P9QW7RdGni06jRQAidoMYGfi4fW1AfV8YZdB7Twn4crBHRnhT6l4
78VHrlt8yaNVHh6ObH3Xp0G89xfyX8p82tXn/Jav0U+0/DQBvzlPN/GMd47ksonE
TvVC414ljX0CpByfxVr4KQwXYDi+wWdQeY+tsFfN1I7MbBOz7dWAbxKylyA8Z+8F
gMd6cpAzr7fP1NO9xdPSQQ11xTUuXCb3/3SMq1LVsY89yzGeBP7sv4TSCv6YVsLg
NZ7BkJBptPxZa8M6+YPA/flbqT7+3TnI7dX964f9drmI2qaxxHJk+VgE60Z9LiSh
XBnsjTcVlYPpgZ9MPaNftVqBi7aZg2wmFQdf8amUxjUlblJLBg28zkbgaCtU64Bc
lYnc5WOUHbDtblIhOdbe++IYqMoAXAEw9se5/JuQpeptcWhvq5HXM9GlwWbo3mK/
8Vy6hMwzG1TEA+ba9xiRCKQ/Ux0CMqZr0S76wfP90gAyFU8MEW+gGT9+xhhQKvSd
9FXf4H2wUTVcFMV//bjvcjUpA4Rdc3zbGq+gm/GDPhhM6wVRsJLHX9UUgS/TemLf
dlA2MbEYOrPTPJ7zQb186KR2SfMoCT7a7Z4pf2Ho/XnLEkRL8YSI5Yhyv9MQpTYN
J+7T6xY8kb0JAp0TmF5KtbMaiBaIRpSOPYNjZBVRMNWuIZWb0618AZ4GieFKHCXe
U2/1YQqODnxLXU3atU467fqbq01TLFW/xS1zG7cr/WylQgXIDsNKErtg6eRr7v/M
baSPXMTNHSHWk6TI83ip1p06Swsy4G8nD5sntBSG/P98vdF0stHLq4hONKE3zEv/
ybMQWdf94YeoCpJOHW1UW1nv58Syb/xb5YlDmR0nu0TFP20H4p78UTMog+rDyc02
QGYsfdxunpsxG68FC+kKv/BiTPsrughPziRqVhm9F+PWXzG/o553SMfPrWECr3pu
Z3O9NMWzfRHUWIdxXVckNRoX0M/ACBTX2+SdLMiPDvhEMG/gbqmTc8tj27hJJlSQ
+LJjELNj56pEmp1OfhMU/zpKDw/OkyeN0443v9pBJsuNW4JMIamaVG2rz/s5cccd
bRqNZz38xGM3cjSe8Uz1ZgfPNQZU2VSpz9YlOdWGOku2sCOlBXe1t2o7QGHipOrm
HtoWoTsPfuSC0t2llgBJcqeXVUU5XBG+WZErEPrcd9ZOQXiUHDA+oR+O+gaQbaOK
8lpZTWmbkxszdn8lcvDIs/0nPcjP3KiNNudUI73HNDjay3C/AVzFMEeDRPg2r0Ug
Sot1W7Vpa1aNr23O3obj1yXj0c/3Y2z9Kidc8/QZMIVuhQBnOjudESZhb2SteGzu
Y760EMsF7tBhnaXwQohSK4Kfrf0aQ6vnq+s7TJ41/E70UHGXy16g5O9YRJvH4xS5
6CMojzWwT0d/pRRzS/uMnzAvetHohL6ij2xVyo1sdpwvNxGNeIMgakiKeeuwGcwc
m2gvJpOSfWhUIa0i8plIpZ8nFD3RWmQ2ph8vI/2ToFmU4YZ3/P+AAbeY59urNb5N
pHn55y7fWu0rh2jvOiquCvkmRW5zEhmsVZzbYj1abRqgTOIt+sotdkTWanrV3hB8
2i082hb/wqvKH6t7rBAdmduKvKvoorLLUC8XF3ywfVvXzmT/gy29U//tsW8/osaD
4MZqxe7FvbLeGZaS1e4u6YBdIMJc/FNMRfFyFxB/E/s2kZRcsNE8YFAmHeYOJqLv
h922qTS7uEdUqgt/EpNLx9oxZ4c3eh8PSSYkjJnYJegJpXcBv2x83/bYQGyghU6l
Dq9MVg6My3T7LSGlSGi+09KAzFRD+4jD0yTZgnAmhGdrycDdzeRI3pLWjd+Uu18d
EGmygtL8Ca2qUrZ3PMhIZv0saHDZfcx12PfSLL7ZGdUjL6kug3NYtVyg0vqHPad4
k7fVjA5Qp7GFNKLxO5U+WDvYok2tbjpH6dxGD5N6siY2sFxJmpb0EcuZDFPuWSxJ
agBoErdquen7snR1KZyYZkYLVRF2pT3dTVdU+xL1ZoBMkNOAd5NaOvhGiRmLTy9a
Trnme8TmoVo6dCJwZNC/V9TGOZ722na4J8p7wC9uFubOgdH/kIWKyXlHirHXwzIi
1IAFiJY0B+7tbT7hkvbYwixf/fuVdd7yI38X6YJbhVwvx97eZNBWHbCtog/rS7lE
3sJ2A0i/CwLO5pD6BUOTtwePO8/cjqd+cky+0SUxptODOOAK0tTh8wKTaJq0z1A8
oennynvO57cIYxq8KMfHGVRuk0tXb2OlJlws5PUhRYBVn86IdXEyjcMtRsCY2b3Q
ynqfZCVNj6MTI8mTXWkitT4Snp0pRjXuQoFB5YQ9RluHPDQcmRjR1KLXVoPa97hK
/SY/WEvd1BdGblBVEpMOcUObTye03M6w+LhoLg1jzM91WXBGDIKRkWGEpoTvqW0w
BNU6qw5iiCO5VfX+DUELAN8UG7KV8/Cvy88HJl6Vf2Sz3U9r7D81wKsVElVxB2Fp
bTPr7kgt296RiZV7c3TcY9Ubc4kJ+ULSxAp42JGoQM6+VH0Dn3JBN325gANKYp2X
RXIr3EVwbnk8k/2Mh4tof+0L+GMbMRfFBJVwPSPITJsgNzE/0o62qHCx+Dvm8CJE
OePYDewuTd0y6Tpfh4eTfhPhoFwOJDK116bFfDUuXO5ZGYwVlC7DrgSw+lbPtYxV
D4zW/4KAp6YILolwJ10aFyR21uxYyfTxj5noSY6Ktj0VL0KnB+QkvWcnvkRGJd24
KtwvbLdHNA+uX+8tf2DN1am97I4OCF5XTyrBBOt0enLZlVa1+YD4X6T7Zul82POs
hXQApwZKu+g7R34kGLdzlbqZr09QxS5IbsBHcESo0fZnbAxOtxs3YwwYqHI6vEPu
F7LszBZbiwvpvaA3BldAa1C6o8ZqH0j42X0mGecLmUpxyFXYpTmpU5ElSaHjic77
TtGOl+GRHN1xjJSIEBBtcV5X6q1H14NXTAW8+NUbX+xl983hygE+vi0YX/8fZ3wj
NvfF9FGItauPCFPhuiZqaIZ2jhodvlOckr1axlxGQMwnuNFGxtue/VdJwmrzqDZf
I06jvFZkgSqHma+Kd++Su4iuPO3aSQw0GlBNYKqAaHhJ11trJd7MpSD/BbREcTKZ
bwXDjmZiaUS+tpTJVsCKtYJNC7/QoP+IRG71qtunttSP0uFBmDJbPd/rRgbk//5Y
2KoNEOT1BUETygof1hWJKXuFjpJ2h5c3+vDp/5Q2VJKBDcRBc6VvPDXkQnjF/Lou
0cwft5jGqsSLG9igqs9JAXGVV6YKbfDkSyvoRxhk4z+vTvce+OgxuPdDbViZ8EVj
tuqMWzl/5QNfCvIyPJ01rCIvL9PNb+dBQ7WCu4tDoUsvBXVz6vC/leydMZhydBUJ
4YkwsjHk2cS5Zpnoaa0uo+SDB1Yj7vLRipcyCfVoMVj1/miCA2DKrGNheyRiDBMK
wT0RKkY1pbsKF2Yf0vbW0GuKuf/2yx0TAiBXBVqE1GGoto+26bhDhVf3EC0X3IhT
SQtYzWeEZJhldDDxZO8tr8IgBeR4PO3resW2eMv4XbnzY2/+34l/2UHBtWoSGgfk
ex6qcBcaGQFrIIP2URvsB3aCYXGwpG87Ba6w0faw8LckcOJuxqT6wu6SLXWy9kCq
H3P6sSX24+fLAYm1c+Nm7hfzD9iFTPXZLJJzQAbLHglmz9/pNbHittK8SJ+D8vAB
AYeILW0LesuIfQkW1elhHAy377ZS4pefp9gC7PsQUedTYkqNhdgbqFn43xCWgsTC
m2fTUbdBwVzIowShogz08QlKCXnD+WSub6vH4VFGyxDYvN+705n9zpqV/Te7dzhU
WAGOrRhlAyPOxrpsiGrBrznxEQIWAuvMVCjQph+ecHb80a1Tl49H6Wrc25c6Q6pT
yQ21T+JzcKuD2HLpKW7PUqWAP4xBpG6Hpd/nzcWUq7BRuoWAA2ibeyvHRt3O3mHx
NDhhGDKwjd9ycRIxzzGx0EtbSKgpBDZA69kWTZb1twHQy7c/u8zrMrqOJO7Wu0t0
jqmQPOB6yQbHqka4/h2FLQMRVH1JkmYzZKDlDKxIqErl1N18gaigTxepWMTkZhX5
ElHNEtRA+APl/FdJyHYvGrZpCLvq3GDx+MHKvMMRavA97gewWKWtJLKSdX03YQTA
fhIvoF7BrkYHjDpLCE9cX0H/q9pnltj2o53ox8DcBFfdKvSoYJ3tA/GlZ+VbQd4t
2xfQssH6/JEi9oR6+5IkFCY/AV2WQAURMm0zvqRgFOV73VzmG5aU+jZe96yaW4ES
c3xY8ZZw1fMnQLRqN6TRud4NFBjIl8rpULNh92+dipFs2U9paHJ2p7ceZPrez1qA
BF+PQA2h54QTcs5g++fOx9pCbTAUtJM8isfR9egKBR0rXqLISbmHiOumtEXfguwS
bZ3b1bHGpDZL1Tz8lVmfVYQ+2HnGCX4G6bhRvqkPvI1RmiL9q+6Wcv5gMUbIvx72
gjOYH/bt7XTeJkppx41m/1Un/3j+G1Kk5kG+Y9jTzUicf9vzK1I1KFAlpFBrX9yu
0h2mDkT5R8vROYO9y2Psq0MmHBHe4XtPCVsgrUnR+6g1vfjm+0riimcTrwFYqUPx
pfEq45CnDJsuZxcSA8YMfeyU1a/ijbtO9PRVv4VZh/Z2HJDCe04D8kcjn1hTKzJ4
3T/GelXaPK4XATMCxmccUT6PXTfAsnUCBZBzLEOysqA=
`pragma protect end_protected
