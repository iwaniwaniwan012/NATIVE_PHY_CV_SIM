`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PGuf/utMkvzenF9WnKVFOUlIXXtaP3/2WyepRfKTjvoPEuC9dEYq7D4RDfCSN+K7
a4LLFYhx2pwk2D+iCBrMtRH4kQj6N3qXfcke9Yl/WZDPRxn/IX0CaVNSKuDqFuAO
n6uyB/O8jh1QXk4Tuo64QE1Yt8aL2w7YJHD0+Y0l+fc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3504)
jfs7b9xVFJlfw0iQDcDu2RCdYzk0qW4eOk/eJOZ5m9/OCD1rz+x1XoBduUg5T0CN
bEId0PnZvufNXFjFVb0MhEv8yIobeB0ErLuLtfyNk37DxwRfojAObLaxr8uz0rU+
1NimTxWG6xm8AvAxytcyLhT5JT9k0hvKavSMmEKNu/T13cJYyj/GchZEvUJxEbZW
HmZRXO12vLlFStEpD7vKCzZerH4HDsshHlcsvxEE1yEBYE93IChoqIrrGOQujJk1
ROqqdiMzuKbiCnzjXW/mlTtCGP5d7KkpojvN65sv/IjZYvU/YyeKbKhdrCZd6rNL
CYilzSVu8p9rI18YhAreQQ+xQwDfhbdOmq5j3IcFWV1sFLjrwJzmTiwoKWShx2nO
YJgc5qpWRwIM2ea9touebQfO2RJY/IUeL+r3jpd3IO/xQRte6gzrbPpLZrPiZ0Ds
GCvslFjjbQRcFNegXc5AfvPEF8Ns2PwAuDxxD3bq9ledNuDchPaofAKPIkpWd26u
em+77vVY7XdO4UpsjiGTsk2OExrxnsxlLGqQMrGgWq8VOIdvqJ+u0OxoYV+lQnQ2
j/0unZvuNVUiRlkykNu+a6iuDVMu7UbNTjUUFUn1k6LUoZIIdmfIDQsiJaueyTB7
20l91+i2umwOQvwMmYglzAzRI9Mm8TkYckHFB6+bhzXPuH5X9VYs3SVNahJObyo2
KCsdC4e0ZZgWeF3ULbN+iXFPgGvpm31s5lh5Z7GD3dm9jHofo7G+jY5/RB6yUwJU
jbleEvNbY1lyWsRLpPUUEzgXSMH+Oz5ITm0aseIS1Peiqg/bYluUrbP6YlgRyEa9
bRqgpTjqaIzYAtcYpib4biGpW3+u6jAlCpl/6qaYVzpgcs9fx+O+luuohYrM8+Fz
RCdGYJvOF945TMcQPRE+j100ic7Lh/qRGoFNNuv+qXMZbYxYPq6qJDMZuLqKHTOJ
slRunUTApIqpo0DAZlIdXIVve/XET4Oh9IlOgj2CSGQkn7Cj5rxF1WDnIsICVfr5
hkM6Vez7WtX/ejY8deYoQfW7SmNGP4YaIlcvUZbzf1gkxOAOILAd2XPkTAMiyz4T
MuyMUGLBxtROmdNQXCO3Pu7DxBIysB0ny843sgi/1vXQBpxv1fJNDlPAFHFsO675
lsVa45z7xsXDq+OC+tjBI4LA2rkqkPn0m0jYp9SshlL5yYTYLVICx0AMrNstuU6v
OvSKsUyyHZMFUO8bmHQmXwaW+kghSbv1cw1sxFAp1KutbonZl7gGM7FNJg0B24Q5
RsHb05SUsM1sZYqLk1nwNfAzAAy4qmdv7C8+WyMg2BA9puKjyZMQ3j1OMVSqcmFU
1rOkLgFyI+6uGBvWOhnO9CkH7udeAeit2NDT45InZ0LUUbChEUrMMBqFECxi7LAx
okw2HvCC8JeSkZPTbLjRVzP2IooftkCo7tj7CQDrxml6WPNAVgasf3EHvkef/Kt2
TzghlHQnaFpsmxNO2uW+dKBFUQzw6jIUrZYXi5wCTEmPDQJeZQmP2lrSFFISl02e
nUaj9cyf0sMMKbqw3aP9MR+ky7735Rrj+D6VEuYI9FgzftFylZv7Av2qR0mfNRNJ
qtB+xrfWBm/1vhPhjmLa4ClHOazC940AJBBnejHEb3KatqrAyHGam+D8jSWjIUwc
FSg0SWVRj+mAkgiWnhYF9vrMPpM+rklkVB+CE3nzAd7R99dPrnXZxDbnZIgmb2J4
L9/LqOZr4BFVTrgwDTazlrIirb1WcYlW1+UPs66aP2qiazLFpLW6tn2vcrJzJXfB
tR8aiPG+Hgv7aULkjEg/55R5erTxmWqfyk30XJXAppH8EafYPafTDXFuT9rJCY/V
qwZrC3Z8sMXn/LmKfllWpM2qWLFEoBKvwll8aLWd09gBzj4GTKIKCU+gRsMAX4/Y
krQfR9JpiqLpX3xryToBbj6it0fVhD7yPsRGHc1Iu/5YStWEbAWMThfMHSFCymaG
NsFV8OpcTsjaj3kyqhoB/Dt0T8RZcYFttU4ZK4gunHNB9QSoVPDTBOIpZZvPH8hR
eGB1V0y8Cycag9gev63gpYM5+Vnn5yCtMQeeS5T4z0tKJwamy1PjPICX9ooOXKLE
WeHC271I35j87K5bzlRy8+P2cwwHgiysqT5VItQ8FyqPCqYStsYampBJtZte0Np4
2cptKA4Q9Ru1RQbCpJNZQGNOeLp4akXAug42WH09gQLugZ6MMyCDSZR83CKlb6tS
mWNYU1xGn8mFnMW3HPPLy0NLa9T9/FibCRLWarbYgwvNDLUff+sBfprHFh7EN/Tc
p1xGE73kqDRvKer8rm+6KjpqLylSRWZ5m2Y4YSqJ0XB2y51ztvpSvIqHBmgayBrU
5dG9zbK/OIjFqR7PGysbzsreGXA1Z15OPbQ40r9m7XcemU59j0g2aI/IEdSuOkAA
hLJGDqNt+U2lAgA462leKziPOn/Rk+gjwgNhfCG72V8TQEU8UaxXWuQVJMn2HQBF
dBh7BvTGDvboFUHe4j0/D1o2d+ugYY5DPD4y58fevUw6Trxgnb1sd1BijCQxhj+k
6Jez8r4OfEAmgaW/mCwq/A5ee0qaBXJNHHx6Ci0t1P52XDbG0E0juOU1THunnBVi
iUE4oKI4sOF6w7zSConmH4DLICsr6OM2Gch4izi85yqJ6CzG/HrSGxj5yoMbbgD/
Z1WdzslGT8Y04S5M3l+hMNHhFzllcX2p5SGOvVcCyvRhYX1IS/dKZJl5eudsUHbI
FsQuxXGFP4cV7z9g0OaQSGSzmOZ3mBxkownc4av0lU+tRVFU9fNhuagKY2BkpMvi
anHbL57vom4xJ80ANkPvC3gXfnOaEykPnqvegIiBqVopHrCc46d10Zio9cWFESyh
o9NAwe1Y79M4cwXP0ne1T84pP4MZli0aEvJZc0HlkGtebSgNAhAAc/zdlZuB5t8O
aRaePRVp2aqkLpDQasZWmYGqaVbSg83M9eGZqHp2TepRm3wiM/k81VSFfC+JGutT
+nExLr3ux1Eb7C97bAD14bJorEc4j8ja2UmmSMHPpAwCjSPm/DG3/Tg5HrG0sgAg
MK6V5pXDoEKhG91bnVxC28yUyKbc9PeyOU560NNdUf6lbs2cmrC2B2ubN9rafs67
rVoMGM3QHLEDdhXkYMk7j+32qL+EMmfpSJg2Y9Es28shTDf+Kzu364pSfNnup1l/
s0d9Oam/66gVeZJ2RPUKAhzMU5PqBW4bQLN8ouF2ZPk76ubI2Oyg9yQEUP8ATFe3
VRDYVWiL0MH547aZydlY3kBmqUfOInl141J8RXoUewLAeaBmArr5Bzf2498DPvqY
6zfTFDALIMxZ8PqP64C4BrbMHR4kvRCYWr5Qa0Ano5Nce0T8Etni7vlahL+7YEXs
yQuEGpC6vaGlV30plqXMxfdvuUXp/OiBGKgq3f7jrTq+unn1OpUi3+SUeccksndH
RReRdev0tYK6b1hCnonQHI2WQjXZYtXb4XjuVt1470JDl/u1Vz+eXYvjovKDdCKk
7kEos7P0tfUj2SH7gcG2Gal1t4Zb0XHkxR51//9YlxH5nzQFMKTe0kvro1u1eG/5
UDllG7PKJ47YYu2yfBgv6T71UNkWG4aC9bmucl/Jv8B/eQ0RLPylgZ3UNZzCkq33
Fif0wX84CCfAZEsNe3pc2PP+tQaM5HMiQMjzgi2jan7ybMdzhF6FP6eSflc83msG
8fqdcb01+pDxpC3QXP4XyKC+9NGXYuM7LKGDazAbSGewrvZd/a9FaDA1xA+6Ojbv
Ba3y1a+wxT8JFmJhXWZV29kJRT86Sk1gXPEfjbnrXbgc56Dtu49+x50pswPznkDd
h2itZhWY9e3xVj3AKtADbpGyFURqji6sPkvcVfqpWep/KkNKEpjLv63Fw+ZGzoCt
4jESNiX9oS8A+rnNj2eC+f+7LH72OCZQcDPh9NWzLNjPt+VPYSnftsXKnHkCFu/Q
Tn84knCJzJKtfk8Gq6vIbLPU+09dW65AGWdLnU4iWLKTVtgJ+OC/uiKbGbs3pe6G
K8sfXXUpzIGCCKLBAJuZVZLpPT5FB1gi0idBKoFrrISNmoMKcCk0INnBwU40SiGS
w/KDYqfxMJmS5HccFr2blw5zIuBOqi5wu5sULUd3PBCHeELWCpQFy8a2zxOQZT15
9pzGQ1FPRdM3ap8k3Ja7fN7ThYvsO5qPKtXXTFrd0JRqwk61xEvXKc10wuCeBIWm
Ni3GrdGicl+eQTmnn5i6dhrGJwJAtbDqn2/zJIrqXNglU2qIYFMdjR3dYAB/fWM6
SdWIrntHcrdOdI7BvCgK3FVxqZm7OEICnhmMYh5CmMLvl26Uw5jPAx6SfwcfqXuw
ZiyhPveaHmlevClSS3IpkSVZg50v0r45hbRMjkZvn7ShG0c9vJwJGmbVIXhXk6Da
voqw6niU2esHeeUp8coEEeHy9K4591pMsSHRjLyw668LyeAem/agxap9fVuN+yQf
+fF8jYFlYqffEGeUIBrQZZCwPJJL8Gj4OxA30jv1tn6WYak9OPE08bX3+9xIEma5
yEMUBMpVMySEtj7WOps3lykzKMRAqOE6rHW82CUNH5S8sFrbdGP+KBZCeRK86xxI
VnImtNQedo9mOMBYMhs0ZD+WSCBkGnPzfsFA1yPytnPAsocYo2RchWgG4+ks6KLb
`pragma protect end_protected
