`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IYHQJIzTK96nlx9FJlkYcYCOXVVroeN5YTdZl0JcePIpZ+YuBPqvrr7f4ethl3Rf
AZPQdYqTa2LBA5Kea18Beqvg+cBy+vT2R9f9yc6uo1GPrDcFx+9aKdzUwX4yMfrA
2OL/Bl0AFrUdB79Zgw2RYnJwTlf6XzNGOWT0EzSKLK4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5184)
SCHTDgH/pvp2Fk0xM9fZSzz4jjbZtQOXItrZ/1QQcugbt+E710YPYZfur8QvByTx
ol90OzOGO3eIzqsSgksww/MlXbcY4w6VmdV0NELTKqWGR+ALkxW1136mNxijAApI
3yVCUxn3MGgNeAN+gWMZgDWOnUquaV4Dqh/DsOSNu9gg7WKj3Pes6I0t6o1WYGFz
wR9GrXuSDIoksFBHXl2w03OMuAlglK7mPrKm/Hxoj+nTRi1siZJysP5XLYqKUoB9
7Wd5+4W+y3qN0WK8zDeBhX1LhWlJkuR3qa075iQshqusYP9xrHVort2U+ambn8It
T3HmXoRagWMxF3Ti96JTHx4sjWgLCmLZfGbkq2K/0IhTQQnM8IlunEamxPlhU2+C
pucSwP7eUuqC+fgU3dfKZvHiOwuHc7Otj8RPwlsjllXQioPqGahADzbi0aAFj5ds
2wYVAKZzGVXSz1xH2zNUAZOLZjhFDRz8CYJ8miGR6ewC0Sp0aoETsJ3XZbA/6PTr
fK1c3CA/0yNk0uLbvqwab0bjSTufaymiPII+d0+c2uupNuZutFtQLb4mNaFu0+TK
q2fI29UNgMsrOx7qfBJn9wjWoGLZB+5RrsHEJuzubnFix73ZFHOt8+ZiKTc24xzT
k8ugnVcQqF89d8nT/gXq/ghlGW7KpOKBZOyv519AETgxQwCHNG2+qLtvcKPstQoC
4pNQheC/nfTJ/uWBA+TEgvuxLKuPY31CHihw7cEP4nGPZBnwBbKYK4Bzvx1FTeuT
Pg9lOP6wJ4ZPz8buXaIFe5KC/DAKDc2NV+ma6M8IzkVx1O/qwoxxzjYI7mBAON+H
TZgGpYJe1jFP0Flvl5S64HIL9pXl+l5lrsqlGxGZ4//f6BNn/kl5IiFkklrkXyFb
MoeQncfN+l2TbRVE2zg9nGnA1yIOC5epvHKj/9D5k/oFH9RT37kfG7D+1ajMfMYk
30m32RKyPPoFXvNez9pIhxYMC5uPmetaWEAcz8RXRmHh0BTqYkVcGQO6sJaA9Oj1
zYRoysSNIA7f4asbMUQ6xOirnqaO3vnQNL+7S7AvbMDc1ZtFYfY5zVz/6F/BKBNH
UEzz3bIZxsJerAJqXWFWVlJUsk1vb9yeTOdsWP+p8Sx1NWaK/fpdhhYQYDJ15qJx
CGqdd8tNny3kUKhY1d1Ip33WSCAgQw5ajmqI25JEi/jnr0TZlmSMUMkzlFATj8F4
F1LD4me30awwxIa6QTx0xLfXbFsa8jM1SAPlwrGpUrHau+3cu83O745o07HkqjSU
wi/Gw9EbGfriepkBSUV4tDq825FCEq3E9ZnAcxrsNYgJggA2WjGO4zJXwNTwHMS4
0pojf68QqhWyywAH8EpjXSwbzMZrfe2MWIYLk81Pji8WIXO7jIMB+4QZ4J6uXlCu
1JAT9xMJ5AdAb56MvqYtaMiWU+QMOhkt2erqxP2Yswci4k2C3QePi5s11zR4pic9
BtfoiYcEYbgIiVwswEfEv2Ocxme+69rvl5ByBu8scDZ864eQmivWEsAztRVSdcL9
Q940nNFm+ufjIU6mmVlbYPJ5tSoQODGvEBJUvVyvH+vx4atA4M27w5gzORp0LIMP
TVZyWJM8zZOaLmleXpX+N5/iAd4fNQgYwJezo6ezNN4KaBn/lV4TgY8dV6Au7OSq
ShLSqsVKPfS1Gn7O9IFNUnfXWLTyh6lytYrstIioPY+gE16cEWHknLy9vn7w7sQ1
ejoDWx1BSgXfduUTGi3gFlWphN7ZX+TLvMBEmqsYBN0afgr6iqPhsmauOQkfO4Ai
un/nJ6GNWLwL2g5YEKw8V+9GMmlvOKmrt2GsV3PZmFZYpQJ2TkakJavAbGVS0yLX
fvFoM+EKrGZJ70GcOWG3m0Xckkjjha5sAAcZYhh16YVI4y7gd9OP7allrmWmf0Wj
wf6XdMITwyrSoM2sEJ0P30rAGNMim6rUVa8b+Mc+3lQwAxEFPKYTdsgM3bKBD3mP
bvTjiV17BnGVxZ091ZkLR/E7Ir3cWTbw85w95VDAWO+Bd6NiFvoLcGuMrQXYfqrO
sqA+AQWHfccSqP5Ctv1npIzUJVFFDu501YfSf/bR3zDzDxUIqbOwIb86c6LCiTS0
hzczLOtFTj4LYq713GWoqzJt2Jlz3uTLnWcWi8/tkJj1FLUNuktXNqHu1DBgTNNe
zOY94iX3TqjFRpq482ctf6OuhOJqoKxeZxtYy+btoe2mmRHe8SO6/kv9IJsnJqTu
8gJDIA+WZqzbJ2WT8UWaqkZ6/M3EgnIFNjzpa16OkQjtDfGNsp0zl/+l0P8LsgZd
wA4LANvgXYCErgmJPOKFSYbnpw5h6tAE9CVjOkiAXv3O9fd+XsBBKyNG5yUutu6y
FBwCuhrfw3ieByYAeXeKB1N4eMxyhLl5X+niebKtkhDtjmQ50aLY4vR62mRNe9jA
qJ2/PR00j7lxWrHpZBjuexyTaXBqPs0bY90iPKVReWtEh8sEiSqYiuimrDYuoeYF
XKFVuKuIhzyz64nUbtYp0LlphJI7inVC4ShowzzajMWNYf5VHrZgXX8fznpfltX8
WgZHt07XiIxCD8r3XfekpwSb8TM82DHW/BGHe4Ib6anzqnjwOnEWk+suY9K7HSmY
DlwgjUMEPFvjUXMWQYDOnINd98A2p1A6vxD2iQhCzlQFg3JSiIrXVO16o9IGQsMl
W9VTFizvNJeQfzI0OBU0Sx4H77haLLUPia7yiX2+96+YVZVG4fLaIRoT8kthjioN
gni4CZAz16/YAH6djK20mV2tjPY/KTkxDRaUxWNflJZ0Y9+fKzxOtxPeNOxlYtyN
RsG/gAKoalXQcQcmqzhn9Gt/mYCB7RwNTCTmJWgrilQSc+a8G4ewv+tcM/eyb0Co
ZaHTZwkbYKGOI2V2gq3JNpjBErQH6B7yxXG+40i4lX0ttqStnM+hbVDiCPWNU0El
QLnMUhPdf1sIpgJrkkP28KBMdVVyGLUzLF1AVLJTejxpe5couwUVRLVIxw37JzOj
wdc2tx4LLqV4GGCiyWs09RUQU6RQjtVyoH34v2CjDb8xpPPhQntGCNXeO15eYKaQ
veKlwsT0fuXmzreNVWNjdo3VsjDdSF7M2/LH+uWoV297482Mo1DAoO7uKSv8nYXb
7ylLTWt2n/9cpM42aaGpG2vtzZPQYBqUrV+sPM8b5XaOGKlpv2jt9ugbwxv6yz7+
TWN7fzvJYWLBcF/i1CabKn56LVwn1h3pFvl0z4j3H9kSbULl95sW+Qk1Dqr9rxRX
VoVi+9Bnmhv+NkifeojYSfiWjNlBy+x2yMP85KUHX9OdaZ8qU35dTHMxxsUTw430
2s6gYbPNJ4Lbew9Rwef2ntOPP3OeuNhc6fW3ID9oI+P0z/TvtAm0lqmkmErE0GmX
gOZMDQ9Xx5rogUHh9FAEBge4iV1RYkdx6o5sjmlowDPZT+dRikaGNqEtGahVMavU
beLmHd0H5vRjUtsHjS6jOL7LYV62DcIN7+sWukZyZDQ37FcoNVk2uKbAbn0yBif0
m3PrpaBJ6PT/hA7gDAn/5Tv9ERHWXC+lO+s6QmEWtoZPV4p5YBtI5HzTskL/p2yO
3QnbvRPgmGwQe2YRI3yeujyoGFxUV1xEnoJL3NAPW6SSBa5BgMcoX698pzIhgvdb
NAIv8t+4jGTK6iBe2At11+klpEVuF7SdmNkGC0vlG1XHHX/s7IryzcjEGLfvNu07
N37XzOe9OCwQkEvtudpYgaFuIYJZjFROEAla8W0siUzG6+YpM3X6CHIuCdu8Qk+2
zkIE+bEgnMERncWSo299tuzjBMnq5INdUoIbjCrkPKkSjkD643JV6O0vDpxkkdeX
ghKQnQMztg5+99U+awDaT5Okjm/uXcW0tu5QP2TOK1neJ5puAcl7hWXhbMZtwmX0
cpsap8dSgIYjZbcW4LKWnm0t/6OV0Pfjypmfeuo94kh8m3awRfSIVp3/tUNy9Q6+
vjecyD0RSgfxveXR9Fu/WH9X1uGTltVf66Nyzg0LjcR1CmWvDwU+WJHTActbFJqH
TNZisLu4T1tQkycJJKygNJ66mTtoTLMWNIapMjMpY+mPQKAlA89ahsikqsp5NkXc
fhMpesfNQKSSZcdRnuvy3IoY2E5QgOW08e5/XUYO48tKooNNDsMs67bo2XYTTa7E
A01FT53nxR0ZAgov9o4Kr+v380iyWlkoO0YV+MPgkyr/thJGOHkoTKD7gNf5u/Pi
PJSiKYmLkVw0Xc/tvTYd3O9ysmFaQQkXWCUzAIlD+FsTmPdOQHCt24axB3I8YDe8
LACKpdWt1NQWyeVm5XUYJShaSkMbiO39g/P7FK45pdsLZgynhpTftGtXfDYHVlxh
4NkNL1dYdSwzyQOh6urH1ZuNDb7evbkSP+xhkQll5vEOl1snCTteUlo+x1zf+mo2
QOuUCaU+W0TPqwu+fADE/8mhWndKnwM6/kUQzn6Tm9kA3x+HIoXnyXPzO8SxpL2O
2Wla1MA1uxhxqi/mbGdNWoXDNa8qAds1h15dMcUg61/CE0p5xpEeP6WngnBOp2om
AFC42XpzkVj9L2icOo1xQzV1Wh6fbcNTMDDLdTTVcuGv59149KYgee5LQXcPeUGB
KLf8hO8e9yLtQYJpExkYTYr0iGMi3quJt1BDmac5tkgFuh0pBzcIPIr1A3IGQSkR
wSgZ9FAFvfpdC4CuqoaMm7lhlkHTgv1d6riWSiiLx6n+BTYCuvLIHHiuFpc55KDA
m2DyuFMoOdn5Tv6t7thg4X6Z16mt7knpuo0ek1QoL4oPTBExVCGwKlJdb8amS8zD
S/4oUvMziLzjHi4zdEQPfXf3GCtKO4fEBpsdyaOVhvlBBZ9FgbV8Tv1nY172m5MZ
KzSDSY4Y05IbjWCDvP5jP4Ka8WEH1+yQHBBW9ydwheGLW5Ls0K6nqv5sP7WHnD+Q
JaU379cQCnp6yTkdPUuMePwXeTaApmbMg6cGVbgKrIl73DTYN6f+JmPnXq7yPKJg
ewpBuiuB7QcELJD+mK1Dbi7XPoJJXdwPQivEunipSI078MH2s1mtAJ6ZkHwGsrrs
/QhoJFUTm6ktaBQAKzCAmZKpzVTraw5EjW8m6P59yXpfuyseGIayhOGEzA69nJx3
owomvEagxqU7xNYw3djRR2G4Q2MEJRhT84g8jBcW7E76ryO1Pm0ex0z3pOpGwbgw
Ed7QVT5XhhQY/5QmOuKcliA8MpV20dHEll7dLiRmEt39Ss9QeFQ/fjJkm9zAOZ0L
RyIrXjRYk8k8rSXmZHpIrThL+/jN8Zcd99ujF9KSiWYrHWdip+i++nVqDDpgJNmt
QW+clMgi1uEUoYkrRb2mBxZuy/ut+b4R7fofm69/e2ZEGpdsEOks4rYEauJtMqcN
RL0mt54cZ3+ueGg21dWnvk/AdWAFiBIWdspgz+fXepjvvG2pClU1O9lZP2fl2NCA
mRMpA18DTQ3itqP9ga0qoL70CN4WfdzzwdZfBiA5hCIY0OtHIp/KY77S6qQGy9SN
RtPpJNShW8wWxuGj60vQUWJp5TJxnu13Yrv4XB9iYd2XSggsytDuTNiQDURH/hW5
2pIp0yyqOju/jD3FmPVmjciCEcNd+rr8OnMSFPNU/4Ma3UVjKgOft4xv2uDW8Epa
D/gIedFSGbMwzuDuFAFiCjG2VL4wG5SGPLYaOohFyQEHrS+sgYCtYXZqkTACfAPA
YpoaFEdBbrwRuzQ3x2VFqyIX1ZxMyUK8X0Y6s6weOYd/vh+zHMBir9Ev08tNAFRc
AYIkq2py/Pf/w9/tmabl4GJ/cV9Q+5ZU4q2KSwMbnWXbv7Kysi5tzkOhFBQwxDh/
FRndvPi2sYmiVRUbyu5VjEyRElwIN+K2lyLq7AmRp8KGZEjQIJxxGutCBQexTY73
vlX3/b9RPQjpWmBOgjEJSucKw90wL9Oe/2hvzt2kKhhQ2zLJgmd8m/qeD2Gvuwv5
k6b8eO2dA8K5wJ4J/2SC2QIAYwiJLp6o/BGsRGMequn/PjqjSgy1ijqPdx2HLRxc
0XLlQvDXn46lqPoVikDOTnJl3dTLeh9F3atYNwcgH8O6Rwbwy3F2hH3oP40PMc9V
IqLmJ3svpgPqdJ36GYELNIglm+owlYfVthZijsjzXnzTDL7ID7AG+vshWUU8s7bL
dwGhLuBgYkFlX4d3Csxv5ylQvmSL28Q7qywdI5MJwyQHesOOyerPIXbDwAb4zdAz
YIsK/IqpJKxlHRuEWdhumZT/DIGPfHo1bU4rSDtiHHKDFndakZT6RqlGzy/AgzI2
K/WzvTX5gLda7D9BihWgYhnbwhcurIPF270ArxW3+Oyf9YynwACKtty/5mZ4I5LJ
rVD6bgccri/t+PF3QWW/z7gkG3yK6wgNzfAntOEli3w3LbBEy5DP4Ah13SXQ/FKY
PRTJ0bzLi7XRwNsCJpGkRd48eBNcDUyfTkiSwNSm79b070dxu7Fg00INuCjFzBVN
8uc01Ytczh9Zn58QesMRD0pjmJkCdRThpJBiDfCdJGoYPa7Tx80BbEDthRuiK7Vb
aTXmZnXnlDTLrGz+6AjiYtxnAUg0V3hb9fbO3/acnl0BdtyoLoCXcz/Dagw80tk2
wqrzmu1pWUaD4JYOOV9akuHO3dY89sIm4CcjB7rYJgdu6cK4D3pfKWpQ6vjo4ERo
rtkMONbDv2IhnOUzSUWPCn0pI+9RrXD610PH2vBVjlrt+tmXhSiqdspXgJKSVF0L
KSrZJhpgt6tBMY90z3cjGaKlOkzn4wsQkigw/rxf4PQaBd3My+a6O8FVNHKptStG
cP1NRBm4WiicwXI6vtDCyzySjsnu8dRMphVqAu/Zw1iVFVq6/k1mlJyEMw99uNgT
opZxSv/eZ9RhvyGzVs6jhrTtlcFKZc7n94mpLflCC4dTtYv6O2nBb86aL7yUmfYN
`pragma protect end_protected
