`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
g1NjRZ5LWvhGHav6DXGfgPz57Tw1aGtDxHLcoEtGmxJDKHUfKOOHbL0NMx3C20PU
z8M3UyfvY0MotH4tMZ5iBnnMTUF/8nUTsKaAHwkox4mRpg5jtWoblW8WUkf6fOKE
UQXD/5uPFm5yQKKXAiGodPI9kPBWmjarK5qY+JyaLoE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20464)
M6rlg9vtTMU4v+6lKmrVpOzEkYFkpuK2UlnIZcplQ3tn/ohP1sDItRhmNTBNQqF6
MsWhJn6Gc4EGe5Sv9v4qhqmuXEqHNEPIDrsAU8rkNsDf5j0B/gT0Yz2jkpcpVTQU
NTrwdjGPDCV0wHtnh+LkmBWY2PLgN5J0aasiNQ69dO0XhowOYSsgMAL+MJ69DAjk
t4tnu8URJ4PtUauDcZlOFsTNhVIETZtfjgrbUYOfXseG2Miy2CH0kx5w7sgKhati
adv3XlHF5uEnqbAGCWwqXkNjUXHZ+NYEJx6evPnczNJ2TeBXmsk4tfcveZtrlgzd
Xme8Y98KJcGSKHAqnSvbW0rdlj+f7Y3JfYbwVMkTOkk6CRHZlme6kpDrfHN4ggzF
dfPXKPzWRoQc6PJTG+cIMPAEZxP7lAKtywRXvd2vzPhQfqRKNohSyASEs+SbttK3
Up5SCoo9jAwlRIUMPIpWL+1w50ByDAgnNVLbExXdRxSYOof9xMjlVAdkLtafyn54
0Oe7gexazZet/Hp//J2KW5lYM19e4DSNDGKP7nCwvFkXgypAEmSHttW+lvy2MP9E
xXw9ONY1ECxeZsSOvTugWQdUjPAc5RgnN/4hJHbrbX7XwxDBA1I0VjOf6leParxX
YDGc2fwgt1olBu+VD/yfnv7tihSU6sOyXHb5YF0gogyXZAezeIgPUfpbbnbGcDGk
vkw0hbD/QC9U1SYlP9y0VDZaWkeUnJXeQgnSGTQcv9zg5Jv4N3xBjpWXipoOYsBk
m9hclmOTDMF8XatQ8+AjVeSreesdO4DPCq5ju7gJYIhhz4LOgZL8kSe0t4yMUSIr
5g0vOw5+WYUi4G2MAnOKDod+2vLfLP67eBAXF3tQKbAoRCWOuGFj8kqN2RR6emHr
hoQcMBCNk1J29qSvDimT18p/+dDL14Mx9142Tn1fTWny00BtFXn2SzC1SWofUaMJ
RZ7NPA5O05xEC3Fad1KHW1pAWgdmABG0+h1Oe/yO8kEosyQjfWcMFPw0AC05YFGv
Mrpgy5hlfyOaNLhwrRJPKHJok+Lm+tMXu9OuztqjPX7S3dICG8ninHrPiyAWojQn
Juor7NCU8z9pl5x0JoZhxXXeJaLoUKxJLb40DV1wWAG+6aWI7e2z0MvyWHl4q52h
VB6/+oWlBhnHLBRG1gCbYfk6DJDDttBvGPaExenGn2fcNBreY72CMUW8N40/kQ4e
xQVrK6JmqwpAw/wKRgz1j/DAjkkr3Vqn7xBkmy0ZDQhHmgBARpR3hdYBZE9Sokjg
xsHmdNe5EX+z3BANua4YpGhfoMw9Dpp26Aw4XDyIQsuQv+6nOmyrZFWk/38/PRsQ
KUreuOSWHlERA3BYmyC/+j3m4jcV2Ck1nOBzMKeNRGDsX26sV8gfjWBk9dck1afI
og1N3siKHjEIs2+j4IhFoauR4UEjbD/u2twTNcCaYHnvT9pEVusAp95gDjxjH1Ze
DAInO8+lb8rJTkKhqwh4fJqfySET92PlK5naLjs8u2ywoExVrXxbYqNHl3vkQYu0
j7dVSFwqWrIAwodrIO96Hnss9hjiLbvDe5d4WHnyvcHiDz7vXhcifD/lQCslOC0O
KO0P5NJyoi2vJmAtqcqaUNpmqWx5Cx91AYpQBeueStFh/EdMiIoQZEo1jZDe7qTU
gvN53zldust4k2K7cthiuWFpbAAz0APAQAKp9eizdKFEiZd6P76y5GD/qAJWiZNV
Yh36QFUxafElVwvBZzUjwpFq8UTPHjHbGcvlyrBE5dUqZjwCZKe65UBSfFCuFRnX
C9aRzUErFgOwitJV2dzBILsA7FBP2Kcgz0zSMWiUfCnPwYk7k2rmmxYMgKdciJ2b
4xO4hnD1VpTjiXj/sA5lzJSVt4JgSvPO+cRPjccUTTN6/g1XYkXXP9LpSDQnKmoq
kI2ZNo7b2Ik0c26YYGbks9hMTh/FWPrTsArhiEQhow5KbAQ9GRywm4vgrA6yvBmx
5BqiZ+7ZhkDNutF6NxM63uB7r750/Ci8lAuNmfY82Dewh0jVJT5v7AWR6+K2G5gc
Bzx2K60WJccUiKPHEDMe2sB3MXDbls/aJWSN/CsOElLVkmBEg16gF6zFw0LQazyn
tfzPIT/JwmaUrLbanoHBi+pk89TMsaxh2ECatLsXJqDLo+Di4P1+SACuwrXX3L0d
qZF77VaswjHyUVYYYEbxxkVZacv/BrdFSU/AZq/a/7sL61XaRTQingOfATkEoFK4
mDKSdA+yd+AgrkaMeqUHq9sG725nGMdSWrpBDLIqsl7qq3DMZvpBUL4dwC5tcfhQ
N11yWL9v23dPnBHQZNxd38AW2c0hHgObZ1md1y+ZcoHAIjxVcedfxvPXxXhNKBVo
y8cwr4xEZmz5HQa0nzgoHrAbWkUyTHVDXotKvFC0eV8PW2mbYneJeMR8Mya1VLx/
9WC3gfxTbCPiUoKeTnWkqhA/4GLyw/X1CS52gQNIm+CAchd1L4a/zXzmlxdT2Kdq
WWYPNzbdjGrt/o0bhK6xTEfDAd5PseVgdJ8WZGZWQbgcy6d963t/vzAD5x2yVUDf
LYuCgKEQgU6842a9a340VcIm1oWfkXUP7p1P/Wju8JAmx2M2tLFTKRd2Kw05GPpJ
6/xbTe4txczaBqk31QJzc5SpbHmGs2dbxWzZK5dX1a+RIkxsc7aFmdQQz31Anu1D
H7KJVStCTR3zXRTjQkbyiiM9iHE5I0v1aGwos4lWhUxAKDY1RdBUv9dxTQgiM8zv
52DUwCmAV+Ae7mZyrINJieHXUtggh7jVkelE4YKjjMwnds72W1vS8i2aQdlTBBAH
REGsG9eLQgCdgZzrLBuacoA56XUAbyO7DJ+3qL/kE5dP+Q2++vQfdMgxzq0VxsSq
sctqjU8g4MtwztChw9uQs7nBRxp/FXRK+Rhux3+UZmO/HAcDrFdVF7C7iviJo8vK
t2AWl9ytOe4MaoLBWUzHJ/4FJEHbkBH52xWMPsWwdDDMabNtA1HTl8s3fNjpPW3c
h38PLEjjsH59Aqi5hCOJD52tTGCErX6T3mIANKG0BiiWPGFOogepFrAMEjWbPhiu
0hPKl94GXG1L/QxG5fjwQyDytiV1pjj+n0ADaN3B/5H8Bjq6vn0xIeEwfTr3BJJA
HTOTan2Jhu/Ld90D8yksNu0iS09E7mxteK8WqHKF0c0S4Fs/PzPgZTqOC6jJ/nWs
Pb627Fu9XV1caL99MV/8ICYkSz2jhxjhT3R5Q1D3JWR/bpJGq3r4DrQSCNIDjgOT
N5lT2zGsCl3u0nKMqN0ObVWO2v0U7+xetl+dvJahyiRnZsqh5jYC8xf532jC9kYt
Wr5DjiygZZtzR87HB+QygTMcu/SLuvtluF3YHqVRZRaihCb20IIqnZP1fhWSeaLv
9jwaerXOPT7+h8By9Lx3ja77hXzy+6DLQzKwlm9NCX4roLbD7UCwAmCr023eMfkh
xjo7qMV+0d/RS5ueHNqW4xC9FIeobwLDDvtVqT/Z546P3LOx8PZ1sU/B/TpIiifx
LurLut2+n3CyNzooPGeEk/GvhWkA6v6ugKVMfZ/KEsgDKSfFWyIcCuFr7geioZpC
8KF0M6qaO1bd6ymnd1l7iTzNXRJRQJV2VD2zrhcCmTf4LRg0125mQS077TKhsgM1
/EDpvIcYKTG72I5PfRthBIELDUy8qcvmFhDs/7yoK6h/OOhZ9mP8Zuw+VgivkExB
gtSj3UhVn1v83iOCkfkti5adBkc3L+kFZU0ZJuXZWwPWHzH5TMHEaQLjhjG1VIdT
Qe6zAjurKYGWGkWHyS6Qc+zjn/RHtEKA75+PHQB5b4yN9hzf8J62LX2nnjrJCA1B
7OMfugdohFiiT3KaIL/2oOe4/ChHA2+NAACIVFYHHlfeL25wsAFEBcHMsfmzh/PV
zEKBzWR7zVVc0snVxBDg0aO/tfzjEV8aisZ+918IQNHFYOpT0zacJGY7TcqvBTDd
Xb/UXlNdb3FEizo8TQ1o2m1U29L03l0WcDmIs1pHz8VIxAcbkY3dQAhaQUaBSLKL
qudq2C1YGOobkTq/B/73O7NmajorPnTljROzpCxGJ8KQZzO9Yy6eQWVxpG7GhIdm
TpZOVDkC9ImyVWxaE3+kO9FRyDCOn424c2Gfpio2YDM3TKPafFWkzEbJUZ+rexp8
YIzo+qYQ8uDxmHcTHBj5SZwzfsms7OCKq3Egdsccv70qsOK7kP3xXXVvgT9UPSq+
qSpArVY07vZapAVM9I/PInOUNtzhI7OfQU4ogoCCvn5SUqV2gczL/zUpLQo22Ckh
Z4NjjgE9xR9M5sobeHEUgCMnItd1zp+EyPTIflLfs0Hdy/GtAEeeVFzuZxNrDTYZ
9+Nf9Saa5Yn8ZvwaAQRJilPzmLQ6TczWygw2vEVCjK1qkn/muPDJ6TrRVNeJ/1j1
27HaMlzyCWZlO86rKURqPvUvItNcp0eo75LcYxKLnIASZFyr44nePxxSw0BQisIU
jNz8xxDAu3z9Ce1VK3zBsrsKTpcCi+uoSKgq2lF9Sbut0WikjYQ8SYx7vC+jZTiI
QjeTKVuDTGIOuAzcPt+CvdQjKhb2eIcgWQRf7UE4UV5K/nCb2E/36F+umL2ApMyo
J+4A/DhvWM/5JnZzR3sL6O8Db1Xm7/NKQVnxgtf2G6eSSZFgMlu+gZ17I+Of2sq2
2OJ1f2rmuya1WsXHg0s2QBe1JGxFrzG1SsrGEEbAL3nNfvRY7IuTjAA1bVruTLKp
FrUJG//fTCfHLa7A1FwfZgYVezXSLjP16oLmAo19X3vOUhH+UpzJXwlUC8BL8qOY
+FtlJ10VPnXkqCfB7WUQK+dT06ZKcoFfRoVCAmthGhUV9H+VBToWOvbDObVuOuKG
lhGW4V3BWm0DppWDoGvfwFYfDjcTLojpikpjf37r1XB3QJn1DJmQzH/g3BKXeqHC
BmTYBT6Ey1B5Ffu1h4fYFx/vIX1vl4kgQs4t9gMjp8IspeFAxqeMkGjzHX4Zx5sY
rKHFSdR0TuLX318mvfVAMcARp0oKi/GVVjA6QRAzMKfRnpN+ffOj0yX05SBSeE9p
fweRPHtXwASztT69RRWxJ1o008qnJ4r4RwzPFzNeYFG792uJFoONwWZCs1d46npC
9mtvSh30p8q8mFVdeopcFs76Idh2FDa91jczxPzUh0l8RkFN63L9mHOZ6YOMzuf+
RWycmOzGR47oUAILZY1hlK9Mtp49dsd/9g/LW0Hu2Fmv8v0RpcHsYZbzFOHsooDQ
Tk7cTuBE2ZqfoghZtI7cJb4gN0aLCJ4kn7fVd1rh1piBksqwDswWTz0fK1dkDiqX
r8rE/VwMBLSgDgVLHbcX/Y0Ps/Wufs1MRf4DqDrVjMpRbgLh1PCKJboGW+dRPEsm
X/lW/Aw2jl92vHb2LxzBpul3WXJ886epVhKDxQ8lbtDgFP7zk4/rxae1oV5T/H8M
TbOA5KOQMseIDL75+sJq24f88RW4ibMOQB/VPmslc27oK4ysf4aFQuuLZmGck6O+
ylNhNyM4jla3Jl1DO2Ga9m8E4/pX9/RCHNg0XuCSgVsw5EOTO6cgfs/GoiWOcHt3
7OpvTxNzqRl/qQ0Ux/cr7HjD0cWKbuoFyPep/wrMfLJdarGV+ldvAMj4ODxjSdId
rdHtB0ppjFqoi2bWh3T8A5xp0zan/GCyMLiLG9nvUJ1dxdvxMQTMuu3HlJZAXt4A
ud7YNdyZsFYUZ2aQZmdBbBuC/AgzK93eB0zQrUCmn0B/ukkXrzcaTkXJyUgURs9b
JMUJuz0OWBjZY2VWf2MSAE8s1PAGYicP9b/gCbPHniW6md64VPTwIuAScV0WGy7d
0FTa58k83jazIpz6dynR2vB8pyRLliaImlp7t6d8LKS6Ktdr7v6Fy9u86F/5rHoc
TKQuAvh12OCXFRZtn79g6F/ovB8TpLiSlxX/RBM6PqLx8lWkIXcQivOSjf5/oFwf
DVIaBfh+T8lNKeUsXw4VBbUJQ7zGnhfMzIr8Ezf3i6LT0JwOgbKA3LoQIWbkvsTf
sVBtKs6EbbsTgITG51HsSdNlK6jJGlfug0RRLe6CDAtF3ah7VCcUc/S+QMovoxKQ
VIgmE1hYYfjvuApOl7OfNDM3d932DtX+Zlojhn661uX3pWz/+EfBrW7hWyMO/y4V
7t9SvibZ1epItIPbRdy/L4+6N9v9B0G5fwe7SzqWtKRsZnkq1IGFuPe7FxyxjbN1
SkI55Vd/rndn0Vlwp4rdyJshpOQebg+7dI4CZpEW5zO6zrb3102dl059eIJw6jD/
sFXajJIqphvWvC3hQe5mqR2W3WKQjSFHMAzyOnpWVFZ/cLzz5fZLRInarQ6JyQBp
TjMpHRAvFUCcQQIef8w71IPEIx0nYiHchgXyaNlFjytHv9GzfkFuVS8+/3TRd39t
+O1bUp5lQU1E/1y5Dm9WlEpG17gMhziFpOsQ70xjCW6dZ87NxBrZWnnfAdrCWltI
YoJwBgCfWNBYkdn3GD1KXenQZscvPca7XCLC6XdKgNocKrVBdl/2vDkmZXAM9tBc
8nZ4i4tXidOu7ugqUmIl/2vTw0EoDnZzSP1ewNnlgL4UqoEB+jvf1E5Su2UXUvhs
SzwWKBIHx6cyVN9V8Svv3eoNEuH4Ua10YDSuNGF/oBbh9bF/R4DJ5/K5sCqNtayi
p4MeWuKwJSPgvRTLsMHtqezMEKh5otiAcEO2spgFpMgVacmgoTqYtKZZkZFQJpT+
RNzd00D8Nba9kK4rPDDzoPGM9fvifhi9Mumzh2BGZnPhi16Rr7NmKXpEvdJDzJRl
yGMArdKUagW+L5UFqqJXRA5hk0hDH+hy3kyAnmKvucQ1N2CqpFKALKoVUtwN+rxP
e+j3Eb91yNzAM0AjBHLJZ4Z516pF7QgtWX3tw6lZdvaSSumP/29T1qZ9RroWU07m
FxiKQtYRbAC4GthTEYKKrS/kicA6/lCcLG2GI9kiOzMgIs0+q2afpJlqFSuhxEHb
5SXUGW47pttzpOIDdSVyJJP1RYLypQWvdyeAVg4Li/S4FNS8skVOV1ewig6APbx0
OUR2WpUbAKWxH+ayI00VWBTKsvPGUc9l2qb8WsIWEF0q1X+S9fgnGP2g7+fOc6Dj
MivHlD79S1s8D+2PU6VeJmnrC1pPsoO/NMXWGc4vrX1mznYATH6Y4q2/VPk0BfaN
Q65g70hWKO9OTKMPPHADAWhAb70pWsdi0BZC36s0JocrviQn1xYH9XUQoc7+JT37
c3X7GSfAwMdXqTAqwIc9MuvRXQ0Lja9zHl3IV9wQM617On85ObNSX+dC16nnZC2n
QCK99lc4cgrsnri2AgCFICQloW7hG9u3JuD7sesuS9Vu+q3cCsu6Wpk5WXEWazNF
vIiB467mEJGMp+RHtI+2aRuEx5mivFwT6TVlUhUo++Qi45Vcil1/7+EQfaAXROML
ss7fzzs+a8SokWm03Fkr8D1xkGGvFNjhiyCnlTK3SCBHebeYvNMTad/9R7RvGyOC
Kb6K4D/78k/Ljl2VHGLTwlQjsBjCHO7msRUFdHwBsbsZaGW7CKJHAGewsKuuke0y
vcXSHdqBguJrffuJirT1H6mlvgwcsdnPfzVdhqYh3XA/ZXc4+v3rNhh9XPsAusgC
a1ExB9Dj4RhOVs0ojylCxnqnaN7zIqQoV1I4T6Wmi6GP1e5CEwPc50ab6QJxZ+BX
eWZ8z9B3J9Bx2mxMCK4iZTo1lMYbr2SJMp+DO9WMT3qgwOkj05VE+SEI3GmBZU7a
9C00/T20SS1pX6aX65QnDmNrvIsYr5tzULzgYAdZniLRcgNw3W8AZG7MoSU0eVYV
DRMqhs2DTq7r3Sb8EfjEYNYlXCtD6Z5E/UI+3bdHZuaaCGo1aM6VZWJWJfDGekIX
Dtv7AF3aRHDxLwiZPjTFLNpurq0pnOgFkYhiW26TkzSNBB6wtDV96bTim2ZGEF/J
HEwGdHgSYmRz5z96lQOSDiw+8CqRIK7etrK0SvwT/0K0g1mVrIaKoZ00IzYNpbLc
wTx74OmNmvsihpgyv0MgFeGNl+RGHfdJd40cM3hHg9plt7ADsJCntIuGAXmagDev
gCJENJD2NnicKu9qJuEaZLfSg2lruUuQbl34vMdGyBuuY0Ps9dK0JJvtGGCSzPwd
Sa0w6HJtpflaY1XJSpkS8CcmBjtZ7sRWEtZYPYqBaVx6IspEpqZARmu7rouCRncB
Vk4qUPoYzJRYXhF8DzengGVhmrqoVyw8WEfMl9Guc606RJVNNWG/R4n0Y19vc0nl
UI4gGvtHtG4NZyWCjqcJhzYCa3mn0e7p1b17plkkv445y/77kjTClgmQgcC9Qqjg
mIvDN//43EQtb94ZenY5EKop+XIv1kbcvSCddVkqe+IHZio4J7JKZcA6BMm65qf4
VKee7TUH+fkJALQOAAgFxqkIYWOu9CaW/VM69ejAcco1HE1biWa6sIL7eIpHVuG2
nvtP/zPo4EucVSegxI8axQmyIfoH/VA5bGZ5ugPPpi36SuzH9uS5wPsVa9xRzd34
13ct1V9dlPLqlt26qQgMuaFpFYJFAtDcLTbt/Tt0BnK6OFVfuwItaZalVRDhFCj6
juhPIuEakA6TYNuwGBbwsMPoJahGo2xngHFrFP9keZrT1s9R7BNZ6ppLDSaib80B
uOMZswC35xXh3NMdc//2I/VQuLGU714D4L675JNpdFalMRBIg4eDJpHt/2d5ibi9
hgrHObS0ZKYd4o28PQZHSfjVoutT4jwKJ9xlpw0SaecVoVTdu5ac0e21vgv0YwP+
LGE9ie/RT8EqtL7Dtb6g4PwLa02wk42tXe+I9ImFN8s7D33VX1WgA08yRxTUH8zB
iN5Jb5RjdKjEGTam6SZuPtc/P1/3DgYZ3KKhUWbAVtJtFIDBHIYWZmutSGIe/GR+
lZ5j+6UCzZSVZ+5PkMlq8e+YqfJ73LUfG0ok1wwmyVThzsKEeAXNPPIrGWcAh9al
CacO+wTkw+gmg3QaseJB2sD2HphgO3ecGAlWs9r8790FmqZ8phJcNLdL+G1ZChW5
T6YITQSYH5iVX+a6UtFpSCYx+VAxqANPmIFZx5gUMfYp+tt9a/T1JlYgx27QkeQg
1N3SPNVM1BcJY6El/jmb8YHYnGbYSDOBpnzUHixoCtGo4y3NMVIaPl5bTvAXp4sw
nRCE4nL+KgA1VsZhKTw76ozGO4rVUJlyPt/XLsPXagulOZo3HiaJ4A5cnmgGmayA
PRjN5rOSdvG4aL4S7ehxY6/EWrjkDJxlbZJn+SWYR3Krhsj21LRxM5fY+Ukw1GN5
F8PGPqPAylB9LnN1r38hXk0j5iZRyfM2YBg+bKhlQfPijiV5zTP8l3plpzwtrAFK
l3hyhMQesCHLxzEckf1pHsNhSUW9//ftY4MoHyFde4OkzckmeWQ2JWxubHAZF+FC
+WKePeXBNnLP+pc9ECKcBNMdK4tpWjqb/579zviBM1k34c9wZUu+uo5DC/paBwrh
4ubXagpcU7cf/7CEcmZWk+wTER+miENxWwgWL/xrDJYtuzzI1U5PSHDbLx9Tkjnn
9p6K7C8udxQqjwdc7ZjNLvjFa/fezlEjvvPtSmmK/Z8kM8++73if+L0Prg5kJIQk
ahjVrM3MMAFWaZZAo0vPgxJbiCWgu8niHs0tbz/LvTltiIblAAqRCmLg20hFf6Wt
lX6vOK3QwMYoOJ2m3+k48z+fT5Fe0BfKdC4IsTb7mZWlhns+y9Bhv6F1TM+FtVqI
zW7CepvLhjV8/jeDGmTMq5wQUBNCdQKGlPYE/aQKD47q8jLQFmz+ShLLPT2WoJqA
zrl5fYKtjVLoVg7ONijiWM2oL2RLqAUM00TXD55XjdTzH4fYOgQljPr6wpzysrkQ
1mZhfEAXZaLsJHRjPfJ2WdxNXP6TUY6MDeE/XDD+2N1pnyh58od3YKPiEcw9wh1U
p9xE1sT8F8EZJSMg7QGAI1erLe/Bai/CRKNgB/B22Ei8iFNwdihcmV3RxDE8a23J
QXHLiEVAo5496KFTCHzkFAtsrw6qj4vVqGPUd9rDjBOZjbUrkvebt5S9xiPtIgmo
pG2w3WPU01rmPU1i5gxr2/teh6VaejXK4pf6PPbFgDy5r998408XVoMqAVGB5lNW
gospim69scn9FPRYJwME7/TyvFeUHqs1l/LW1P2V6qjh1yaElh/tvYLCi29ZmHMz
bZ91578QX58AuEiMglDSuLjxed7bnvYpUQ1B/IQqeJUwcFA51tV76NRznM/06IVC
GCHsncnUSCgorpH0P7dYKR8a2jBLAe21ufvoOiNz7gE2Idp9QodtnEccnj7PXhuu
ipbpC6MlnM0JgkJgeKJjYI1OGyYxIWalrs8icUVk0randuztmzISYPf0ijXkN3qq
31xEgAfNZ4u4wiSMVopY9K/v0IfDs6ZQqf4w1kD6UZtsY0FxKHynFSpLkzmTV+0h
TiL6JxqhTh7qiB8ZkU7AVAQrOS/eMaSM+weqtS+y22WJtm5r9fLfZ0mObzBSGbdY
UvPmh1zuMbRvdHo7f+uztq/o1i8H1EpNbhmkwO/7AFVn0N66QrJk+/tMfJIwI9C0
ZorymeKwB3w8n+gPu8aaIK4BZ0Dinlx/WAYe/F6omCZKZZQePeN0Ej5f6KOkbkXN
Tk7KPnZg97KwpIwB3ChKJomVfOqlB7mha3prEsC02qldxHSfaCfH0LFczLY9d4mP
I1GZgRnQwbWmqBglSDtww9nXvoTU1f6jM5/bUvH9IVl5UGDhOkem1cCYN0ymS3Lc
5dgPszOay+ZdYmx97nLVL62aZicaLhxmEVNBhGuDUJpKggTTUhx7auu2D+NiVyZm
sSk4DuTPkg5zqenyjdMtfWM1VlpL3fdCZ2wbzPE0y8XTNdFrA8MHv2z55qhiicqx
1LLtowtKpF5FtzrdVJUzWE+dD9dnETOJMzaV95HYbB1rDj8dBS1aTEQIidfrxrsI
p1mQncWK+1dyjdD198iJ+nfuILZBoaHZ+k8MGLR7fWH7WeUEyZ64bvDge7UbqLD4
OHsERS+GYw3JMP/AEKeNl71F+fQqlvL+fjijSyKeSGVUqV6yLUEpm2jJ3mgtmjgG
78bC0kbT62n8d7PjVG6B07y65gYQizcAmNQKI1K3AnOAuH6NVaNjnB1CoEOjZbAs
oGorbLUdO0NWugLgg6oaCldXyvrN3ccifrR1wtfNkBlovXA8l09GVX8SsLVjJnn2
hJ67qXNpTTjjO8prm+8av9WCKCTUiPoEFb0JRs41OYD88FhAeqZ8O0LpBoCrC7zu
/LXMh3SK5+hiC9dO/+7qXvaGmytd7hMNx20FWYMUqxtr0PSxo+lJElcyKe6jdj+Y
tac3h1OgL+Uc7x7ZIfIbV3tv050ht69xlRxmdrYcavL16ORr+5dK5brEao9aX6zD
ZB/v29fvzzXf14tHZzX674JwOSTlksryOdOeZ9m4PNIdXujmCjlDz6p5L9YxJzEq
OnJseZFbYsEu+yXpjx6z7lAvsSSUH+PHNWVKgAGZoa8hRLryfaG5tI1sFardyS8L
Q7DUoblRWz8/TM+ghD02mrMjknUugouuKE1U7mXg1Q/maVrLCjMM9izqsycT2Owa
b7a1PdQc9VW7mIDZBiEoh1qMpbtcF9A2uqa0bJVlpyEa8ilaQZKgRpLH3dhU8hr9
4Sv9PFYWCJfqMhhWZ1cQi5pZZQio3F74AkDrCpxZKv+kOfrgI/C5SyWHZdKVGXaH
+UWiVxtszZ9RU7U8t3oB2GiCIrPoDJ+H9oBO3A68ewv0wYwzUwll521zdA+58wBL
No/bWDBU1l9PVKpLOj+Qbbs888R0zw7VwNcZ4aGPZwM0yYUQMFUSM2d8tAhDZIP+
jL+S94NTj94XvAzewMUN37Dx7IZa+7h8pTVgeEPli6cRvZ7Y48Goq/4TqnPbNHJs
NM04FIOkqqObVfqiV68ak026QGToHdv90/QuA5EYR3www14uesvcjMcSSSEzDLIO
i2FPq4jkp4g2Yx0oUbYN8+ZcF251LiIdnQnmf6uTvml0xHoYkcGuNIThyT8TkLlO
X6OCQGWzY1k85GtYP7ydx9Vm7QHs7L9lEflafzpqmvRGakN4vfI8VEnrR5oaXe6Y
Z0OBBmOowuFqEz1LvHj8kdZONxJccPRlCQwNaKGJpKcN9Uit8Ookn1a669vm1v2u
k7eMEyVr0cJWDohCWdM5/PcPI1ZrtIiaanqEhiH7E0s5A9PG8PmoyGm5fDixtXaz
gPaTLOgycbiqjfsqlA0tjXrc7NEUtf0YTyjA16ujOgytjnyWxnQEFgb65y/IaOje
ZBhU3mCHtcSHJVqARTiSvZt/YLVE0kHGEogU6WPGNT+h3O0rt1RznRcw2/gAkXB7
j8u/Z4ai56Ny4kR2tIGwxnZhf+gtBPg5uYmc4r5U6vB0ESJhFafhNlGzDU1gIpqJ
pNgRYTasJ+P2wx/IgQU48exHLzW5ijjlEv2X5ht5t16T+W/38YQg9h5QniahI2o9
x42LvxJr1pnaYAtrFVwY0LqwCQwQxOyRj2G4+Fnm826DJPk9LtCI2jrOPMW+/SQ0
ik1d/jEp5j/+HI3l4XEARbR+gJxE7Ztr4UtefNXua1uUgPdTf7oVaNMdf7Gh0rEU
QIlodCC7QHkoivqM3A4M0HtMGCvJXV3MxwdcGNoHDZPoXfurvaJLmWD1MeG6af63
FAoY76HDuS2smumwwO6KQyubCOqupHlmNWBhyARwho6Sy7oSxQ64gjpbNrOR7VuP
RyhAnT7tUtWX6tjsHfSJ3A+t+o42i1bYiuO7CkMj23jdEbWHFC2tmEKPMEcJmWXp
6UB8N2BJNTQGrCbBd7xIxPv8me5LXJUiDhulIbheO8smagVSRJsSNZcl4sMZM61a
NVQceC2mVfcPwgIEaHhuPOjZtC6a/b0NtdKuy8s8MlzW0poqM+jqdyFHzR22gfOS
wwZlBqJQxXAZwOHyRCO39QOEwOJ7nOhuIUEDo+L8LMjbg019F3vLYC0m2Gem+Lcc
qh2BVeOpC0ct6DUY2Q+FtdxBbU/4Aj+nud+Y3WVr8sMfNADIoceAvImcMwc1rqJb
Zn24qW4mRbm4t4ffg96tsTkqUYPHsbO1ddgrSXGYShjf3mq/+/GTm6Gw7M1WDyX3
fv8jsENJYxezAx4loD0V7RefaZGHAHZjroqCooEhVFSW6zIZvWq5vdKdyAxVr+7P
DsGWwcYbsXmvzzD6OaMiFHEAN/LBVDOLhk5oNcJ+ZLMwTi2RUAvYnJGeVY4Mfaw0
lVc5FnA6ODFXiW7FdqDN18Wv3z39aeEM2czMPJ9Dkv241E77m8GSN1mySZO5IrYS
hFWF0KMN8Xsy1O5sXqFZd7ey/KTb1doLJVoEnUrrghIwCv1mWTzTzKCMHVz5WFKz
yRP8kxanma20yhU7cJ4OQlZqsIisWUI+alyQ+bBSoe9L0/XUt10rmF5bVBBfMfgG
LIykD6dr3p0frgi886EWoyCoS7Wx02Ic7aaNcN6CoMf8SL97gjXwH9XMkNWYesgd
X6YbHF+Bb4oMAoLWkHGgQNiVHpRuCBC9zjXyW7+uBiwxzbKBRweX1Eu/d0xzkHp3
eSwwsA08O8ve2ZD7LDPGQc4YSpAOptKyqEdTmO66T8k5B90xxLSM56UkUdIR9cqO
wpRIWfu3KqhBVNSWg8FoV8cRSrrP/evD9hswxRzyJmA1GeIVO13yc4CV/0hRLYYb
24xvcccycs025Q99JONjbROgHoGflchRhlNaYjOPJ27zIAtBX8s13GJZNelVbuKp
2Ghnk0sjHRsFRmErg/ISo9mBjBnyxhznzn2qxQxr0PZkMUM0rDKmKXgGJ2rTZzXk
GH/GOX4xLIcDLEcT/vV7Dm7PV1C1pcQDe+JjVFQrAwJtA3q4uRHT95jVC3CxI+8C
UWMcJBIr1IuosxjRoWfHXkDm13oL1JFWlFG5AWpq4egRyV2rXeEQOqP0YfwS11v5
xRwXVo8prli1NoMzgcRPISB215t8D0N3930pUeLj0GBsXNWSBP4J0XW00Dlj58dc
1PWAQdxflLnwQRzAOwqVrtVPCnSbf+5FSCIpcRNythV1fsiQG3MoFd8OieZwWvw8
AvRgY4IIC4xhEHZAtLG6SYlF6QUb7ipElMKJW2F6ZOxFDOwVzPxlXZRzH4jTBZ3s
HmKGhFpOnwuNo3Q8d0jTFe1N2smBX0UWQ/yVhTl78Et9q/uLvHp4/tluc2IFoAbK
uGSEoWfcwsrIOdiaH7VXH7nav4NzdklSJnsJyctk0JJB/TD4rAKyvzWREX3Rp4vJ
GYBWMF8ygLr4z8jPakshM734Lqd8UN3MgKEEYneLNRwIlESHEPVZ2IjU73UPreME
yPCna2owBLaHlvWRrAWgYlDciyqXjMlhYw0ypSMNp8WeKRbro8DMty+cRpcqGcri
R2O0FJC1kfmDj4eo8EoCabr/JhDVarBsJicLGwyJhPW6dp+uXSuMyE6UTIvQrHhf
bHm2XhRmXmBIyv1DA0WBb6NVvDJvR0OTpHsZpUkR3hltyskLRzOY3ea0eHxZTIGC
dGr7AwPXLE6XSDss7XTFeSczdTybCgNmQkVn225inSkFUFR9B19744oWP4MPI28h
dVTDL1BUcgfY+DtkDjKqE32CTf71iUDsbihc+xZViE1mu/yaaBbWLcX++i7bg3YE
FYasnKprQmO4B8kJ9Xr3YeGaUDWrPPReuXaTTu4J+JZmOWtMZ/m2MMyqmtSjUdnO
uuJemhmIYxNnemJv9bTvsc3J3l6Qdspr+zUE1kZRNVdznyUdk4TJfSE4jq9clm08
q8qRHJtzB9YwUsVfsFsD64oeNSwLPlHwdegBZz7hNhG5wtE7Ith/Dv7wdFATSgSp
jwzSAnk4IuRg6twPoPVn4kBlPrF6a1fZ5f8LtGJ0k3zfmZPqmA9ZnS7AYFwbWHm+
1LUkzY63/k1g8tD9SRPMUlDojFhW3vx8copL+rYklK0qqAhoTQlHA0rr4q0MpO9k
q8ynIpzWYBcBEb2p8UxHlZNmMLjlk9WjNpNSfupv3ELM8q/jzvBXTmf8uv4lW/A9
JRusHLAbGP8Rf8eyv9pvK3FceTBCcwzYIiAH6TZBFNsesWcPa4kiXBo4EOuqVNa4
1qCnVQvpRE6dEu5RyYGb045J6W1dMZDcbtSV1fJ2sYTr1CKBTb4t6VKVU69dTT1V
5H5zpyU4DaHkBfSqpludAiCC51g0VWmSsAQaHiVIIWq3mw/qTSFjSl6khnXXAXHF
UYAobHE87yFbwUJwCR7XuzlScHCaDVOqTG9YmxHAcSb8LddpylM8MjrGOwswmyoC
Qi6n39SM7yaOv0ytUuYmsJnDeljLarQvWuanrQgXzY9yoBnUo1TY/fjRmLT3YiwK
p3pxZ/QzC5ZrxI8qJ8B+CT74NGJlgowubdr0CKhevtN9rZdcZ4K9U0d8X0YIkcPl
V2WV4gttKRUaa5mazWqY7AX0IEoXfvGztJhLomIxO+6Ygc44G/QE8EEboYpf4lNM
4b4X5ijSZ6aeq/pXVLKRWt4182a9xcg2ZFOaEjjHRPgKvYXdfkKCeVZDP3Ah6H4n
PCeK5xrgU6c6ShcVU+/Pahi0QIhYCQscquXBoJWvtBs5PGiN2chkKNoHddDEx7sq
xx+/s8E9x7LP9jU4s3RF1d8DFFaF/IkPj+VHPVWxMuKiKnJJo3LnUXbpNVcLgXKf
dn7F3bU6XeHEvDqefxoQAw4/PhMEQKZllF7GKLJ7iK5WnDlxpNpGqHu7G8EzQFBM
9up57S8Ogm4kboOkeqDT+M+PbRfdoN3anFvNzykaDu9lv87Xco0VPhJFyeHrMU6L
xoK77QORCZ6MxHesy8PxoEzYckyd9ozVzmp6xo+Kf4X14obqHT5nmG8+8pK2UYqe
1Qz4e6U+fhaXs3Y3jWk8qKv2j2EhszQQAiXQ0N1/rR79JldqLy4eP8Il+ruvqghU
mMP8iVoUHw5OGd/9ClcCNvT5O8FbVhiFidk3mLl3FUrwPV3dM4MpBQQq4q+X1Doq
MeW/oJri8c86ksV+3I3VrllkEOdkYSQfalHYDdxAb0kE4RkR9HFaeOSTAPioqFTt
7x3R6P4NDlr7mlbVLPFe3OoKZsD5ClfmotBsZLYpOCMylU44ig31efEX7JKXfzBk
FU8Sj2x7yjXLZF4j9ZCMKRZGZvp/HCDvko6BbYq2erGFumPJk1vjYuO3PPK8TIuj
LLeYei2k3t17Fd3iexuoApxTd6p66IMMllzc16h2t6sx1Z3u+awYWC6VH3Rf34QK
0MieYezGo0axDAIdCPeB13IyubecBkchrG+8Erlci2DGo2cznsGVmX1AKVpcq+yX
pja92AhpvGm3vaYaRuHBeTd3dT28x7yxdM3wjzMArajHO/4+QbOkmoYleDR8YSxV
kF6TAufA0mWd5DhktvQMKeW/QWv/atQ6lV6KdX8uj0wjmZ+w5my2wm682frxko0G
963BWx0MEjBnN1S3UuCRDUMTsYLE1DZJ67d9EUX1YqY8wdtTiRoMX5BmEc1Bw9KH
PWbNoWwpVKhRjHS9Mh3Fz8YQrlUewsmVNGCh3u5W78dTa4hW/FB9U3nfs0bWSqOm
kUG5aGiQSFo4Zf5cGGCxCUL5yEByPaiucVQFqt87pwC0xfFwQfFJNsor3yzjoQBK
Z2wSrs0Mk8k93Y8oQz6x3tbj7HfBUKhQ+ve54h2HzFzSk0DTyawecmphNPrnJa2d
YYM45HFXaBxEvVOEf5SZyYeLJoaDDM/nJ90mfbsSIGLQtQjcu/UPiHsdcJEAydHF
LGa2+4q9YYXCcCr2HNaOyPrY2V/BnF7bJF38Reh4wowebyeurwRwcQyWxMmW34B3
/SLnK1slSIgV4UA56olyosCNuP/iUh+z0r6S2i4NloLDNapK/Vs/809HClOja+Rp
TeVhU2W2d1jmnPVpqMJDkCojb+9fkF5hXxCT80BtVpyh5+FcHGXihhMXGQFfSzcH
a5hVKHdYRaxs0huNcl4/vRWvZVQU3Jit+Zd5qAcXQmMccJSiZ539lAJeu3WAXdMY
khSm8BHxDICAvP+2slqEqeOqgRwI35jVmWCizW7xjJdUEkpqbZdjPXYuJdLVEBFD
yx1i7bDUmL4Y4TzK0BM3jLgKaDQmmx67jhr7KPLlotFH/ybVMd3EhD9owrzXNg8u
iyCP1jc0N6a5J0X0NfK/VcmjgV9g3zE3INq/zaPJVTLBYU4V1tngDlWJobevAvYT
u1ItMLVoycRRJDbiAFZdfYgNsuN29SsQ4oDryIfpYur3/DTJ9JwFSJeEPIKRlAP1
IuCtSwpEuuJhchesalNRtb7g4h1SXhVGFjZ6cLzm8n7xSaLNoFohUQgzPAoPLwbz
yBs64Aq/FFd8OCmMUMOi9Fy+odvxHybMQ0KNVvgmL+EjzDYUmQV56JYYCMuiTADs
+MSo/Grb+sMEvNB6ZRmOINGXoWKdgUJr/PXEiQgM0Y7zxsS4erNO5iStqFzPwJFf
mBY5I78DIK4vCTmCIuH0GoRzzaaQEbvUK950QT6+orw9tiPs16qJECKoX3HCRP1R
C0tTcdpM3mRnz25nyxEkVQ7DR4pIavK9Vtg4QqcWm7i0ivYZZRX+vGR1Qc7s5/wZ
gKQZFAW4uQ2sOJ9PoJMKOALhsCGOp/9Q2FyEA/aQ4C+WenXhvgkZTzg4vPgToz6t
bmlQWLCxjMJTLXieG7Ucw2CQDkTG1WfDdu0NtW8jXdrDnwhMsnwwFpJR2Qs8zAio
L6zfOO50VSm47VBE3qOITPBHkIDGL6COodS8c3QEbcYl63lk848KJGZEotGR0eNy
8Daehnt5GdFdXWZNnqpOYYCaAJrDV4owXVS9fWGIWDQ9zr1Ynx2gtFJ4F65m/4dZ
oCPKDBcrvlJms1/lS5v+GT2l2qrcXciQgmC69R1dC5Ys9X2SlNPVW70r99Nu7Ky8
6jXt/sbnLL6AuKD+lGT0PhK5KO+xlu0ifWXDkhBgTi7AOLL62pZIAN6WmaYr7lF2
/SH9NhCqhYjyNYdjCbLyvirZnmjuD0H482uHcf6BMZKwMSbBFIZmgrv8mh7ZZ2a7
BlUzEweXDegOR8VujVZv5p6VV18OLdo6Y7b1qD+EswIJ58ZQWaFjGfalfM/975ql
sOf5EtJyxZKkFUwQei4oNf4XrlXJiiCjkvs2aJVdLblRwESxlDcBzdncnRz1Ybdl
pj6gsFtRbQLznzifzOy5EcuR98BmHbVpbPjd+fKcl9kqZo80gJ6iNsRrMhhggNWE
rSYWXLn5SuR6zV1UBBERXZnW8ILns1c/o9PaVEyJ4y6/rWQ6slav3cGV1lu50hfd
J7DyHl+BUAUm/IMSbc/gp3ETFnTsgaErRev4gnJ/h0tXF/b0MRyuotP+Ip0wqW07
EHR9j0YgmTwikxdEhVJ2MpEm3rhZgEV4BG6mbe0vnypz7+AHc7Uu1sOW8BYov6S7
5/GI97++vtfGW41sD7iim+CL4jaZvAxmbm+H1tXDSCIg/7UGO+okQNHN9SnOdpua
8KjJ56hbhN6ZxyTksNvWa0QpoplnCiZ5ccZbelO4iSpePd8Fw1ZBZ5X/+eYJQ1jG
lFv9UyZzPO7inMrf7Hknj4gglSBHp+w+CVoQYNP1qLpDr6vK2vdAlwHeK95Rd/Bc
2DbtlWP4TfLoPpBTdvxuiOUjK+Vdeo3+kQaPFIaIBGKQ4seXAOaWt8uSgJRqOlbo
LEfhg1KOkmLpMql6fE5Uog3ZDjMzUzhxyGN0fC1D35GJbHWEpnjnbJ0qblQ5vaEp
3MaT0oElw9BTwhdglGKRo2elEI5nsjAHMQsJS1B1gbKTE/Cy2cmOANCo6hk7B6Cy
YKesOMIUzbJnfF2doZzx86R5UeCbrUg5WFRNfpRYG7n09wxsYxwhZ9TUa/p+Ngl+
FEP2Zh4dgBxfVElmSLikTOqe7KckI5JRxTcCfW64OvtX7VblpYqYNMr6SqOuFTA+
6Kjsl1dsZY/Nq0os2OPIuh6xadeKVAc7WMoFA9sUeZsKeBg7h7k+DE82pIPUbp1B
38lZX2h/8HC0TLj8pFFZ8t1cLfMtRpBJZgqauHWNO1bD9ErX5Sju2dXC0wt1XdHW
I9+mB7jWskwBGaR44S32Yb8/VvQVCWpxc3QrmuWaeZQXvFjL6h1jX8fuOizsVapE
xW52ktajip+kcJfpn4gWTmorVXyd5Ja+ReSo/hoFg+IBut4TJbJrqyPhqC4991CC
DBkKNLUONVwJnh290T/rS4YVNXXHhyKb9WthRdL+nZMjJC781Ir988YrGLBLjIa5
0nqsZtNAOhNU6r6GKzDNN8gUDndrC9frfs0Gvq1MSTCkmM7WNRD8DN5N0KF+OMpi
Oij1mHypgXLektEG8oqsfSPzU4HYvp6352sns2FlzOctgvC4oo7shmD25lwXAidu
ssx6bmv2oh7an4NaaAcLb8fnUA57hUWdtb/OZy19/PjCDi25Dif1Llm9Y4sCQ2ss
Sr3Oj4+Nw3UKnF6dEmWopKGnskq+szjiboPzq1I2/Fd0fXRIWg1/I3tyD25n42v+
k/1QfxKtfIgbikf3FJl50+RylP/BBD1ahVHQ5skFZMgUwVqvXfGzqXiqWNewwVig
es0K4I6vOV2/IW78qk77FB/pyhgkl2aLbcKTzGWk92L41zIIwf8tTEnHitso/cY/
urTwO5J5UkEKZUCvuNTMwz2NfJ2bN428DLIBLktlOe3m+HbFPZogI2sw2Vf5vyqt
HMz6SKIyBR12HEFGZ1565SX7twXhZsO8tSpfheQF8DHoa+TbgF3jK4nAh3ly2Aih
BxDo8xAHohcIoAqt1wtOXZ0Zc6dTTA5AY1dEC1nmmgBWG+HBLLhu18joz6kFt8mP
UJ9clgy8ArRvflimXO30WRQY6uogwogHrCiSBn6E4lfbM2YKDGnEaeRQYjFtMQGv
AG4fwJZg2opKkzQuFSs31awrKxSI5NArv8uB7EthVK0WXNT/DGWaVuCkDpRVhGKo
ZmBy1LqY1FjQouhUmeU4fxPuNVZCRbOY0LpwtR+lephjhDHrkWJGFwGefVy4XtUM
wuRunak7ScgyOt8WScLUYwjLyqlzf/HYTVkn4RxQVcqY9qnj4rj81QhV1Z3uoz5+
oGbR3Ydc1WpBniv0Tz2cdtqzs+kX/9wmWqgb78gNemVM7ne87kw1I3wbBEn5ssxX
h+ivufp0APB7cxmCMjXsGr47aGUlndXY41LGbl5biT7pKHHULSUpcFaI9AkAu1yv
QD5srws90MovFji3sss+TjiLoHmprzRo5cCEH5hj07YjQphhO/+cEz7XJ4s1HEDa
AH+QF7sD9EXgypeWqE9amGFp+D0xcHNv4M3IE+J4PqI/SgR2Dn23c1KOVu+HxcC1
y7YLXZRotYw/xhGHvXARMKjCx507ibdi25yXbBSOSBfgbKREDoic3zbblraOhUuY
oi/8VN0qpEZOZ0CMAzBHKDd0fzfrO/j0VXkfiAZifN1jCr4BQFDFiIxmfgO+HP5p
tYTEazDMsW167p0e6t1PkL9+vP+rcDqAFBuuCCd4TyH6x5wL8gnzvbZ+UE3h2mya
EWbObBzBx3DzaaiLEMipfaLi4ATzyE5Tvr5O9eqATIom6p7+qy+C1h+lp5CH4Yuf
xiTvPxh+L7WxU0uWLZb8ibotBgE+oABOtRdVEn3G9lSYDNdqaMJKIRYNMWhJQTXg
4b/c/It+Dly+G7fT6WlBB54dsKFbLxamd1s6gPkjEF2WcKEZZt0rhrczx+mpiK2b
YrA8LdkNAfjMP4G4imzYGHk7k/QqZlxVDa458e3c8ampxKMlC2WPuPPFnC9ryvbs
W1CS3Ei2spcNTVi64B2DhCVgjxwBv9aVT72HF9+2pfhHHtfmjpYbkmgk5l2yFU0E
J7PA9pcXpsSPHoDFFGZ+xUH/ElSOClJqdtq006x/JZu4/8OQwIHbtv6XvCRsCqLt
0oj5apcZCA9NElGJzGEaJG65xyjthRWi28ewm9jxzeyMCTu5egzVtp9RjyxoPnrx
SNCG1xUVbvQwLcAplzn/j5zXjOW6PAfEUuIgqLjx4Z4Stvg6KBskPWeIOZv03ZmK
P/rWF6gTAIVS/CoIcEEoLVcL4nSStainBR9EG5hAAl4a5Efc6Yy/g+Ij+aCQ/xFv
Dy2nNRtkkRDWbNu6+J7yxCQ0RD2f7RRE6wVt6OqngZjr8vQRGKMt5FIzf59g9VNZ
WNjFK52n4QpVrZtp8Y7acnVepzf4/cDNmpr7zR7Wog/5vG1DUm94s26ROnHlGQRD
JJ40+6QNM9T72d9Fr4dkxSo0GK101FKJ2XVIkmLOamWgDQJdf35JL+jrJcGJla5S
Idp0dRqqMVvCVjcwqdapVt2RzzRW4OUO1GtMolNdvbrdmyQKzILwTO2lDNTuhhfV
CKp+mpch4MhVtD/R8uPNvkw0AwLLP7ayxbimQ68UjJW0xA2u0BnrY+ndJHAVC6xB
LNSirJ5FqeBUchWiGLkbJ45tG+avYUtPCQUNOySMy40OiYquPKO8sQAok4az+hIT
Gi6xTT2+h/yIXLTT6WCpfT2qk7vHDh91aymBjFfA+hjMBdUHSERWasrI5PHjfYTW
bqs2l7Y/kU93vq4Rkft3W8F2Z1dKxVGxWU3atlUSMjI/YvEM5Aky1KNSnUor/mQG
Q+LXoBLCBSoJVP27kYPZA31CupuFUaOKbv1kKrSKa2jt4k1MWzqlhLUPmIu6Q8+Y
ypOO3+0t3BEAhPDZ1TEEEeuWfmjH/tHCRx/dSsHkVt6ymzFwSwiJj3jS2K2g3gw7
k6hrZWRnJkh3rpu8tMbI569eTE5Rt4LpketyGYtWY8DTcLRM2srIW4BWOxPplhys
Zvf3DxdqCd3mcYyiUST2UCbR3ZFawlPNkP1D/1Srpmqwhykx1VV8tvRWFgE0NHzP
xq5gVn8XHerrhjkUU7CSbwZcFH5HxyDgxQcO9O/+j6Gup7UShV2bLDZNyed+POOv
xm7zbz16Rlri571aDquG9SlQ9jm86aw0D0xnqoWLL2n8fEyrjUYKXumKL6RiUccT
wE3bFowTd2MRFPkuaqsN5OOnfjOGuK1KcCojyHzyrNJ99da4CsCKXNkgJeqq6xWP
7vdahGH9kxft0YduhPhA1Uvo6kZQyzxi/Rn4X1JBxo1ltcWfYkYE3IdP7VIF96Q7
BnD5zpEFax/qlUtQMWZpEaC4h+NnoYocTovwCBwadixwkc12Y98cm84BWfg73gIp
hyAAM4/SePUmLfvDHw7STsc7k6rXdc+Vo2mN12gKOkVeXxZTFBmpLxcDtEfjGX+w
pMQycZg9z4UoQvBydnHzXuHORo4pLbwi6CdhGcn6jNPZrBptDxLBcyaQC5fFPDwI
Spoh0Dg1ZkM9/+W5t2F9HODAX7q81CMkbFy4CrpwJbXnTGHEw1cy+WsZFv4PjrKi
az2152poEOh9o3E4LEAP8Bga74M0Ec/k9onjW4mrsSZvCUNBcxBY/r3iRPQ4ZzPl
VkXBT/HJwako6W0kP04ROX9NwQTIVlqit3RF5hx+0ot9rpalJeqL90KFGgWeQjTf
iS0XMWh/rYWTazctokTyoH/nRE3+HQwP8pelzGIP8yM7vbAtN1UKVCdc86M7t6Zp
jST1tulZ/WlVZr9M/P2MdUWyjZodVo7ycvAkQl8dh2JFdlVY1WPdTX/fi4P8QmZo
b+mCM2v541aaPiE+6UGQ6bPjjN85yGhSCpzKJ1VFt98QCxJD0qf2sxUJhraPmQGN
Ap7v0nfEcc3flSP4hyoB6yaq/sK0/NXWjJxQoTPbCrPmra1c88yOJn10/tZ7Jl8l
kGCOBV9xuW/dO8/ctKc/64MhlYo7mcFbXutT9BgJTbO364hkcL+DqnUr9cKKvAKA
grm4HKhXCnbTsKJBcbV4ls6AWEE9oWJFUvhJ023ZpqBZ4EJjyixXsin/O0QVZXfD
YxtOjgbde8Z+2EaepsY9iIfw+uOIO2u/l/8vb3TkxItQviZOY+06H3LWVLaN2M6B
EhpWb1AQXm0FxZ1UZnRnWbcgKreGr3Gxc9i9fIvA8U7gjqqGEUe1YDq6vb2Rk06R
3aQteXqqlvew+Xj2QQglLQL1ckKVlafLks5eaDMLZZXSotCPpljV6jiH1k16PzBj
0kzqPGVPkJlRz46fP+5VhhwPJ1CFTpYuGzgjkFWfyWEMjmoE0YC/IKWndVF3cE1i
wJ7tN1nFClA5n7QyGzp6j4nkpKmbfFkJ8hkONlYIaatqfW7xaLEcgx1kVBsJQOlW
iXyeGZcFwarE++XYRnrTe3+UlXkj18l9WlSzOlbxBu5jgwvaRmPRbFNhcxfa2VMz
Am5jK7m8IcNYN+/da4w7ZYDsXk0T8f4Q5q8PItnNUxDoSes8YSDk/dE5bVD5tea8
vJCIDdPIQ5fvRUe5V0pBIH3E3lMS5EaTv65+7QYrO0V/7WGce6feX7aHdudiLXEU
N7vrOBgv0/jcL4NtX6mbaKW029tqwITyYAgCV+y5/O6ppp8q/md6sNSmoabDq7DX
IwiW+8+SdagV/lwUSObOjiZPBei3jQUJt7fVQa9kK2hWIoQlSoPMkd7eTCc8swge
csG+4tZEqSiVgMQe/79YevpzkjARzFB7wiJkon9dwDOCwi050NYUwZdlf6Ajh09O
p7ClX0n2S6D7l+mCqdM67ANAK4v8bxmjwwe+7sOle6n1XLbv6tC5RXHteowbGI39
7q74vsrrUEZwlOWrNS2x+S7RbRZlA+7yUjWdB1qnwKmgjt1yNcwa0zLF5nP/bjH+
vxuRbKPIFoawXLRsfI24n7R4baDWrl6PiKksRy56UVhu2p3/WZE8U6QH8g21PVXn
FDrvrwdeOtM5fYbiaEw61WnjtQ9AV5ugaXYVW7S675kORi5LRUljP403rpzlB6ce
qlKaXutp/zhTPWui6qLKwH/xKAWlp3yr3SwrRszgT/biTzN22iHXOuDm5H2AdGnU
BMvDt4pAkDmUbwO+fHgsvabqiCVz8DdXtocFnuFTGIrR8Sz63qTJAudI20R9h6vy
5gqL3K4qQldy8aWydDxY5DUgvA9qkdz0HrjLdjxpFljkahMIrLAZRfKkF9kWHh17
3RRTC1xWKrwOfTQ7Nabnzw0XbgG+hT/P29vYpmuTW3vTjbUsYOlw6XwqiNQn/MVm
yCn89n6l8U4gGoF2qBfr1gXoXRbxOdHGIGLiicyjamcgszjRCQcuYXflcs36urFN
FDrWqUF35djip2cL0p78eH5TVtnMjg85gvafGTrxrIVyguleMWyewC9uIi5n8GAL
na6viMzUB+Vqy1iyNChX2aj6DeOayRhM7MMAAf3/rRhMXU5lLIsUS9MRKvieN8Qf
r0kr0hKPAGQbw5L2qCx5YFeffu/0NmV0onlqt+w3lpqbw9cQAbfhdyp/BuPu+O/k
c1oaxyzCsQx5ZHCb1rOsAwG06TMSVTJUjwNmKkIa4dAoKZXY7vjcUGKvRgPbmQbi
IMWnlOZjuALaPUO6/Q0TZvyklVcfFot2xbA/iEFNRRvLc+QijgqVAgGjlC4rf6Ne
ThFdOU2wtb5Ur2tdoD37PCwDL26MNQH+0OfcQ9TzRm8Jfx76KemIVNedfn+bCgFA
0Pl/G4XSYMJt60Tmjmn8EV+pfUQo0NFRXI2054VDjPnoqMnvaogYBBAvxFh33UN0
ONg9y/iN/Zod3esSXyBWbU4TjRJN7mxW1aE/1bv03h4qvFY6+z7O80rS5eNNVnbd
bJocCPvUJjN7QH/Y27oja+oHvgQIvdxDtsTJKyS0c4QU5CIeScyg16qmFvZh9Yj3
kx07ab9jSVLXwKSLRzgZUX+lXI6d0yE4AbYf8YPOKTEJdw2/8HUwt4yNpXDFTsoY
4kfehw7/q5wRJsRGqyIwd+0LU+3g+wULuavkT8qwLOkriJxaPRq3K0vBdE0PQAwM
2mNfS0UULP4Hduns9DOXVSflHRcRxh0mRhbn0BRO+pGp+gLE9Jw9Fa7aSUaYZdvx
xLQ91VtV+iz5PH6p8l6d6ZI/p3CjHaTS6NDEc/Ikj8hyE7Rc5obBzbG8dvtLXpya
5AGlRBKO8Bk2N7WdDgCAKyaCHuT6k9T5wbMIesSBqHG99WWnN99UZb+ugw1D33Cu
xjnsdXjWVbgEWaiOpo4FPSyBqjPv31ORwxO+ajInEW8nkOWB0yeSvtErDnX32qgc
Z62YqjHs5gUBBBJaXxhhnFSbg8kAUnOUi6bAfGKU3v5NCL2Jd34scxlPcnEWDi4C
J06oU/budvGDqrxkcecF2D4vKwLP31stpNjtS2KDAEtH/Khih6s8vP3sEG9h8+Bj
YKEMvY+VwuFsP31TIw2YE62R0T0ua9NKQ0sITInO4FGVjogJ+yqGzEz6z4r3D/8J
1c+j4I+bAANAn8tL74jHnQDKZ5HUOsvdJM0l0x2vjsCNzAxgqaIYSnIdbj0SWfsS
wrP51dr7pExDFrFyKDTPznfNtVL3eF8lhOT7O/mfhiPucPHZuyiZoV4HroRe4M9q
QlpyK/i2MGg+uHT8LJghRw+sTImr9bIlLogMvpzbQXluDZgUP2+rq+AJI8hMJkL9
v+l4TZs1JEs1oZCpnghC4kK+mCXjMYtqs38RoSWumjmXgJrD4/nWqPCb/zTPwfmd
DdZIyl7kuWs8a4V/1zHPin9cwvC/IvU2bhGXTw0sQy6Bc/L7uMCfwRiriFvt1okC
WqiLlZHMgFB+IweuxTPSX26FbxrBFT3tb3npI3rdjbsocRzlpsE3HmTSRFs0Egvh
LzV/SMGsn6qHE6A7yFQq1cxyDXvJzXTNvVMQcXpIvL59uqZkOkRFrf9MXYFAO/UC
ZB645rg8CpV6NkEfN0jzbfo5st821YTf70pvWbJUKWqoCebDDpnnNdYrRvOPOcZo
sffU8QIVwyZyfs6pS4UTzYnuCkEryssDwos31jYxuesly+KzL7U6AGElJe4bLff5
wX98UfFaqeo8kqZFcO9oq9Ah+jKmLRstTatnojvnVg9Cn3TzrrWnUGY+pbNrRiGg
K5I9EY6hZB+MXwdCLIAdjnH7fqnB7AbVvvAeKnV9buJcK6BaPjqAMIstsFRCWlaU
LKmk5GvC7RDimYE6iTqTuTP/kSGT+2TEUDh45FeCNXDgyZnxVfvrHAb2zBjJenA3
0W2anFSHocQ+LTIJR7ZGNQrp5+puerjT60Sh/4/c+00TSOI3xqAHtk582MpFF7G7
kt6puekH9WGJUXW+ZpKy46OZtMNfac2NI6LJCRYkGsVtTFhXCh2Y47TNW8gSCP1V
mEk1PkBOUvWt77E0z6DAY3iv/2W4EcURUXLwJwHuBkDLJDM2bM4ls/4aaJ03Vn2R
dfJRrn9hSSrvKHHmNX+ODDE69vN0mHS/jxhcO1Oo/Cny9wmrQnp4cLmF79pFM9a1
N+fSsACHbAkhwEqhX1oYMsLSDEsEeaNBQ6XDetgW8EYsVtGj8fim/D2ZdwEHmdEq
xv2Ee6fQ3iqrCyvXWWBdv9goLDIRby6YS/ZK3XlHDTqSPSSC1BSIQR0XVXkwy30x
LXDC2lxy0+Dg6GKj0kKKLWPhhksdvOQMuYMaGsgScSytzyOPixCK4ZcYLVqIDBO2
q501GJicIH9ImvBHvj8pHDe36a2MUEZ2ch9DM1r2OckpCeCVU04izld0+z5761eI
u9mIy2zq5lFGH1FAYqu5Lr5X25pAoELurA9hqMQ5KRg21sV7erY39/ZoKP58BTPY
nwJsJwkKNmGmjUZTnwYGK9YV4/9oViRVzqnU4yMq4nH6GsDfx6P0IssQ9ciCQgFY
drttBw6kMdcaEPMXj0fvJ4/5hIAcpKijmYgRZ8uHYJUG7lsfe7uiTA7KasyYJDfO
Uhzvy3KFNbfPMvdZwUHpsvTNRjE6RpXoM5HqVbJ0gJqbujLVR/eQXm8pi8nlBj2A
ipyh90WYN2h7zQYjx68h7c5gn/pwoNyfo2mkFs6vGaQf3ZCIWZI+RfuQ8HCJDC89
dTsD2luA3XFXkW54h11HqGqbD3fA8n+L00COKnYa627s5DO8EoNHrHKveIDmd3Tk
1GxtStz1Z7RAYaj4LPY9D/fJzckQSK4k8tPxD6+FdAe64Fu/gaI1lH/rWs23UUIK
5ZJ2cxedUy1xlDyU8IJFx655VsJk+6ozYNuDYWw+fy8+04qeoRrSpUwoE6xgmnZF
yxRXBhDFkTeOWrIOealKNKQWA4hactVL5zvCL4k4DEDldqrFai2uoNRxtLHoBUO+
V73fGBpvTQszIub6rJtlf0I6GVXAas3uzupPY7Uh/Uds2LRYOD/sErSEK/8jbgQ3
IS1askqqsZEhEOzmStnGfw==
`pragma protect end_protected
