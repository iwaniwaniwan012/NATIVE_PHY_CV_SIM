`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
luUE7yQXoA3NKnvDrR3c90mrlz+KUh02mQvNrdBx0+X9eun8LKAjPdedW6i19c8V
4LQkyiNZTNtaMAtuxpZWAAUrYs4SZpgPh/Lz6VtCOUtOVxJfATERx27MU+J6M1Ha
x3ka7VsjnVMWzgJbZ9TZkUB1Jnksu9aqpICAoPL2iGM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13104)
GyI+8m+Aqi0Aii3DxYnCBHKQAWz/UoMmZs5S4+y+i/QSHAZWBOkUV4Ik6m+CaOIf
ccfNgvtPi1ihVwcI0Qo1y2f/0SjXqFdZ0ErsV91wNucKqGE3faMNuiZP0s5nwfTP
RdV+nzbFqsxCPkOSF78UWwoHNnjwH3C+ij13gG6y7zt7N9wP61xQKlR3kt2Or5P4
JevffkDBHhd+jA1hTiI9S9+yK2WK/+WjwkC0xVFhitq+wDiVOCQFswUd9OA5IHnN
Ket4fAxwt+jDk/fIbrZ5/+NiYfDFut8+hmCtJD1wVN/TBKDh3/YhkS10IFQuSkBa
hHS6+9Y1SRd6H55hQZr+AX1ELtzHfmUKi9KJDGiSCyykJZ1em4gbsAOxmGpE19Pt
7LvdhWY/HAm7b3sh8ARQCupx5qY9QbojxARoZ7CZ4SfdpjWclTBTVFFjOQpVSwHE
aWd070nG/6i5Wz3vUV/wozvslfjfKTgBrxGKnLuxaMaaojohEglPiHJ8d4dB5lma
QeeZGwV9oZxymOmM6dsZVxOqzn+biF3xeaXoWH3guVkL9l3OGEUxGlsIodrK3Qy4
v2Il5KPhXYzzSoCujtjyusurdtyEcLOs5DgMG1BfUb4kkyOki9pEt7ecZlATvQMB
/5xwk3ezbdnozStGTuzO8iKIoRsQw+yu8yQ2naSuTMdY/zMx/SQbW/sMfEhohG4G
FtJAy0PDcXNtQpe7980hWxZFus53qQ8Uh5uOu/23mDo8zhGjs/zdCuy+Wj0sqCms
zQLT2nupMeGw8aB0/9MVmQ4hKaJjgtd/49NfvGttYOZ914dL3bayXyRvxbAQ1+//
lJBSd3rebxbMZzlT6h7CLk145pIhx7nWj9q/hrGA9KovwAWVLv/ANAk2mr37fNeB
zjJyace66hDkHc2C2Hox6Tj04ug+K1GNeSC7zNyh/QFznvsY9sk1kSYylRA4RIAK
wE1wnBx2EDCJFetEjO7+Xa3XmdXnSDw8z/fYUjQ1/fwSN3wjb4A+6JLtrQlxqP7w
qnNQQLFzfQ4qTcFZpLtOSxcP5aiA6UUvj1bQ8m8K26K/dfsF1YjrufiTDICaQVWt
MlEJAMihlTsTvttSIwF5rfVp4UDlPru8OklBhw5m4yWPz3SYDIGwVrF9gBz69bzb
hVa2S9QwQrHofCAkp2T2MRnVQKBTVqV4i3YQz07ayuT9A7Jyyi6nYLNSBCqk6UCy
ugOJpPNrCMmQZkvkhab10BSduFLq+95HYUdgXuHvy5Ja0kGD62WIWtdrs8zY0zLN
hS5Qb9TXPm31bmYuy8mQdG4rsH1zznS7MoFLwKkOO+sXN8nqEICUk4eVBZxPMG1v
LQFDM0Tpb/XicCZFYoLeG5W4QJCgU4dGKkPHj26k4+YuphkI2jAo1oSp2sjgl476
F5qnMpVGmuqYzZRZnohXwqrW3GIUOw9GY5keltrILaTERz/MhWRr7AsgLWC+yZVv
pz9Pee4yYxf22/pN6pRSyiSXzbxupPOTg30qxwYnHjmpW9NXghTCYhsaXqsJIetl
9gYmZmWZyHsOg1QHGiCnqVcLlprERNoJFIURPSLUs2iIcX9d0tGuvbRy5j+c3gLC
3dztFgVxp12gQ3uFZZlWQ1RsSBIYYzR41brmWFfyFLqra2w9bt7D1+wCifajNo3/
uXJOI4gi3Gt56Rdy2a0K+Ojrzb4bqkg5PZHY4DmfU7mysT0Dc80F1UwFt3+2H/Hv
jxUeNpzpBh9fNZZJj4T0uk17BKToNQ8fHOR3RK/Rq4uSwQcyG1Q0XCi03uf1kQsy
urf3sI+6H/4DyYKRrDypSoVKge/sqao3K+aFckGD/DZZNNcCVivM1EZmb7qvh7Oq
GzjZ7lUsU8tlwbqcDlj/zsw54YgjnOV/bsdf5hNluZ66GsQBNDTYxLVsN3+mJCVD
NUfw63qo4J1esMPLzyA3UtLxRp2zFne0h8oe+edGYrEgapLCOASvXRTfKIqxuZJl
MgRmAACXupksj9kCz0Ax6Ef5E99jAravF/PDEqSL/KlPxtKXIUhM1aO1hW8lvwB4
ux5cwkYhLiinoH7NDmY0xvSX8+YSewoVUVS3UM+SbXq5cTdzt4Yp7ABQxoCxa8hm
MMJBe0mWdK6/qfPIiDuWcWjoBHAbTrevySA2TViuuu910qNpopZYKn0viyIYGWCP
6t6ilvmRdGxh29k6TU16/qh53tQNE5QjUjek2F/8smwDpqbiXKK1VRR7DVqsYY6E
o7VJnOhx9cr+tEIgY7ydWKmnLtFedAESO86HCwmcvZbqRyw+RIy90m9JzCF+bg+b
iJC3BmlEZRWbSfhBzW7XKbY8mGCM7jjtIMhRBi+wviiy5im5tSNpMh2zZFLBr7lg
jGgpp32ZLGjfPqYdoqUrCvsBNAk1E7Mo8YvgHLic5S9Q1+Xv5kzHySMw20tQIAkp
jbRn0Zzs4Z8OGSL8OkkLJOT6xK+2/VH762WZmqZDzFSSZ7P/h6BnBMqmkmbxYjkn
w+/49Ugb3O5Pg7X9pkIfAp7NpoW1jejRNw5a2Wl5Ya/3ChPrPzssUC1KotS5EIJC
yvh000jdk4VHOwxZCllf4zvpaOS2fqPgo9gEkpqT4IhM4gjSujHOmZGsg1MgmFHn
ZBfoaYxENxUa3cDCYLqqvPsOUl+zmdFN4Wh0mx9XR73rbhXi7f67jhGq6xKWT4sK
jURriOyfvv/ynYLPFMP4BLIoA/SOVUOerNKhyr8AnGOxIOuAkcJvCJQb8L7EKbXH
k6xr01/9pAzM1yvq8oJbbNTngbCJGXnhtfZs4kgNAMseaWKqdTWuEQA1iIdTtyxt
wXzo7VlYF6X4lpp2pHTf8k0z/hExwJZj5NWLhc9dIkdyn9K2jmZJoXDC2HOfGex+
quglaXQ9EQso23hZh22ynu15sxgY1nVGQO9N5JWzms8Zps9CseRu/DO5fP066W3Z
TiSUphtXUsSF+e2Ps+waEwHvZwQ3r8wPk6SXDICyyYYYEig2Xvxc2ob4a4y4i3QU
HOk1Z/rC2dKOsA6KE/lVX+Ph+IzLSTCLHQrZUI4P9pRGGv0EWKoBncj4InM7mIMD
gBWv8fJzRcYp7eh9E7AKOGXsRfMtT9/IcnIf3Yr/acwQMgnS8ylxYlndfq/4gVD9
lZHPHVrlrY8SamJMothJfY9ppTybwUuiSUqOtUg2Xv2SS4wgFPqRHz0od8+ELP7i
qq6bIh+Sn6eiAf9IBlaargIZp3nqRHCpaVyhRgvdidDzw3zDGePikvjQ8cDqu5xJ
l4OooUMsCSOKua7Yj1JU5dcL4Uut8OCdYsIDvL+oyBSm0vowuTsDXlvs8mX2tSy1
9YqsMteLc6Nyde3q/PfKm4+z5NFjZjlXTWhKCumXTQ+H0ulB8xibKIOsejEFosN9
yKaqsEKSsdgJ8OJPGUDL9zv789SZWqZwuxuX7BN97HJeHY2otj3VVnCqZu6PqU6R
PcNXtqNcxvdte5AqbBynv+lskmw+PT3YcdSEUG5NcX67PquLF8wwu8B84III9WMH
PLHB8PuHhsl7g3TnOwl+stvXqQumOJGTJPlcKe8ixLSo+0+5/J5GaIBS9TKbLYyT
useS3RywoFq1p5mM/sWWIJ+BmCnFHEkMSbnZqnbCgBdNe8RIeFFc+2mOHOdqg+AW
IsfPq65teLgwjIZdMSsTEKMPripCGpXHbKDWgl+Q4vEl9M4XkpDzcisi2u9IOmt+
8h5REKz5RQMaJBTlQ83j6c1o/4zlczd58CsCz6o5qcvflYG7Mb27acB9tLHd5Y9h
MXTBA1orcMT16+lh9XzDtBg8Nzz9nLw6+bQ2fGCW5IbXLYx0+C+mUL47TqPFyDtG
13K79IwW3s0PoOF3XDKBZuTdAeYkM3U1jL/IJ93eQVlOb3OERApFF8LvjhzccbMg
YbzgtGOjZuyp7YcjvomOYzzz2oTafIqylaTLHe420kzBEhXdRw3gwdBAVWNRlwNI
tzxv9/pYLBtEwjKGfXxTBkIM+zU1xc3YvVuIQkZ4MBnp19MxOX6KPwJ2Y6eCBLZG
Vvw4Bg06BA7ix8xj/TObGcagrppa7aemwKthQz2oxotYgsXsEVFmrLL+N9dhkgBx
xdsHdwM1dQLyYoSRByr+4mgJKghI8PG7AGbjHFsyXFBcdrwlCv8T5xjq9F1ddCpz
ESHrH3BLAc6oB5D5WNVxX0osNTghfTQ2Ch2xN9jD5c9MHw2PNHwL+URMJE8yL1sc
fcyY5ZNJcrbmj1wKqDfhxCLi9Nryo/9KVQs2KaP1vUdP7+P5qrbfdr4XJ92KD80L
cfKrzUAkcahCl5dZE5gYszuU/dO++yGuFXtU7emxGNfnro135OJmckUFQfSc/WWu
BcIQB51kHb6lDCmlIcS9Hp6YpNMzWfeVUkdbKVl7IhZRBnlO6LXNFPbaeQs5Mk0A
OSwwIhQ6txfsJgNKFzcPZlkSmyEKfbZnsbML9tx6f2mx7fgA+FvLUCQibPE3hrho
TgYRC4IDvZMiXKc8sJ9p1tBqbDzKHFGZKkVA6qSX0t5sdzaHGPOdDfi+WjEOgpCy
OEe6SSKhH1DTgC0XrgiKWVt12iMLDB5X+2rdVmZDlLMzsFkLXdYn/19X8Fztb/wZ
vHFqlxXsh/13fpxLddnIfkzQ3G6dsAQtZ4g/eY/gzt0FQ15nMEJe0tyytqwIjwQC
ZCybDPbxjyiQXCQTJNiaFFCLiRd36yiisF02Cv20i6qO/TK63W4pMmK+rKqEtIc5
IwUes+ukVD91YER39iYaseWsnod/8ugMLFRYYoBiS54PASvI+P+U3LrKlZHOhDaz
mRJuNxDKsmOcC9LrF7aoYCxHLPlD06ZtIE5sGY/gaewL9hrHrWuVrL+BDKYw52aR
MCR5FhAa6q7TDBC1E6R7FtXRLIbE1bz/xFtiZGGahgY6MagjkuCuGzt38UqlCdsD
u5/qMqA9IN7Z8sXDQF7ju1SQTVUbG6ttlHtxM2YfwNskf+IVE4f1BmSowvnjw6Vp
vQtFY6imt5g3ubKYkzIia0LIEVGNhlNQy913GPm9Me55/iyjm3rNuAPcc2k1Lymz
uziOIUwEUbGptALV2xmFAnGBnJx8P5eRFYoMsyZ+kD+DFX6ICraHphpzYpG+UJQY
6vpyoUjvsjFQRrwH12Ji0WWXijGkn1kLLHqlEwjv3cYfRoiRNWBujgz+cEsg6C9t
/3kiODVLC5D3JfVWSL+o6BCn8U0d7LbrU480BBzagVC/KUWsiatOi1mveMW3HDle
WJrwXRfDyZuJN0a5PCnjjFc//hMDLp26ROhwrj70UxONz99edjPxiLB6m1BlViVP
U88wVqIgrCuXHlCZC11VmudN31qpwkMP82FBx1uNuJdM23w/5TDg/mEzefNIgSfV
U37bGxSD+Uxm0CsSSf00RpGO7R0ZTxNgbZYgMIaX0yT80GGYM/uC+Smsbc1kL+mZ
izdrP0GJg8kcFx8x6ND5EFfBYyvhXSojvjIJg0Z5mgVykJKo77CBYOKLh0nSx2jE
mbPamzXMPYQjKT1TKngTKrcBcSH9qUb2EUL7oCfcL5yQ38+SczlPj9BwHjeQDzkU
b4WWMzU3M4SXorX/12FnDOACPqKkDWYGUfTelXZjsrrZubw05KcPUbmanVn9fx4Z
F9gjTyaxipa96YU5HlUWkRcZ/uOUkPK9tehuhbmHnFx7gNBwlMsCu+ciXrGxIZga
PE2irbsgGQj3ftG5/0hIDggNi1EwioJX/FhQvdjrL4l2XekdfViCaxR9gCjlOcae
U3/wl/0MQ0bi4wh3z0PAqhK5/HlAb3ysiuxcATeqgyRSxk8Lm7Oj4d1LA0HLnYdL
BJ/5LPVVzYym1olgNnP9l2ARAa5wPgJLZBYspRP11DmeEZWEx2m1Y5SdHliY4MDY
LGTj2LGiuJcRvKF0apSsHidjlHeBv9KFYWOUx4GBBu6gsS/crHCrtRitmy8shHK7
arQY+wsfKRjKQjk7aUJMZguLA2WYNoIlhDqic6XIs1V2dbtzI8EstJrOYnexBpCS
fWp0FgkqMauAEkVUjaLhRA0SepshY2d+2g1SPG+NnUc/PoQuhbB1ROCNrMu/hq1w
7+6D98yo7E9pemoOpVks5X32T3BxZegDEBaFYPVKPgB0kKTZHMTpCNff/iS3jwu3
kwa2ZbELbyxZ9Rmz+NyMz0GGc/lSyw/+8Yp3GtP3sTnw/jNb2KlXhJHcolcAgEg8
hkXzsK7/PoQxxRuMPSLF5zKfL8o1zXvDlNGfa9XaoKiewX9NNI6r2gZTyGVj4RFh
zw0k6PhhhEG6eCFtAL03+flWRv/ZfFLe9LX7ZxTTw0RMGKKXG9rI4xrlmhY3KP6a
yQAXD+l0RNDASI5KO4zixLCUyjPSIAYJGmbbhJT5YBs2yxJK58ulZ/vH2jMMVG1K
5scwDcILn+QfT3OfWe+qJxzmVokv13uBaVs0CS8ei4XLfO0WKdiZ+N4jegCOxFtP
3od3pzOSHLsio9D/7gPgsgbUZscNYqtOjpLLD7HFDPzc0Qofg5mCWfTY2XuegIIR
tVEsV+tfsjlZTFgKM3W4fWHVee+b002EpvTt0mNWx+GlqSmrSrJXItQdFpu4LuH5
J6xnNtB/Z10OnK2pJVWGk5x4vziK706/BEbyFugkyhJq3vh7s0JX4dqNyCrEVJWd
jZ27WNKVkSNZoE5Cu7DdmtNWsjpwfRXs3GsknhPMNS5pb1MeI+DJvq+H4nr6xSs6
fxmt/ht/rziNeC9Y+UyhwgBGOMIXpxgkKOuTZodGWKq3ws0z8KXD+aXxpxlC8Teb
um0oVpKHkqEJQbAwwIj8YIMwPGJ4W7wYV6/vKy2fVc36v8sMf8PgFL8ekYo+IE7k
uhOtGyNjCkWoKdabp69Eq9ovXuyGRJCWmhvHg6cthLNatqtqL+QXo+XolnlYe9uG
Rf2OWL0AMyWmnmIBT9zFT/ZlvHkQvl7mvyvxF9l5XE287X9pPHfv9+STByuZGlY/
wiifcxWffRQIWICLj78Z46ilG84fbFrhux5I4rlObOsYWI7IoFsjhTDnhEFwS6q1
NRwuVVRNL1EL3RgrWnjNzifiHKXEqHeLcfNBoHM528JM167bspkecI4vnFmu6yXM
6fv0MdwAF4KNH3UW/TvrDxPJMiZijT3uOVLaEiY+W5OQUVefPsmxdQ5vN+YLNycL
WM2uvow264xWsI/JDrgBIEz2f4q2qJH4yly2EBo0D3chg7O8ZgBDfc6RNE1gxkRL
Hk/NRG7qow+6GN8OPUua1Zl8+m9/CtH8Laetp6cW8CVwVweUhAagynhsp5nZ26nn
Q4n0Y0f7beAHa9Dz+4F9JN8EBqYR/NXGQwxi51cijVNL1ZDAWeVC8+9nMpdRiSv3
DDhdIT6l9kQG5o1H4tkt2JnRiGJjQABYnNbth+QM6W5BNNPdP4xl2xMPVaUToAra
b5/+dcvjMhdBT8LWHKGEcii660f7PK/TA9cHYDPg7ObYFC8oaiEjzmIDSf/HiRVO
l8/Cd+HobqizYo87CFjNKoQLt4EP2/iNVfR3bF3vNW5dRKW3HylMZjZTo2OTmNCR
Njl/PKtAxncaerHrVnbpbFrp5HIbwFeewN1JSFsdYEGQdeyVV8BddCA4wyXMO7gM
jElxCuOdBd+jUY4kTDS+n39pMIi9lz1WeQiTgs0nA2P6milEEndc5rn1YM5fRSLO
kI2glKd+lQITbBN91bePjrND8eVeyXJ+ZUjVOJXCwCU32JAsAiCsVnb6ksfjHnCZ
8eO75uhIeOIW12SefBhemQFZnSQgrYCl2De1mR0S3eBChwgpBpkC8rCnYaq9KlvG
Ci6MTLavc6RT86cDt1Gzy+f4Vyo6NGX7jXaZURF+iSRE8Fx4ASU+wG7peG6n+Pw6
7TGFNjWmD2CKrcHj5Gp6R2+LGxS5JMzn6BOrTdmuL093Y6R2LVk/wCKEgT1DqAkN
Jc/FbxevF6IXwOCnZghT/aQzcQasxGNQx0CE6pcuQ1tMSaIcUMdGrXo1m0YKJSuK
WOtyB2lR4OVNxjfQaI2FmXQlu7FXsANmXkWHSbpPxn5qd/VQARN2mteCBDRa31Fh
NBc+Wc0xsHvLA581RCPV6VQTjjD6JP8JYriHFXBq2LGjbkJ97wiqIjhzvpZ5YE2V
9TpJS6ial8UbSaiR4iBJGBCpOauLpmlJ5WqA7zeXhMhlBUV4lvVbyIRQy6f81IQC
ztyxumWpiNfjrPk47WbcPiUHWCLBiM5fNd4G/498ipOolmj0whQ5HKBpruAAghsG
6WhHmpezl2QK/aWf6S9d1M7ShLC8cIl1WbgBWf1WrQ64ReuQIJK23H0oQtxvjszn
TvnivWaRgE30iI369fTb+y6fRIpm+xfHsZ6BI5j+ug26vdmlRnx23yCB3Lg1Wfqa
iwKa/ZM8jv+VmY0nTMj8XSj9s4nedwBMW0zFPr+5xs3qF9zNscLd50oO9yWwlGHV
dnyQ//jgwQGngV2EyNcb19Q8IUMKOfecGkEKZYD4iFnxf0Iger64HMm8Iyrobt1o
X4Cxclv4gqbr3Hyj3TIE2e9pWVzUBgE+rw6jLXf3I7UeF19e/NzkS/04H2ZMVYnX
Jcp31XAknGZKJXuaAfik0lYuxlDj1RcPhCW5hyI0C57sS5ZYfX16v8tcHCP7TwbH
zzphqo+puvBiJvBPNLO50jlwgEOB1i2XfjVLSwuIlxGn5Cf4CISn33ZYMdPyIquN
SF8Br61DOYSAWBIrOjahFmmzloEKhU/4JpeoTLiuOozqUBBcPQITltsTnkYANxW+
5v7Dn7DmqNlA9RlXq0PiBSjs6Hc5jvwJuyWZsVPjbj+JfuHgHzrZTE0xiBQqk8Nw
oaw7TP1RXG6Gbu8HtEbUrJ0EbORaC4m2uZ+CHCt/BDTPdZw4S7aMUz73Zlj8JjOK
R7YD6Xj4to31u7SClNmCOMbuz31kQKtr7DvW3LL8wtpNLimejq46rNR3wALDXkEL
IQQvNDHnlhsFSooChWrRSZdP5mTAIuECkMBmpzNoZGQJNNKTe3Uo6jynY4CdUcwU
TDJgt97KVZCMpra3yLWekIyQ6qgLgZs+RAVaV0OIA/cWqWjf6rcyuijCU3wXjbyX
ElgKRdWoJWN677AT096NGuAtmBMH7Q8dhPNNFC+92IekWjgWZzkjeatiaOec5P10
MZaEJXbJEuNwwYvye/ANLoJLAcRtf9rGWY5XlhbXpnIm3GExicop6H8ZcMQhk3hF
40q+cdM3f/tJ2UAKUt2C275GrXFOBbJN+DhU208YInlQMv0pNqFp8WIL/ZhGUc26
IoYo/0YEA3Q8Jk3XD5iKaCAN8s9cpbYl1oPppu5AbMQh9+aTIR67pCjj8tBdNwKS
VPx9/tf/k+76hL7USXtaKkNENp/So9NrwtXmOg2tg8FWekeM1sAfjqEmocpo/05r
1sWumo9bGHhlTf2qsubJ7KHx+HXRG2IOSz0ld1GX5kUkZOMC4cTb9gLbsFeZfGjU
0bAd73AoHVhJ8Zsei3m67gojtw68xi8fSP1pAPcW65WvgBmXoZ9lY1+pob96PPNd
2/GXF895JlK9RQwTM5hHK9PSS8q7z+Dc29JRu2xCz8NcFHRHBpZsehA1CRb8jv48
MUQv0c/E701fSFb4g9sQsxm3PiP5pjKMigf/Z6ULPbOeSUa7YfnAh3/7A0izbRis
G6wp/x3a6zjsBJFMp25+netODcQKmbBskeCy79nYu3Cj0CCQCXPY6+fELAtgkddl
VJg+lNyWMc2y3crKUmr+4XH6A5b7GkDmwImoSVXANkwH4BFgHQ+wXtvoV+4efjzu
RSuKhA0lOsGaegJ6WPkhvIIld1cgS29oWfHmH6jgFI8/roef3YK4WQAqaZP8WHEH
Ztx/L0z3skYYowVOxd0IQI1CN9qeBDpSAfsyTJxqGnHjxyPk55Wn3UY19KEhJo6e
BZeaqM3Ye+ET7JYHOi3HUjdSommcBFuU59pDyixxTIxn2zwzG2eSSQUA8YwrsgSX
QjhZEszTJ5E/AvYz0cJffYnbvkKaQiwK8erXXrdw6Zq1poVC/UtYrbEpeh+7609L
rMuBcWYuBCE2RNSLinsKXAwoQnywYUTocbR5zxSBBHw7XKeeVeabSod/eGWjhROG
oOYUDCWFSuwk9CvSFr5PFHmGTH1Wru3D4HXSCthtpCENVEMIarbydZmQOqEcqA7V
7Yzy6ze+Ag9Q90+TIBHK2KhDOtrDTKNWsJ95YWDt0PSBft5V23yi7jrdisNFLvZ+
PW9Q8Kji4TXV/+Tgwxez5ZdQwWWTssR+V6+t3m7j7YH4iNpSzgT/ufMA0KNBvWak
+qLLWkdm+M/gx4jCbuuR/XCIjzu2zVNoQjg40nUj6xaR7ZKGd3h7BXMNNS0DG85Q
sBq8hJXHjOypAdxkJivJ6lwPG2BcnI4GpFqZYb4D1Ib9/dRusp4wVM7aVEr7uj29
X9LExJsGgKiM6zALCCbIWliNtikPEE+AA7ZQBVix1JBE3TruQg9ndxRV9kmPu2LT
HkxIEsZE9HDLIlghDUttKzoPNTylEO11zIxz7d/0ifnJVC0qlRDA/j9hETHxoKFy
Tnc2tG4Ksv1Uov0QwpZiU6ObSFGbhm0kdzucgC0HTpIeYGYYWbpy8l5mUKewMwNH
ENQz1m8EMXLD3ZYCtnymK6Vkgp+LOButSgpgSepeDJQSUho1qIr+74DG1CWQIh3h
BahxT5QKyQvnde4cdt1X335fX/yTAUZ7/6eN/hlt0lNZHE66Dcw/8/QEoa46bY0S
/CVW0ZDBs4q5vRmCnnHKeO2v/auV25bfy82Y/z20nwlzij3hvyvx+t7eMGWBgQ+O
HsBXOyg30oUTxBzGQ5GAc9PoYNiMMmXnbS9roZrcwzK/wAtmSZ8//l4ZxRNOCknP
utWHV/p2U8GNLHX8C1fTuxsQl6csRUeDoSjOBHZU4PPGQp0UeKXa3h5hzG9IQ0Z6
ETnMpdOm467Wh3FoP7xCeVnlBRaMVdl7tTjX0Pb7JtrOdW02y2gexyWmSXKcCNTr
O2k2daPjGO7j7jEAry/KzVypuApNEBEuYNjI/iHSBIS9UkA89e52M91E+p9OsVmb
xo+K3Ujhpgl3r71une5fMGJJnEkm7iSDZvCZwZ513bqoS3gkMXQ28/1yY8YQbDfK
RBx3gNWKS5deSYBM7ApcCIjCGp/JM654PVKXYr2CiQlXJn06POHHshXYaUg/yOwh
m5hy313LsVQwJ0fU/b7HUDUrBnHPdlyiupibpfOmqlX3IXKeZaeJpmV3jlfSapvu
xveZVTYdj2qhCokv9TlxHtP3d30qxWwwquv3vj5It04gGWwU8ieGnmCfVKsWl8tW
NQIGUnuuJNdaE0IYTLHMjJHgCSsx6xiEIzUSBtRfT+F9FO6N5gYDRo0RwHREFhah
w2DHoEPAsstMRkT2LhiD5RooHKReFHgj8NVXRVJgZVQRVZJXDhgK6aecTHMgvZU4
EDodw8cfiDnm483Lbepmlq9qGOVoRGR9LIxUe6973hmu9y5BSeoaO1spe8teBPAs
VFyIn8LPzwtKxH2bjwWeL+1YVGZJHux8GuGfLUl6AlPdrYdh6MSn8/fkcJfwTxXa
3AiARJVhXD98CDd71mztQ+eqgb/c61Yjmv+jU48Bza0uHe8OL1Hi8mAXYgIaUytf
+218PWUz9gWcJieVk9FiSfOJPWiBj7Hf/xX+MCNA4j/vtFh8IZTH3ctGngN5/Yfh
ZYTJ5BRHDp+b79elTsPZLcKFiRhg77yAW9Buey9UYfq0MXFge4VOxaAQwuxSUOdY
vdK9yMaBNVvRceLAN+6Otu0Rgh/iZx4EKUSDiNKidOVLWo4Jd3IHCJPJdKlmZLZ4
Z4iR5QsbTdOsBAECmCa2o7D3fDTl09i2m0lk6KIjPPjxVa4BnE68iowqV4FdM/9m
Gqrgz/5jJJQ1bFRnkwVqZnCJCgqbRKDcrya/NlG3BCjjBkM3BjrsNTs+MB8dyV54
wAXk9gpaYqrU/FMxYbIif+3t3dyBFVSb70cmsOZwh6Dh1IBvZrdJrWwHI9yujfzx
/fsJ6Hmd04fdeKYQhNpsaNYX9TWPE9hbISIcu5PmUWLD3zbE+oThqeUu4t5blLjX
9xqcpxowTUBwhnPJkbTYzstEx5WyTE07rqCwdbVTzym5X1f644MoZoP9I1S1xMtt
tzLnmbswO9a0rACuWiCxa629iv+MZLxYHnhn3R2zVYEqdg3rEZTgxyRkSfRlmFbO
NRe6Lf7NEa6Q7SW8dacPPxUW0w7bH6o7n0INQcPQ4qNxYUMdoLdYpORSYsnTu+oU
hVRpnFZ7ov8c/kZrLSMvNlA/JNxikYylba5jskC6YqtDuCtYNTQH68WFfbqdLjUh
iB0I89wOxU8LTVQ34TuxC/uRoObAeNA8nxgqW5dmj7zo+IXkG8xBPqcB4FLlk/pe
WL8Y8C8HTx60CAKrHYCBjO3n0LdHiE8ge1h/+1unqzStW2n1gEF+P/qovuQI4kFt
5W4u+gFtcKzuQWvpw9ILjyMG2baCVsf0BBbjo6eBkhptHx0rFGPaIOw5wL4pRyWK
4y9IGgFfsVmuMq+qvXxXc2VBYXtWDUM+OC+JQeMTbr+hKD56u7x7dX+g3oTi63WM
OlSCQ4UgktPA9Nw+PtNcAhGAI1QuNNv5MTqrNXt0jcfYa2JBL7FamGQfth0AGiR4
xtO2MUNJVPjDsa0ZSZ0OcwYvZ74PR6g4e942HTowwqEN6Xvig6Uz1FCR5QyFFGKd
WLteF+4+xMq8ZvlrhGm4YOQwHRzsmiPI1TgtfIcxsZZ+5IjU7y3LFnzRutpLT+8b
zREQ8mR7evkrN0UfS2TzRK9QYM7UHOetF3F5TanNn8B31RPPxjiA60moT96+Wztp
OHCkjEHQ0+HIVWsiRnD2VuyPXqxLw41BY6vUXjP1NeyIZtiG5jbgdU00gKceut2/
ZGkZpNMNOtyYTMnzVukLYS5jqciVeFb5SHR2LWqn27s/4QZ+YJqFwT20XLnHlDof
GyE/tVgomt4AR2sSlaww45F97FpfStqCL2TPhA2bmOkwNIRgb2/QZafITDzwjjcJ
uFPzaP9QLCtg1gsDoMYBahNn/1eem3OaBY4tLVTdIjcsUmItLb6mZ1d0EYGar+7K
imYp008gMkRQeiWFWB3sObpEBsainNpF83sglBzX8Dna12wq+9+BpI9rQ/F0eLOj
fb6M/kq8xn5XoIAXd3aOWthYjnufS879JTI0Z9tYorzwkhP/ci+0V4QPPRFy2l0I
ZH6iFq72uZGOyir0aANyfaqV+IZ2VK7cZXzXFRouoJ5JAL0FljoEnhrJijr6Z55G
OBcidg4JPvPKTGqE2XTCEkFFLkoG240k498mrYMRxx7ktBhkbtG0cruXpjQifyg4
S8y+ClVOo9nnBcsyRoLcu9ndvupdyzSXLreBLCMlc1ZIUWS0vrbblHpZoGd/BEil
QQrpiCtkRn28WhoRKPbW3N459I5LSkpY//JwY6DcnEkD2x9KsOlWPYJcc9nICeZn
XCx8O3+OB7oufbvzHvRfFI2P062x7WtVTAAFhet4Wt1W/jppx+IfKXhub8SNf8CO
WlLnxK4dBk7IdEuzyv8KZXTVCC0gehox9S7gb1RrypWMm/8W1Hq1asQ2/GSF7vK2
FVTo/Ok/tYP9F9OqJzIvMO0XP0ma1JaVDjw+KR/Z6dwEiXjLg5I/nSOX/Lv1SEWu
8BARiJDu4nJjzfevc7kyjcug+eIbsG/DzlB/pPpHQSz74qCBgjf/MwTfBTLFjlLK
N4YTCGNC8+ZDtVpjd9KqbL6IfDFXtI/wo12GWA2benEpgFNFJisRZmTepY1egFoO
46FJQvbs+21hVfZFbYeRKuaps5uz4JLEl5YxT6bfe7ohxIpqAtIOOGNMitTHv8ap
m0tbD8uQbyVNJhE8c8S5FOZZ1bFy3P/0ATVlAWesYbNYgxO9O5FnQlVR1jgiy6BB
RyV3RYwxvN/B/ukm9ZcYADiIOCCfPxFc/XezkJMZIcS/iFQfIfVCg+R1CkZfyuyo
I4z5TBPGU3gPSteNuLhT3l1QtEdoBMIYhrfqFGAUYXDIx6Zmnq1bZLPpd+70cTQf
gMmWqi5FkLjV05ImnlEEiC2nC2IGnRcG6l1YsZ0ABaokYqp4nphP2I1S4LAK9oi1
3PidPgeb12ZNKx4AawK1yLLW8FZD4fgM6DDxpyr63iTYHW1MwDJyhKt85TRqXSB4
XVKxbGNHMCwd6n7x3QnzOiFAg6GyipYiHNcfabO7HoNuiw/vUmerJEwXBLjYHbS3
eVu7sPAVEHkdwMoW5b5lU2oBD/ahMdZ8vH3skD3bf3JYJgE1k5138wGtpEVv/df5
vOlgnXY+d8KE4tvFhaNbD7LAlRUbllgPvemX1fp+p2K0ilQIKmoK5QCKEkfYnIJ/
BIm9WCka+Qg46iJHKaftr+Q7NOW7cAmtLazXJGmTBpKnJ47Evfzfbx2j1vHWtlhQ
EsZkBrXe97RY4nJM5tA8pRM3+k74Lcv+zjLDRYTzr/IgdoR/vwBAcnuk/uGpK/vG
m6J3q1qyHk4js7CXg6k8NViG/Fs+RLq/nEwk/DrB3+N8xqkSwewOWzd/f2mUv/ay
nLGAYWHkjppeLQrMKx8dVABOi07f1pyYmZMY9N/Ck/DVITWZZvtW/jJNjSY6xIKK
aW2yLOB/7Fzz4ka1sNdhu5Tkui3dbVZQ1jclZ0jdNyVKjwZuKVwUYPQhS8GJ67gr
rEoke07EBYH8Yvu+GUyRCFdIfXz/Po14qpoV9jPXHPT/+E4BwJss+tJNbFHR5VSP
wqjMiyYt0J0dww1lWo10M55qIFPqvHM9kODJfTZScAOegF5l9eGgPMfMcEbW7QHF
xs21AQ1vh39C0n/DD0sTvzXst2bpeLZE7S3QYPrpJffG0WVzmexYuuCNLsQNQn7N
tLdGefnVYStxlMSAROuxfg2rZ7hQJtWk8QXsx1PXQHQ2I85yf5ImBMX+MJtcw6wC
nt8snWwErGgt/WUH0Erhcr+bxXFOxGxj+DA3Bpmh55ZM9IbaA3H3ie7pmRMDlyWj
NahIc8X7X9V32uMNz6ldBjNFlIHtB05Sgmf2JNqppWVIEavjIhfvCxF4wMcLEWFO
GNibFhsgwEC/dkwHJk1YdeeffvnnjokBM+eIyOC+Vnipaoz2EjmkgQioqg/ILd5s
ZSbyYQp/dZ8KJd37XCo28AZ2O5pLO5DKZz2O3wTHxs98lQaiHipgEo9iXrh8wWdf
JhuMEyWhAEvcZZZFMASn1WKtAfK3AK1EBbZ46VL4TEUXjQnqs1EC9soaSyfY4KTx
QITyy57AukKUgxGuHqvqmD7OvJTswfQ32laMB6Y2ziHtmLMlBpLmJBh3jzpxOXbS
KVjp1XbYZp+Hkv+Go+Fh946QwlU5cZaOHClG57nixaqSQPLbWRQQ/yGIFeuxHiRi
f1E+XfIg8I4udbiOoYJz/XnjF8ZwAmIwBPdCMP602noSvWNGECr5bpQnvxxMlLlD
+A1sBuivc0lyhhXkqu/1NRsweSHv2ke48h/CJ82VL/nEDePcfg/suB8qlbrrh3M/
GEsyAJYMc04qn3MNvrggpNx+yIdtz4IlXZoPyEjyJu8bj6pmQevPpr7avvyI0TiE
ktHlSg2KuTPRfj2ssQS/lHdgureYtzviUXX2WyYcQmFsm67R7okjXoppXTZXMC2I
7q4YqnQcaqP6a1xe7VpvVeEqiG2ohKqF0EBl6mYntyBmTGgRcOR8WxvIccC2Weyh
mUxt36yJQqUOKQKgMGzSx9wfghs9XFVxPDn+VkoroigB8hcwFeytUfASXKr70snZ
pcTwq69SBoVvVSdOU8cyilEaMCortvRws5+hzHJc5zOvgbeive4a6T0QPFT4AoCB
azFuaWG5g9lYedhP0lOtI/9AgwU5vPaMAISy6UWYCa2jCngXJfvEcG7jn7CRIqI6
S26lJuvj53/BKXelu9rJhVoPesaHC6SeLtB9CYviwuKR5rRFrS67iYikVHPlAH5H
r4CjlTikd3xUGOYuxrAuiW0eL2Ft7KXriELAo2Y6RsN+u2Z6Q5CkJm3boldvoExZ
5hyGy2Sq8e7AQqYQvL6fMZMyP4a6J+dcS+P2GrWuCJByVcv7ywU6+q0tReiKA81e
saNuUSwmmORvvdPnyVNY4IXP4PXKw1brCzDfJ8YUsHr0o245OSjeEQIBFQOMxyxS
DxrMQ3R8jzcpcTWgxazfolJ86ttasCLuqaFGEHIJtIkUjZC1BfV4vliW0fJwOa9c
GVpZWHqbKg2xC+y+YTdDhj1N84x9aInFerdUM6gfLmoYBPXmFnbJjc0rb040imbP
5WQFkrGEZIE3HHvycN0c9zqPqc38weub2VLADbyFso5oi2wrGbi6TRu3Wg0X7zlf
hznBrsxzj2/xG5cLS28A9oe3AlnQ/CKV3p729enVs/KZTNTjw+co36r/zNP6kts1
YfO9DQWiTyHtW32tAQiZMhVQFj1CdCgbJx1PoewDESxzKDx1CwU8M8fwzyUhqzlQ
fBMimSx53IcsuZ50r7ldu58CY6MC06sfhrh+G9DDPG5GJyxKg22GwHkGoc980QNP
8j2Waqj095XjMvG9NKY1pwbS28Iq1b3DDMf3wXQ2gOpZsKVCl7fzPee+LtihuKgr
SpNYpR0EahoJLTrmv5EJHASygF+S+WKfC16P8ve/GrHrrvgnEhwKKDw9Zg9wFvYn
wCzOWsZzZSfGEThQM0CagErxs4W/WawFfSK2ly4oXtIEyhbLkANCVSm9azicF0pg
oifjQrI+3TL7qrz8zTUbwhCO4SGf6t1xoNQeIjRMdQ0hR0EVkOtDHjf7IStSe8+s
9Db5NqhvjJbzVUp6AxTLLtSHoD+3Uqlk+/c8PC/Hqo0VYh3pJWdMjVKw4I4x6D1y
YwZpGX06UDT8e5RD8UnS5nPcr4q9EebMFTDTfB26Jb03ikave211fcW3l9n08szX
/7ixgUrHkSITmOaUOzRVW3fgUpbwOSwMC203Dj+umbYfuH2JJJSadynMll5TrM6E
47Q5Zj3rc8Joby8W7SCQQopVz1AmzTfxLYq/2mYQisaIdwcvycUshZn1reVKPVP0
zfng7i0dhMtmO3dUZ6BJ6+wUb3xnCTCdVZF33vLjLwYEzaTC5V6+t1dxAURK8Ssr
w1lkrNTwp6ml4Pml2ZtXU0Hhyat86qZS1UXAOPAGD0q/5fIC20dWMzHGUj1FY7uU
pnH4giZIxhHAf0gGhOKjO2BPAHhCoP6aun04xHn+IwpBviEgOvFWQartUV9f6R52
jx3Pr2iFZTPjehzI1SCLpWy7KBG1Oa8xXD58lKdIunfriDQY4e8BVv1bGmsXNZHI
Ua476GI/4jLxXY8ICMj6zAMGdO9yjQSIRRf7OxdxOIzTMcm8PlnS2KPHwTQFX8jr
MBDOD1zrPG8myqgNeU98X8olDHKmUM0vBAF/4WrKm5VSCg7j8TM2RirJ3nawNt1W
`pragma protect end_protected
