`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UmcX8HqLV9AF/eW9ja1ObWpicWB1GHM0DerKOnhkubaWStficRf81dgCAwGinJaV
cpcJZtxOkeBnQBvQM6hFykWdBCHw8COo6IqLSK7HNtGio1Ity3BVbTrCQMsBMyUo
4Gw87jj5dOC6xJsVK4twMp90ZKUM/2wwqiMujY8c5W0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5072)
GbbBzLEXL3vYWc98ip64yFPWzGjsw4dNYSNsKgzw9TtPY/uXbpGFhI474nE+wdsH
Og5/eFVBZEZ59BxZXFV8V1jsjSZwj4A5VmzgWuT+SxQIGT5WaSJTwjnUL026eUJe
TrmRqrgqtjCidCNdg/4iYXFLcmlRvUgDFAcD+Y1vXgAZhBzAUoDMA/+ipwXpARsR
VttZyLeuBGWyvCVY9Y6UOfXGsfgw//sEuf43BqulHvrL0dRCaPdScRFjKixXY/6d
9QDd283jrmA19VWZw5Zv98bf00iuklHvOISi04jKYOwR/HyGTB/4a2R9Mjc+ofEr
8UAgA+Ot/tQaB4ykfSJN+bFKLPI+x559hojBoJm4l/U5ui3CT5M6A4Uv9i9wsKjB
kwmswNqdF+xQhTLLGJlxoOqQlVm9cMnQ0ThhPJ7yAQaa/JtuDpK6JmFdPsFFA7U/
eewCUc/5GZ+dRTw0pfBiLfwGdL53dbIxNFIP0S/24CKqBt4iyR7owoaRcSNN6J+Z
4x/vXEYXtl/hBOKbAD0nf73Ke69BA6zt4iQo5DIZ27W8mVpX5P4MHBZjjTh/mwdy
6OXuFTg3sNKeQ361WInUhbLtMdrS0DIo24bTsxf0G66Scaqj6XNGVTc5QFnO7Loj
HyKkbi2dOKHo0TxZnXfs+KIm5GfJVFz0Oypavr3P2LESjvlnT2eUFzAaLmqY/a2m
XRO6bxFlrMGSdNJSvk7Oc3JsrjWGmXgCAHE9yLgRjvfIuCwINx2T4z7UNj23FwY+
BUOHXb3/jxpIriRAzAeGG1dvQAQkLi02xBPwHPeUDHU9vi9Jz8RFoTYN/STHPL7K
UxHGXYIx0m2d72ku4d9oebQRp+vNVL42Dqj3aWbgXWGBGN2rD3xrnnqwQUpLlMAd
ym3j1FaxFi5xo5GFQKEx5P/b71fCqOwwfEZ9Ww7cxouoKkqS6zvgoOngQE98VNk+
vo4kmdCs0pZTfaENwdm1dvNTYTmHiZCpiC0p1sTm/n0ZvymdxxZo71iE4QrizmBS
MsCk/TyXuQrtuAYDWsXZMZkrsApqoOYzarWt9TPYyv09cJGt4mBubVsxKxmguzDw
7iy2Leo0Q4VRmb4SFQcP+OtYBaw/2/3EP/YD/jd14bPSfmxYXYbFvFbtRLWTX0+b
9/UN9yOX2TaxY2kmtheg0RgD0Cq5kjM3vHjmZny+F1s1NewE20aLz/U8stTEe67Q
PgkKGCkBGDGgXUgMVKq2m41lcRcINCusDKMwzoa+0p55nJLzhO86YNqSWVMXscmy
fM0zpEwTqYTKfC0kdavYtyjQ8HhaThfQdCA7hEb4IvdB/6J60D+rD+K1ij5Pk725
atyvzEhSUzDU+3EIQF46zgCXGjCbjhBOmKu9cpJV+9rNEj8j56hXFKGJeFFLFVTO
F+76czKeRgx1vjGe8pyG8vHcopA6CyQpVlaVdnnSeNw9BLrQpCLDpDasSrrgzCLU
evrGkUL6ErBkPO58IRf9O0cP8iKaAhsvh3Ooibilqr0wJVcR7H0lc1jsTeDgFea4
2d7vtAWU4JiR7xtmh8kiJeDnoYYykRuKWZngYkku6+xVGBlyc48vyYIh67uMSdYB
dTnA8PQ2GtPwrb7FNZszI6EdW3vXDYnPToP8qDA1t1JrGdOvgeiDtRBYkB+RUnrl
oWFm4GVMY1ngaNQUzFY0CapWx8R8taB/Vb1NdA3zWJC2wUnazNXRqp3ThuHlaXQI
audpeElY4+zR7iVXhIrnrf1VDxoa72O8b7AQfwhyX5LJ3C2ie1QYxPz+6BBey2aE
xgvxYrQRzxeYJf5Njxh+YXrFRJiu6DO/KUB4jqsBDX/xU3Wn2Op6IsfX8kzMeDJ6
+0d6oXtvahjvXCykUcmcZvmFYVHEkzo4WV9lv41Wz2ciKzY/pB9b7H8KJJg1IfmT
Bk3Vs3Ba8xRMlmYiS6rQ2QJMffxPy86tP7jz0JKy7GUXBTvkMhzxehnpivNyYNqi
wv9Di3kUBRNYjZ9wfLQ/EIc9zKzr/QTvOxGqKSub4rnG/xhNev7+Jprt+ZnUGlfj
R+Z/EJZcFLmhBiIiOLngo8dx4q/2XKK2WWLKT0ZsAPX/9ArCtxQHysTxJpB7rg5X
i/Uu3G4fVRT49Sr8hz4gjj5hy5kH+PODYt5/Pne+1ZPAgCiltQp2YjbWVdSMODBP
dECFYI95dg32nqXyt+yUrxMhJfEYqXLdrd4FFAOU0J0aWsgqOsPHvWSn6q1JbDs4
h6Km/l2ZrvJirSl3P2Dsjq0Cau0vOp+drcJ4HUXYjDhmyQ6M7zGONQvjh1pamBQv
bc/HogvuULEQ2bRfUFjzQA2xem3vB3OJdiDbAXbblrOcMtK2sse0GztEz2CrTyX1
jyrZI1cHvY4Sbe6FuCcWWvYS6qd4gi2R7xcJReEY6UcdIHEtdN9Pv7VzCWuycVmV
Yxm2v6+viAUjt9U8VkWPA5Qhgb5UF7NpuVOd/VDwLQrbbHtHyjV7LdOV8r9Jizfv
45+8GrGy6iiOK0Ahgd2lieWhcqUrL/xlrPY4oFSPBIQ83VRQdkZNbgeF4jt6hMZR
q5WF89NP1pAOY11YXEJxsJoa6yNb6Bh3NXDivz0W++cVeq97AC+W9mUuytew2pD0
GEmXx9CNMn7RL4Vticg+S9iMSsU11rqslC7R8AjvkoP1HBg4DsmotlhJGQJsvSJd
GoDCFbGxadwXC7WWRfIkcZR6UY0wgrJz7TluJTfwqsyt5ACYVCr2zuoVgEC0L1dy
l+L8h5YwpBMthHcot+m6aX4xsp6AxRnbJujPJvgcyj5QEOALrBXpp44/sSl+tJBA
K2C2JlK+Td6FeqrUucdQ2494UTo2a9eSjfdKs4eBNFr37ZHecUAcUNh2wr1OFp8j
rdmsDS/hHJhtxHu6dFRrSXHuy7d3dOoskUOzUMd+w41oqBm2hH5dYIa2Nm0SWcUg
Ngmp/hNGejt+dUaDL0tlhevBAStAO3POnqy4dQdoIVLkPCOt7Bq0TiM65M2XtBwl
9ncPeDAr2WY+OxsQzpjD9EsUSvgCmlnOD7tUro/Yie0/PmbMHcj5YN+iKLbutW/g
8WmtCONLBm+/MnLQoQsfC7/hQVQaz5elxCPfpFJGAPMM0hdtYkQQQQTP496NosnG
wt2JXjaTLaeyj/+Fq+sYDEUhtMhq2RwvLk5xf7Oo5g/mVlC9Eo0+DWsAOvRHde+Q
hoGFAQx7n+pKqW4+rOP2+oW88Blvg5OettwiflddAzmQRRuLjxmTqG4GfVe//d5J
uSf0LUZuAV62gT/GVdZfBhVxOClPKAa3qjeVpVKp4YoanX4u9iPni/aZSFU7fdjy
+j/+vN0RNEpwj563IDBvba2kqYSrHYeuTtnSUATzjvxMof7jFbfEj37Y4HUc1aUK
lHQeli4Szn68Mgv0YRXcNa82LfZ1JKYqW63/cEZzGYwlapAKFcaNsUMsw6KJArD5
PT+9iCRZX4cacHoz+HELK7PPH3oxP5aH7w1X4+NrKCz96PE3NC/4evV6eb/qdBhx
c73y2u8HnGw7YI/SjLo1CeUuBV4kPBmikyYKLC5+sO/3XxNDNcFb2wpXMxJTj81x
8uFm34LSMStK+uPeuJ+1pv6wkI47sCiPcCkPCKux9Ua3CjlEzdDmXMMJtENC53Gt
kYeoIZphwZX/ino4Nm5uV9aYZXYCDeGfHY8dcdB87cC9gzlfww4sqz4lvEFYGM94
xxyenkGDFlyQDuijGlg8gWXv2Mf50a5WXViE/J5m5lkWKWi6T6HAsi5lsPa3e7FK
JpR27ltBbFQdlZgHB9qRJys8bjBSGXBS65+b0agCukz2gDH6/vs98xlHhcf+8+J2
6/0Tr8+eMvcXQzP7I3ug4NfCj11p7VATgYpJq5oKsUDr8fB43skMXgfrCSpFHFtD
aRLIX67/FDv4P3/o8figN5XB7FYDITnHP7iK+ht2hmT6Zr/fo7RXvB7O4LCX5b58
+j9xBv4PnRFwVVVRjJkahATnb6uNik8ZPlSULBkQLCEoQrRAZ84mxxGYqdMfJqWR
/3Wf7R0CedKjvSBz9Iz93Mi1iqN2eqhnIdhjpoljKQr2Bk7U6XLcDnuGUOJVCc4H
RqRNXtlcAlAg3hrcdSZmtG5b/7yTtotduU+s568rDN/HJTbdzzzXC2GOaqYarG6C
jxGhhClV3LA3a3KVqO9hb0CZnOrOaCR6y0M1XDCGh34/RWAq4KeEyNmiR8wKF6bU
E2CyPv8DUPmaHJjMsWZbC8Q5/3jeFOnhcbKO5NKNA8BJkbU3cG5+VMhbIyJHuWVE
GBtTS9imSBruurGSTnu/7q8MxXW8hyyXdt5+xMhW8tm3h8Q3vRS4/WYhf+WZOJK1
+37WpeBvei79mutYBMBc2XT/3FKGxssYPHfmNtvdCo3SSPG+vPYz9XPNU9yI1F5f
FRwwzL8aFpRNLuLj+n02ltAWzgqcvBBVn3FuQCogYZipIjQ9QEMApelORo7a+yMO
aEW7hhV5xqDF0T5D6s8Tagm6KQrjLraZp5p8zSdgkaudiek1xsk7F/Y9sMeATsmM
lUdA/1CJc2RMhTBP5NoO8mq3YOtLBeh8FHRV14MSxtaNQTy7WAhdjfzlLkt4Q4/0
D9OgU+UrORGWRWdkdArC0l9ARazpEYLQhBVWvHPzofXUSWR7LZxV8nFtH3L4XI9o
Hk4/K2yiJlyAEUVa91XD88FocWMVCXynpIsX1QG9tXVopV3F6Ufb+yCrPdXW2C08
bH64k+YjqT06Zvh3utgyaUiNz/b+6G8jrpC6luMJA8eJtbSfL3to6OAUu+HdulGg
DgQFZkGtdYcXMXSz3C+46x2Kqus2g4/PtAvf+tTF16J8kGsZD2OE0/mVNCZ7rdGq
GA2hJih/73jLlLLB4JDGsYVWB2VuO6omHsIEnBQJyeGB6fJKu7NjP4lza9J8rI2D
AolKfvwe0VD4CmtGEfA74pYGgYTb9Dxu7SXjl1V90GqcbABz8kBd0VkrlRJaIIou
FK1KYYFX4cPHi6hc9JwI+TgTN2E6gMoIIJ23HX7HQ4PHLoHoOmvNpNIe19VhH9au
jY37+YkzOJFyZYDvlmI0Azy00z8e1M32w1vLsMED6KUDC0/Jno2HbuX0a5nFMKrq
Ak/mZvSt8luwyQ6/z6PyZP//e2MC+hoZyUoADjkhulBnA6+pMI8CaCsMpK+KenQr
MKDJ9sdd9swLx0W/ND2Mz9KZpwgL9QZR82YGf/VrV9M9Bur6hrSRoMWwEzrqcw6X
Y2DK25zjig69NP+vRICuiNesaZv13mzuiiXqFAk1Vgfpk6XsQIcchhtXt4DULQ1e
JdOoqvZ5ifrJYudZ3riG0qAcBRiCsm2r/w1NTF3Pbz6K3CPCjxW6SSA28ys9//Un
2P/S96wj3pjmIVobPEm3i+YAXHNzRKsu7RUtQAzn6WnAvtePKMAPbUDQE+JoZpj2
MIKR7RctnQFiIcwzN+kZLYmbn1hHBxtORMObQWD2iaHpIVbttOsuxEU5HjlEWUX5
VOBUws4y2cfZYfIEBw0NwIeKaYZr408p4WxwuKql2735Sh4O/eR3VZk7B7E/JlCa
Ozii2ntU6quPmPhWq4lhOVwLKH17AM/hvDJeEotWgILEI8z6nxPx8zKhCr9OZC+g
tC5zpZvci+zM2zWOPPmuXedcRi8q9bSz4GCHPHNml2dfzKnYtmV82zuY0EUcivKy
FqIkqC+cecZXHSyuXmvFcvuhaIIclHUIy6l2D0FvpoyyUHv9sNUTFGaU34jZ7e30
TeZG8YBQ59TA66qwkRpgWgE+V58a/KhzO/4nnpBnN0QdBcuDyMnHlIneAZ9WFqqu
FJ8Kq63b9fTQp9oklcf4gboLr3Lpy0P+nWSKtZFGqj8+BqqZKUxrXAhhveMwhnLL
g/X1YCvKYOGqi35Iv3knaOtvCkd3ingyBzDtbyh1LW+kWNsODlP9jXi6ET2WmIHT
jv2M56XcePr7Pz/ksSJl1JxRztsVFJPlOXQZdcNCy+x8zWFZ6QOVNzRftmPiPxAm
vjMm7igdqOr1c5kLKuaAXf8XVzU7zq4hTLxVj3XZATY3HvEaKuu+aq+hZGmdzM4B
YRummCnSHISrUyArb0mNcXub4JGs7f9GO0twG1OY/LKFMcxKr2//Ua9IOKCpkV5E
i32RG+QBGbvKMOAO0krvjL5XLzXL8jMUdm0tFttqv81ykr5I1y+T7XLNkxUeFnwu
CZXx7tmdyUASkzXyE2tziJWH5HG6rr+bMFZXRBmV2JTtYUnwAgsn/iHOvtzYHODi
+2rxOrfVkSr4rianJtZmATwVDm8kGh1z/vo2XpHUpyVkOy/rpik5ahNZrrOSlirD
T6zyg/maeTBCUxv0Jsyf9Mwjrp9SIeo6qnevlgnGPNSXuabfhbIaKvdMagd/JOHq
HKGo3AgzCL4vVCryzMFXTQ2XqTk6wBBC2E2JfWiDNh6oIRLRcITzmrXadyKO640f
QAczlgduJkjErP2xenoF30too/GRbq5TTStI9Uzr4ffw6aP7YF3e07SXaDWooPz4
0Sf8oB5LmOwvQ06IpultCSNAkVL3JlJ8NCB+Gf2yEsjqoR1wgTPNKAx1s4fvf705
G/hCna85tQHlou5wQz7cInxu7l5pnNUZmhhgy4bGwKUNKvPmIrElkACEYPBAUr0D
0wuWe/+fS1gkglXJFDM2+G9ts8zxJtgnoB13LXRmAMPpO/TTUMZEEau8AwmMX4MH
ecybGsfK07Os9lRRVQZEd60ugtPmWjHL1Wt2fL+W+Bg=
`pragma protect end_protected
