`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bCAUndH7EQZjGo0djTHvCzh79c1Kx7/m4d+gx35QDRhPDPM7os6EawsYOsaio9tJ
ocKOluGqNOSn8UMCfufRa/wQOwKVKDf+/nXt5LVKDxG7voaYLv+8EFUT/L+EQZKx
7T2mMLOjBwjPAZHIRPs96ece17Fkhk149RVQef5iOH4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8048)
u2OM15NQTQ9KanynCEh1HZgV7S+GxQDu0J6lCD9JK7zuYEcnk2ai27XrUNyIvMqh
8usW76vA22uMibou1AdNZ/roJTnoxYUfDpAPw+5yw6LPbbmOGEyFjOVk0ZadXvff
1o5+6Tp3jJD4zbo2k5QW1Oq+nnD/TzyRSogUmn9Ltw+DDpzsmcpgEwN76wpXSgzH
4jXBEqcVKzeLmUwrSdzqL23DH18kIqVkuFS3qybwd+XnoB32lKg+cAIz6WdQSVLC
Q+hDtn+TcdXlmIjhtUP24Kuz2XxtGys81OTJ2ZLmNl2j7u/YLpTBy/Chi8GWzASZ
d7qrv1sgTjXAm78MGTKM3ZXTodU03y7F9HkMew/kbMwX/Jv1Pewj0C23NUkTMXY0
1MxxRAmjMjjthdCxcDTPoZfEV93RF+njFX/eNj/I35TUZh5mI4kj5oNwVeJisUCR
Gl340NlW7UXL/8IqLln5syp8UY2FlzH36kpOaGb4ferKKINYUPc14B9CTvDpGz/f
HKRoRfNjWvphAbins1tazQRKYejENQQnnj3k5wvMjhj5hSWq9eIBbkZBQYFmgxI8
qn+0nbiRG8hAOozJkgoNZEeT6IDsq3Q5MC1h9ZTTCYdYRZ97AVJTm8GtGjXLNgpP
ejjUxduUro/deoVtJ/PYbGPSkB5U2wKRty7uw8cTN1uQ4pQ3GSiqMTLUydXId0D5
X6RBvW4MxhhygA3wP7a1S9XeRPY76qYnel64pMCFba6bxkP1YGiAN2L/ZLowinO2
4wE0fHgC1oiAJuj2jElzBqxKRNz6tgYF45vFW7Evv7piEWJ1mUexdRL1ZBEBqWVC
BbApK84T7cAQdnzU4Usqu+Fe6xRIQwwlxLbBytxPsziEqMP4oMUUcTrZThvQmEXp
+Rl2qnjQ4I3B0DzqHofAdSHCoEJ+CIBB+CDlv7qUQvXcaG67cak7zACL5vUfEIrC
XVdKLqcp0u30YnCk3nksxcj3V0P0rSetTR6gi27QlpcB0xhlFJgwQRFYmXOkQo+R
UfXX9yAY9ubUCrZQc/fH5oiUS9FxO/pck8C4w23rsv88Q2rOJce6gwzGwuPQ/FQ9
3ayHdPejm44GEQVb1gKdKoeYlv+dToVtkkUid274fdaNDGbADz6/DPYlWGejGG2t
d1qcODV47lEy+BOg12kjWXjrQjwDuBKhzlwxx/jegFyFsv1bkTQfF5HCBEq4OLiZ
3+2OGth7TLER8OcVM+GNEO9FkF3MRLBMlr5ENdQ0mA9c9TSROp83/iEmYUR9tjj+
Y/T1FJO+AZ5N5onKh9felzNRqYRQlxf0JjnpRPl3QjlKfEQ+zraoRKDOFWnUVhdc
XOxae56tnhTH+PWqM0i5J+80VfNniuPynzezzhfJ47FtBHTDhkFta7BwvtE6RG6+
aDoGvLNEgI9FyLxkyU9cbvQCWHCIvbz15CRXtzH0+FIqfdcM0PvOLDx9Awq+Mbs6
sO1VqeNxY+5ocLCPemWemxgTw8Ne6CaZcXfvvwYEasidDlKBXebHce3rcYzq5l2p
BVPll0dA2ZuvMbNeO0Y0TgXrXX4j8HmwYmHbTMyyngp5SFslFVp6c0uYM92aq2AA
L8cH2Oh90Np3bYTculbGMlo2If4FPX7qiJPM+8tGqu/kto2rgEVxgze/d5Filkt/
/D90JNQL/LHyiBGvopzglo2s6VwmEo4vWghRpBX5yF0joDbUaXTCvYJ4sxXALZ8N
RBZTeNXTdaSVUU93w7xFrDK+0VlSqR+JquyTcXUTuNITNUoHzJInL3DppDEU5y1T
tumWxpQYgApsfjbDd559lG30VHYO7Y6FxU9BSPA04x289AJcrSFX42PM1JCPNT6N
ids3xYZoSCYZfPvtBt4cMqjnSAta9jGG9B2SXlqJkQGwMaECt//2NML20DL2Oy0F
lwVuTIRW4Jbu14qlhDNf/S3vcnANv+O0iZz/2Zl39yWc+trcUJlk2BZe14Yb8Mrr
uhz0yuCZrzxgC8z+DOrb1hr/K3urxD7UQfh+32IptZ08ONMW9XlyNhaahqY3y1tQ
VWAh5Q7XB5UuWdhnzHZoEkqMIuOysJInoh3DRc9VgcMEXnEdTHZ41x5BDer0NcIj
+AGIEOKLJPwBu0pQOrlylfendArrnwvFj/EDRjhQqPddsZckIhRJnBA8U+pyIKOE
bYE68xR1wcPnaSeQuUR5D1J0rPf7rPztPj4CkvxL5L2viJWog+qXZV6pJVdO31VV
pi9gQB2Cr42N/4W8MGj6iHTsSkBsauugTuJvjrflc+HRzzAL49iMxR8g4mGGiAcj
49s1DlHOiMePY5T396yZzC7YKv6qYRspmo5SL6vTtClMya40N3jKb+MYGO/pIDFR
McttN+9jdvvSIodq+S3pC1xkukX4lA4w9csZX0i7VYUv4h+Ro8pIYFiFUyyv3NOq
BnMwEicUJZ8hReQbHxIQ3I8DBebAqK+eSsr+0dGiFHvnay6dG5VUDyrUt2c6kMth
Oebx+OrbmaN7/wDOMMYoGmC5uR5kEL+f6yvPPjcGQLkQmRgnYg8rnRNNud9FfJM1
fiwz/vHx7B2IR66TSL6Ga+ctSVsj9kdNL024gCAhHVqol/lWscnV8n6QtiS8SKmz
OLv02r7c81BcZ6FgJhCcZb4Uk4i9CWfT1iky9IFPm2qbbVXhxsrrDUMW2Q1e+vLE
f7PjbWntIsyHaVe+otf+TbiRuIg4aOtt+x4rZO9U3FBEKkAuC/inXYNBItv8sEk1
I+HwFB0wytmymxLeFsyRxMsTNX1Bb82dYNomH4eP6+vsoVHQNIubEQY34Mqx5OW5
C+tOM6M+u2ZbFvxOZHFlpjmAE9wBN/VBk5ngFrO/80nghJiTxtrQa8eBHfnzXK6s
M7bRQOUYzqhZiOw+pVBE+KG8Z5+hZS1Yq8+ft/J8vanQInKa9xBtTkpfCOm7Ht8O
PHFsg+Q3SxVHNeXPcDqRax6T+o1BeZ3paAD8tBNNGaaZuiKKbswRJ12ILyikMNb0
6W4gnv+QiISJxFi1gOGPjJauBnBBR3VEDLo57IPB3Txqj6gIdW20WEgivVYZ31T3
VBZVpnUdOuxiU/V2DGL/acoUtQ7vb2T1q5P/bA7YQkRjSFxDaKK3v6679gOBOFkV
0O9mzPt+4vDl9WZhqaa+cu13u7zfm+B/XZul7TkmQPPANztVF6hIVBq82Yj2mttp
UYbirSNdCVPrEB4wYtVBO+Yi/kHkM85+zXBD8ATKWDiY89Grzdm2bXn4rYxlJUgK
Wt5ibfH+6S3vA3gj1lTG/wEMcQvf2lOj3xNs6KuxjE+PJiJRmC+82TwFpWUsRHbF
+K8GYoUMP3ufC/sZY/87lR/GTrgSQpEG6aEk+Tjsh9QFmn/nDBfPaLDDdWYGcWNx
hPSAEbgjeoLiQyvho5S3jlh63YZINmYlN9C5gOgOZydwZLQkPwXy/+EJAvWW91z1
gRm1GuzMYcvFd/3/kR+eAg9Z0h3vRgSfo63ZS3H52uTUs/ERYHVgqEs/pqZw6Iws
N9HqmKiozcF7FdIHTgOh5ZdkXU5fkZ16XbheNHa+yxp3UNGyBGqfkMjJeRj0WbOr
RaUXyQidn4r6hzhbxxWpEs6AeC6v3PlllJelv1FLC2KcNHtdKcKO/MaEhswj5y2g
svrksHRNlAOlmyRZYZZT/fRojkrPAPtI1ok1ixLIwVdfrkRDn2ooEOSqNvePLlYd
IK2PWJTf+HyL9jZKwLHSkoeye5I5B+BMfumW1W9WUkUBCE5WnmcDEsiN3ntfH5v+
DCMr5sRSBAWUIK/LW4PqaEf3VKAut1fVG5jBY/3wpUOyr/fDOqlAfpTgUm8XkclV
91wL3ymIpa0pbaIHdiYCCBjyeloAiLT8uKhaR6gf5tI1DbdAVxsrZFmD/BzW/LgU
DYBxvL0VDMVb/MaqlPpCi5cVeVkxCVLFOA05Iuvez3dyg81plZhXB7c2s3lkcCOK
dxtWCs2Fu0dBIMG1mqkBFAFbGcLeUlQS0UOC1Y9t+yNzjokQzpu0+hHNjujmP8X7
iLZR12/IYHhXIUuEnkK/bQVFs+vOD+prgJRg1l4XCOpgeIbhbhm63XHkYg36BqHS
DsBlMB/5mGg2Cwaa4VNIU1mtEVEXeMuh+RkRGIfWKAcHPbLO4HPzSZbAE1EsyI47
oFgCaWUgK6zv6WTHV55c7LpOtTczPN6sFXpmxY3lvZc0dfzP4tetviiYuc/kyzTQ
XaJAgeoEMseCt1i89FZHe5njsaSqTND+TlPGHOzUAREQ4n6c8bm+dxiAEqSy6PtU
3lRJga20GsNdA6qMVni/2DgT2Ra5dZaUpXf6zcm+c0D/HmI4mkX1ZFJpNs3ei5ih
9f1P08Gqa3BqPVJCzMxXNzesR5WJPcedVBXUxhqfARgRsdgFwBrOzh3aA5gWVfAn
7RlYy95v33QrTsGJPv9ej0ixFNRJVrP4UDkUxiLjblY0bJNv0YwJCif645wHaY04
nVYRoyvcdfToQPrZrOg2E3QYTIhjVQ82+WLdQnEkWnaR3QJmImpyllVRa/icAztC
cCCX6dCIKJYplYse0DQPkgQsHYcOd7LE/MwXImFDVJXFtvcg6Hp1JUmg+pUaMnmD
HZnFy3cOT0NGyN7rjC2P+dXB7nc0m1U7yZUELmBiFFByNg0JyBQsWKNB1epkK8rd
e1PPqbsjgNOMbrhyqG4UFcYNX0b/RI4sRYX9Etok4LIBNnOOSTd8vnZW0/+R2JhC
80PRuHOgEGaHB1jYV5PXyuUqPYfe/l9zC8YYG2qd0I7tot/yJEpyQ5yTpNjM1Q8I
ILdQw77741cASIqATQYwxp4AmOk7at+ZDZ89F3XUnNnt+ge64/rkQhhP8LHL8tmr
PGqAZTy4DuMaPeMeXWE54SRrpgwYH51YQ5MCGqiQQ3MNvawcmbE5uG2tKBvGKenn
TlsV66cXNiC2XC03Zw1Z2U4g7U4ht0oo4mPgBhM9IvY8oCDAtust60gOaflqg7Wj
NNSM94GM+cghSmO/DQzFWu2owxHipiXwEDx8FNLFBT5Rrl3UZBXc9TsriuScNYaO
fifVdvJpuaGMV2e/UksPdEapzlKpKJ7NisGiOd0ztDdi9eWzTLdt0a3/ZNtKC5YG
fFBsmdz7ZpNepHh5PnC1tzdukxBth164zuwgX5v+ZYM4qGG9ypL9j1GS1h5BsvH2
1iFJCWQg8ZKRtz6AILgqHAWZLrqehCze1ERozCkqoWQIMrkW6Gk+SlcjUAkWuaVs
I3uPcJxQmY8MTcSUVyE8NstC/oe+Tr9LTssicShAhv1boVG7gmvaZghMRV5dSPcG
hpa9wPoGaICgeu1Xsimv7kXs/kuievXp3qpfPVeHSTN2PPc84nrSvtF7paY0yYI0
iiZGdmCVVSff63MYy4Rdbb4BbPkm83Vjn0ozmLDVf53IzwaRcnQp4apaTVIXuQ69
rTb7EkkVXd2FV0siajOy+ef0Dw/dkLP0XJPDymkFDGfPWjaeKdrjj4cW6W34XaTj
9GKTgzKX4dChI0pCdsnSNF3qlgp4qKRyM4VDGrhxJTD2CRXW+rjmMFjO53xjIw+V
FaZ7UiV40J9CZ0fz6zbOq8+uD7jr5C0PGFEkEc8WGX1fuHtCwcir17h3lh0BHPEG
XpaWZeV0ADLOOFZadu+XhaLNo4e1WPPDVcAz3SHZ9bpKnQoYvLK/YGdgljct3VJ9
WF7sL7L+f4LDNX4wkOTdXy0zbd/TLUt6serjR7NAJorbEB3T8jY35uSO40UWm6hc
0F4oqZxHbiro5Fu/x7k4JAdvwVGAJ3agB5Tt0qt3gpkLkRa/rUwWxwJu+6/R+cro
iDjuH1EintsimW5383CYJZNByNhJk1UD03NSNfAK9RTLhB/EtrEADu/EIrmPoROi
ER/3wOpKkrSgLq6rID4dDqd3CPPtFIHiRYxe84u9c0UAJELTPYojffI7iGs9KVe4
IDcQDjhLsFHUjlRVpywCllFYRn/JXVPKAqdVQQBqrvUv8LwiPXgKEFfQakh7W61L
OI7AHf62PbVLEBBW3TSEH6xIMkTQixBCAVCY8fj5P5HD2m2y/wOCd/EPn/0ZKtDe
XXifL8RqpCuSQagwnimi9rxOXSXxckeg/XgL9nnWK0NsRrc96Ae8h4Wsa1tIC3vO
dZ5dVxNmRTtHTrN2nv+h6YusXn1A9dM/xR8CWhYYrhXy7hu1Bjk0qyDlkbbgcOc5
eWz/Hu8+8lJfkOBTcWsASHRoFw9q6LKTtylbkjP2Cu7cE/Jn5EHEIqBd5c3q2zWk
ImKzgNDsqv/iKAW3QrJhD/7eDsgvnKQEEZ21VoPf32DI1a/DsAOlJGx7B3gCYw9N
N8fckhLmVm05EcDGM1fKcErGTWY9lP7zjmKxtGi1K0uSRunFmo6XfyjFN/WmxQ7/
Ux32r059PZXcBtcYd9UtVy24x6CFlMUIYZHwvWhBtA2cbovWA01VB6pEDXRJDBFv
upnPz8gv4iCKf0Q8lhbgOI0Uub8Am/xqMoIVtg2A7uANTUWkOy2waOoaF1VehmAI
rVf0ehYm8BgTWYaK5ZPi/uSAZgOEjsZVgswHgzbNOD+h2hSE9kpOR6F46F5vvWVa
JruMO1KOZWj87Oo4jPWAfcDNv7iRki8YsLDqL0AxymjLR2GAYUZ3Jcm5QWDE83UJ
8pRT1PmOvIwq3+eQLV3ATZF+u3YInG/Ef3rtHESBGo58zRLjP2cAbit1nkfKVILl
xuEnb4hVMRlpF9BiO2VPo/Z9XUXpL3EuamD6GcBpSd+C60nXhBZDBkosazKiGD2g
LfhvdPTspsrmxViBaBP4h31m1N5qEP0hMSqeHvjw5vJBcQHRJUcgjnpjxsFsCYsS
BCfKXFxun5IWwwqQqbDDVmVXFLE5ImibOfPBdjVb00fFd8n6Af0NORkLCfVRIzTS
TbEegL7UKz7greWjztFO+qN6qj1HBrNM5IdTjT3msRiAKObI8M7TlRQj9mQX+n4h
SEg0toJqmU8RbrIkIPOloIAeyf8shmJXHkATEjLSUyVPdgM0LtNssVuqopASVGY7
s6MNJPLnt4vF/s9t9A/Y5aYbxNU3Qmtk0+Oi+mLBesntFo8/hgFlLgue9ClKDvmM
aRxQA1Uy4LlsZRPm8ALiwz2cd/4A7ESOsaKq1T+ZxcuBCOOG5QXtG3BbA7ouqcxL
D+x3gG0YwwOgCp42YUZWbHwTfEJycTAxWSgZK6535GpLHCYMltGJZdi21STH+K8u
8m4dqlg2RJGSoCO3uN97Opd5HOWgh95nApNLWNDvUcXcb/nOuAs0rzP/Sh8anE60
NaOxj4uicnxLs2SaS4bHB4mGJiRMMshrpeMvVlEAbaSq/TYs2YK3dNpJEsMPJJXZ
rsbCrAxc0AtoGjo10Swx8XWSuapO+Ao7Uof3bpdpZgVmXxUzuduqxwhzLQrItX2F
RN2HfKjaWBExGpHfxFERUSlJEx1leKcnGcCv1VqsJ98twD78R/mCNgLeyWE81vaA
m6pNRFbo3jTHNPmguWGU2UY/mFgc7DTKgJQpuAmK49VAVCuxNibM4oioA9R8UaMc
q4YKP0q9ZvZkX1VxBCxMsSI5AY9kRM9ZpO2MIMfapKJDzaQhHWyE26Mo31z+8Pcm
81KbGeYF9sMV06RFD5pa9SEMpZtpPJ7TI8hSLszK5Af3BKJ2KDG6ByTcSImJJRbQ
VqlS8fEqQfxitwxLezx5NdkkuDgWJ0mN1lAbL988UBXmYoDhXPOS4X8uZR65acD2
WNMsw7siCWyxBy6QWamH/bn41Fb6udAW649+DqJoUZ8mcPtJj6Ih2Fvaan7jF/Or
U2kWTrP/teX9WFdkAPaBHykwbiRTDMFaA4PNl3sDZOQvrHGH1yEK4t+dhjZfpsw7
L4EsCLYVrrEJ2Ot8OW8mnwrZyUouZ5cZY7aQvfCjDFDNhDRRYcj+uujD77NsdLuX
gQGlLHPhWeNp3TU/KsAUo6KyoV0dC+xVmaN/lBefMc84wRSpJPiclzunsfgtvept
Hw887zHoA5dBiqwxebT/mbWke8fzg4g+/aSkdgLDe7weNLdt8TpVOq6ID3OoIlDY
3RVLIV/NPvajvTrDCWNlwO3ldvj7VUEMZY8yoedpwVjae8Q/NoJw1jT4P0Kj+UvC
u1AifzwR38tcLIpeg9uVS01gCur5mIoOv8NXeX/IpCC6BXMD+NDbu/D48RW+sQ2b
qede7yCYf8uVYxnBts4Dt0fJZuVEX8b+SdoOBxVWLnORkI2Bk/llrCPl+KY1Z/Tw
Y2up3JIYkJOmGFhgQPVdvT25xGhd3Ukr+C9XPN27lTR6STR4AuwTJcEoUkuWLqBX
81AjRdbAu6o/67Q3NNv7IZ6qUTM2lFoZD0EZfxUxsrCcmWet3aCHueGetheZp5C+
X8KBJuyJx+C2klQYxKlnb6uIwM7CpKrCd39Iub7DHvNBugJhs1r0745EEnS8fL31
HyvCKhDJ10NWL3t+7gcrO0IbAGoeOCgwHJOmMhLvrkUl0Db4SMKPruwylVt4f1Jo
idJ0xcjd5QmuH0ZOa/1V8A4Zuy26iZyz7VvkRE4D0opW3hugZCPAwAefn1736XjI
1Ee1IsmPHWpjG6webtrA7EwAYBW16owYO2DwC+PZhv0FoZmlMZFiT7YkOKD7uqtH
BuyKFxpyVzBq+kslTVrN7KjEGY0vkIFOJsC+Q7kf7A/fIs6oQryzjMkpayasVLHf
gj/Kz779rxPVt4+x5BRN9pL/HZ5n4zQNaU7W/ovW9zKIVhxKvoZzFcdSnf57ytdT
qcBDfleyJRFI8guYTjwp9hxmAxHmqMQTn02+8jw3SmGxV8XcTELz2/O6eeB0WxRR
1qAovkCQUmL0aaNLB407Ye0DPWphWhxfGQwNNhIuotLEhsuMbczpgTiKcQAfZjeX
Z+RCXXNVBUqCfLX/vQ+ZzPxoiDEWjtdoQMRlmE2RHhqul5eDjTMx7QlxxfDrUXgO
O1qsb+Pwr54c2POIAvfJbXHHnTtt4uBImJe68SuUedUE9ffH+aVqXl9lSVgDzYBN
aGvCL/MAelrovRxYYs3nZv8j4yCagWTbzg3FKGWjZenkEAD5epYINQB3KSrY9sLy
HPXmXsP7Oc8OWui6X1m9HOTuvKW/kYI2DbVsJVgGRtsNm0bKt3T9O9LF38epgnsf
N8cfcXZ480xUEJ9W/ltNVt32YrlahYYOOZYkVsdHZrYU8ynjQ+cVnG18DdXnLKjv
FblZ3CswLrVbDqwUm7H6RllXo/7GFfeffgSdvUidJq0IqXAPrmuwHCxu/5kr8iOJ
L5qEsfeAyakX3aX16p+AbhcCDMmb6szw6AseHuA0jdidwczosNL5ndUuczRSW/e0
CIS1LXYCRF9tR2zfuqodbQyDSd0dRh+FgKxZe0NvYlNHXqgzLkHCilwS+tixBjuJ
xsn2IqkilKv83mvhnbI6SDRJtXnF5nCzZ4UayQjN/JawG9fQx27FjTUisGpKUw7S
F0fePpIvS2wyMPNjXdwxP9Em+gNj+jJL60vc5LaFnq2i5QKZUf3ecVqSiMe7hiWV
y2QfFiQHpa3lrLFBBDcq6Yzyzm/EF/XNjvzDNcPdId7f5ZGdnCz49yeqvkIspHbv
8FEdNhz7raPd3oKw5r5rMjKdINsDRmSxice0w41/tTVLOfj26zBcA5BfPqllaQO1
BrXjFrqkWBkuVR57fChnoYdL3MhCJBBzI0/OUTGt7lpCInJnRCPgNEupPC8kyH75
KAu25Z64arFRgC7dvR3ZZvTobpL8SOgYxCPwedlv0atUylHCfJ00msxxUB2bX+V0
ytwawLtEA6ozXhEjEaEGKtcuZgCfzNQdrRRrOXYE9m9bGtklFjr1lf1pBGqpv1EY
h+7GTE6HaSYxRzakztX/0Ol+LEaQpqIaRocI8cIeS3vgmWfbjeZ7hOWqDztrI73j
Gh2p1VLGbNtGA+bSgQ5mkpXDJWZlKoapaTKeJYg2tQH8TnzBKFmHTPs8NmMiWUxm
UMynvWQu5wR68fIsEm4yOYDASm76zijeXOMc6I+yRrSoVCEIoliTkxksVA6zmRWv
sLVlqABJRS5jhop1YH8iesJupAoFgfa7Nv1M5td7w2pQiQMyV+IB2oIR0glSCJuB
A4Mbt8KBs1v72nGX/U7teQgyou+3zbttTVkRAKStpw5yXoBZDgHYrmsboUoACJBB
j3eUgIcglk//jVAawWgWDmcCtwrUetkXlgqNAPf+Te/aFJaeSElc7GSsKsyxclau
aQOw+OovlBpgxBDFcQej6cEhohuvEqMxw0c5dHqkYrstKuaXJAIlDWMzXMvwbRwB
WhaelXoEvFuB9jpUncBgCTyzx48U8toovzcCFyn1ANtYC5PeoXrKD1lPr9/RYNlJ
MI32OQISgNCZgZdIX68/wrzsL9yWn6ICfEtjfo3jzya0loNTTP6hu1ncXSvH//wj
7M2wz9fpAT08H9xKScdBK2RGXjjqOQgblsMTUfWnnlkGpKzekDP+AAvIdzgoktoE
hA/QcygV/mVhZUjBk8R3sUXvQX4eJY/NiGm5F5VuO95L/lu6cX519j23iRNyCzcS
URE57uSDqTJNi/RWpfVwoa6M35RjkG82E+dgYhTOKg7PxxBizIZA+HduD/uu+YUi
tL9yPoE32m6C0rVKOBssVWnQj5HatrvxDcjQBU6lcwzN3tBnj1KVXoQPnM1/5v48
zvu+TUQILQykBu3yHdhK3pv/8Y1+VcK48jCQYTv+oN8=
`pragma protect end_protected
