`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aAEqQsn8xpQLRyUEGfyNAec9DIud5DB9AM7fMZ/6Vd/5dkEdIewM7ZkyZVClKkur
TgDrNuv17qkvCEF+RCdwWdvllBGFFtizjLndt4d2BWB94eA29Xt/rH5PxCA8Lauv
7Q3dTjqnOHf3o+K89m2LQDPyAUAqoFGrkcKICsjS3cU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15600)
Eu54mp33kTRW766+Q2cxMCA++z8WxYR1dPZQoEhX3JItXJlqlNIDVP1cj6XCLGGz
ZvcQ/wXVideiwAVGU5hjUjW1gqeYULDPAK2xhQkmupycZom5l7/CkTVOtSaL5ubQ
Q4CG/qEROqZPRnhi3MxAnEGNRwdAf+dx6pRWYKIdaZJYKRiSVI+58Ul4CHcfKPzl
g6+woUINtCNRNw9hly/UsaCuY5+W/IFnxbANPNZiSWCpYSH3HoJ+GNBysV5VEV6i
6TymfTF7X9hFdpzHA+349ucZjEP7ql9JqyKuzME2/Y7zYSe9GyvKkdruqjQ/IgkH
gRFiPtNQOSKBzLRNHYvgKlRyhpIo8jj2tPVFf7ERyzEv999TqRc3kdFzXPDnArGs
t+TuiAGtRBJJsdNtM/pJCHloVNA1FQS2Snzd7vVPW7C3EYs2Pj9ZdJ0sEjQ97jqv
WWUUa7UntiinnsTGPUqAe3CkGmhn2YL1EDVThu4ig8g/0+ONP00mAYDn5uEVqvnX
DX0kk0tED9F3CLAcA1IQA/2UD6Dd8Ef6sbjXFFsesnp1hYNdk4WM274RYZBT5iB4
rEl7LjH+jMJeFPjqVdHc8XdX5PcFU+ht510i2ESl8C0/9wQx2MIZgJ0tsOYQRPlP
CuLINBH7A7Fe+jZzDsl65kQfl7akuJTbnW2cGQ/P0PaGbs/M80MOdxRjoft04kzh
gmYE9JTQ2JLTabYCVa8WRBbR32fiwwr1LEaIlHTPVxbhK79VGjAVLb0rsWjjl3rK
AJwBEnThlZ9nub2SwZl4R7ulQD34JvBKf/e978LOCqRLlTSRBaA5cFrDR71giwyG
ReVBXCSOrPODdHKPgJcfZErwUuN7XtaA/YlD2xhQoaldhIiv3YgTM7+BtEynT7n4
kw9bRNZf9HxsCvB+0Skz4TzZnjABx0JErYnnTiBpupVg9fAYV/lF7GJpxGB6C6pY
JXSNTjABQihDiLCyDpxI4HCWzoDk686zu7QuJ2L1IR2zRP0W6uhCMb68xkBI/oLY
2Ho4Lxypjy96RjE5NEo9znm1YjY0CqzcyAGwxPquIdHiXwTJBUPzVQAnGMdfznq7
Ra5B48IG13oGR/AN1OT/ODCsHlU1SfjyRyMiiKO3rC4yOLBYcrKAm9+fawBVIk1Z
OS0U3URWIlBWdlsAo0U1LkNphtuQa6v7kKHfBGJLXwqe6meu/3H0lkTpJEnLn6+A
xOXJ7MGwYsW2+kVIPeMDOyabIFDol69FbaGZP8Z7QpROomaDn00LiJVz4pZxZfdX
yD93zG6VWyc9Km5EhWekKZLLxwqDM6/O0vTIUXNXwgPe50TZtajxE8k7rAiemQzP
lgEZeSQNPi2TRo1lEndJvLnd95VF1/1M2O4gxrGsBnppSXdcY8z00nqq3Hv/W5on
Z+Q+kf+RX3VH9O8XNadurBbH297nwTqtr9oYtQYibZ6qhZTsp61a5e1G6AN82okL
5CtX+h/Jl2siou6umTsCJ/C06Sf1BhJMUB7DXCGwhkYbnAQBIa4Vmocl7nTQOywG
0R7VUmtN+8+fOJADyrVN77ahXFOtUFHEZqUrePnAznQFs7+0Obi5rE4cQfp+oJZS
xolnLaKpm11ODh+JKAqP6AFZPFUm76r1b99+k1DwUNN+vgi96YfFAJg8/MGh0zTX
1nvCk50oyrG7GWFZUQix7HHgywtXUOcNJFFo8OHUBfaRO6qpkmctjxBkVFlHOXk1
7d20n3gkfwqWI5nueQREOXPBfINuODejigv7uuKj0/UwdcVhxg3vUT+2e7a045nD
lzVfSrzRUg34xpGiChp+uqhGSu3O8YBmdojJw9sE0C71qBFWfq/naMSqhcxQmlQ5
5tk6nkaFx58JoK7d46yPPtmTeoRtUx4vubuog90APbxrXey3Bxdz78goIjXS73m7
oFF1n4q8g90Hc1WYtIoyRkFtBRZpP1j2qXyHJs3/SN4QuEqXmJDwz+3stHbOQKbP
zsOBWGJSXjUG39/BPCIfEG9sudCMVPHixKmW6/KuCarXdQpX0JGeeNHPVlbVeY5Z
5sXfTEbhzPx9Ek137CpwB0jj15nqxOUR/za0v/m5F5Yc1gPf+O1JA92ACOdBE38o
Q4orrROGNXFlDyIEyLnfmN+dQD32/SiskFVbUvSiGae7EMeNMapAIM9y6j91dgv3
PILvLOjZ3j4BdfjxSZY6bIf/Cc/XTV/SIXM9B4aaoL6TPOsTwFZErivZS3mqb9Vc
Uh/TzfRCgDPzRG5TTXo4YYjLYCPjY5oB5gEzvrsBLUqkzxCQELv9gOiLtmrCSJlG
caEedi9x2XseOSgsPuIObEokjTURJ8WLySL8e4hLZlAgmjiFau06dtveG1+AqQWb
MhQ9UDnkzcP5b4Nd2ZUMTiFaHUnfqkKLhsKpVVUvYOw0nvqXYT2GTBcMgszUFsRK
c9pafkC3yI/dguU7XPcoX48jSaeAbAcF4UqDVMPdNsWy+dwVTTw/uipkX6jxVqOQ
BgxFpPHcej91kiMSkVpQNQfUtoJtJd96Vt3koShEvkX5tqissuj/BqYAdOUmhkTU
sCqiZ2wHWUy4Ohi2mLQIFr/lQjf8JD3bCmzDgiApeHo36FsZiXVBTp8upebFzXBU
92YwnQBVb2TKuRUWwRQW8mj0eQmj4+DbSHDnoOhgya+o0S43X0QtsJhkqRmkAjdE
My+6o7AO/Y0YlRvirs4k5KtduEhJhpNjQbGtMk85DpB9RK5AnAe/HIeyEt4aP3FQ
i9ErfxP1cx4SFaqUogHdHhZ666ofeQnYwwJTwOvF5sFUL2qKj5rSHK+0odnFuMpR
+CdhJZUA6eY37HGPDq/WU0pXP7pi0N9q4lHcTuZlZXxfJG/EkqEWG/PHmb5nXUrt
SuVyqsowdqIpT2+ubpj9mg4mxudwk02QkzQ65mNEy3zfK3s6SPnSnNU1Wrjrcl2E
ThCC/exj7s8YBJUmFb63/Y0XNCNspAXhWwPkjzbdB5z1J0N5OV5u6XrBzVXuvFAx
3XtCMvv/8ynFOCpcmnQbPEB3PERylcPZL1ShvgVqt1cnroq8f2WgYKBsVZbCA49g
BH+xDGAbSZt0UWZcoPRV99WuWZ8iwtTgspNncHbqrnmAELU++Fy8meQO6cvjDUVk
5C2bLA+0Weu23rdzj3vZhZBfBwCCs/0BwRbx24fhJOzwcmnjnd+tlMACt+78iLRy
sSPpfdGtx124CkZcD6h+7IlOe1PN3wO7fb8sdIOpjVQ04U88gd6Ffrwc/XzKcHp6
Eqn4jvQiRFVDzcIXvmodZ1QkLYPzfzLe+lYOCMYy4UZwXPkbNi/0W7lafXhsTOVJ
OB8N2GevnmWI0t01gKmqNymGPtjajwg/7hXpR0X6sF7yV8UCWwZeeQ0VTOLuYk5z
AqI1auV5EZUQkN6agr1/UQrGLn+O3MGSikY3h+QD4+82BHvNOGVuPsGEUxK7G7tL
SOLG9eEn4hqvGXHcE01aL6PEUuJNhN6de8HufVVe5TVNe65kEE2oARvUTGrxa/QJ
004NXPfhPunukMulK5NYdQdv+5borPSTmdsEoTDigVfj4g7E7b4oFmVZptByIAfS
MCjs4mcKUNyT9d1j7+KrFjt3vTysZE4Xo+kXO2iuZ2Ltc1V5U4SNRnxFvhXwZJxp
WGXtsqF3wkbzhccR+EfRoUdaSo8UWAXBMXtCsTL4dnKDhTOtA3Zp8mHv5PAGtn7b
jA0VAMsW3mloq5tNzbUNplIALV0XyfOuE+tBlWTlAkxa30IQlnGOPXA8ORvFiysk
w4nJNWhH9nv+9JrlqDZZsGEtZrI/0PV0uqRdK4eMdeSgr1fQEflaSX9wuGwDCDkr
QU4JJQjXQI7S78XacjEoJOEEe/BGDzbcFj9FhPDCngfNrlIB93VT+X/E2LVwv8hk
WPylmEVHmq+c1qvQdSy4LW4xzOSg3FHs0+H3+bG0T8bl+490pel7TMF9EXgOJPsO
s/5eM4Os/4mOUhiLUSQOP0cYiAQc6B+ycS4F1z8PxwetdjoyUsK6ID5u5ni9QN+Z
4Pu075/basdTRCWPC4SlaU6/acdTiQHnzWwhnlojv3+bDjSSuVCEX2lm0graoxZ4
pu23fOoAauq5QR5T2n+baIYFW7Jau8iSnWdHiYVEjVfm/qPRvj/yXtDWl1lNu3KQ
CfH/vUivG/DLpGwZAugJyEjfO/+kSzR8DLSsn4jYNy8aXOZAOGisDGynZzHlabij
J6ejw3o6711o6rk5EDfX30ws2/wNf/v/ZPIHt5koGQUUBKXols2Xmvve9i5T1Fw7
UEd/fZPN2noDAnm0sh6zsTk0NpCZcdjJ3/8dldXr5fiLRCBu/QHyfmM+Zpv81+d9
SupkJmTLyaC2T1i0vycJZte7mttL2oEKwHY3ggKIiZ7/msdW9ju6tBmAedXe9Rff
eJywCJVrgBr7cNc01dVh6eOMzHeelwtdfLtKyMdWOSWgL9FxDbhWumbHTsdeahoh
CRi4TyfKaa/47t9h3CH3e6xjMGFGTMvw7qHZS81SliN02TSdscAat3mv7xkFSiXQ
uHJo8/+Ef54VHakHsR1m5k6VKcKLdYuy8ZxmfvUZywXRBf+U1nKlYZQeY6puNsSo
igrHEFAejvlKy6X/6A1gZ6ld9Vhd203mRiFF/DxCfbTlcK0z/UTOqIcu8qkz5whU
tPmVq6aeNU1TWH7oTpRQWNRC/cCZw0/33w4y/7kklJuG8cYGbAGAg+961KxWgn4T
HIqACmE3aSO6nb/Wx0exfpf+9qb1NDxdQHXFNHcnHkiLfRj8M8tYVJzJLOY5z3o5
amJ6+q1yvTaFQyPzs7sq44QFlTs6H7WgdN2SUjlxVE6PcJx8OT7CaZ2flrI8G9ie
ooGmbbDWsMEloBS/ETZq3z5egLrzGCndus7LvoFMyqZfGKVBqRLCRENhbFqfZteD
AeTDTU9xwRaz0NJeEOK2trT5gHcjgdlybTdk0QcFvjOPoGMlS/phAD6sXA3wj+U8
lPsMWCVZw033m1k/WHqiHFVnuEwKMWIuePaLT/51eWBUNMIIgBIXbh2Dbo76+iXB
DnT9HIM/pShgRidwq+LJ7Fm7QVEUJcuxk+vBroU0loavOAfgcn5UWL9ZyYdwXvHL
6e9rR1d4rfOWJh7atCtiZcoxEeklVHCUmfFFaxXF9esw/v4sbIkNTxQH7SWLSxEU
JSBS4H5DOWdBpgrEtEAM6GSMGMzrtrXztPwrEDbnEEoKOqbZSgzxJHrgc/mfHzOw
nl8hIqX1SznQdx+spfrlU9nMWbbvV6nJDL/FNcPH9ldgLtE85ugZVwIbnyUiF1Ga
Hs8rVHbAlibd/CJ91uW/Lis1B0nF/cw1BPPLBypyzjMDciNIuV9GadRudMkA0+Dt
rkHLf3LriaSNhkE7f+32qlpuJ435fw4V6aq8S3sIpJlmF87I9Nm8oFMvEWn1jqN2
HSTP4lDfffKUNlGcwKzD/wp3aya4n6tjPubD9rjBOJG8/jWyBOaWNEb7lrRRayHt
jsYGUInY/R6peMuG+O0w3nActYe9G0JroIddpn4uyiYsd6f+0F/ZadJ035a2rm7Q
XbwSr8rxVW7ghoy1gOXabIzqey8R2rd8SP/g8gNzxKMmYUhLfwazndgaYT6jMe1m
VWvD3iIjRZiNw4y6xTfM+MVkZ9lx8RtYLng2SdflaSlNcLEFdd6Qs2XRLFGxDBz4
BVF+cjl5DSffdPWyTL3srroVpivtLx0svvzj0laQtj0FtBPmv0AUq0Z5VyBN0ng5
etQEoleX2E4lsOaFWdlgHR+Dr5rQR+nmf3JqfSD9x/9C2Z0Ze95Ly9smwmGMsfaz
KLHLvF3brofwGd8kdTbS08W1n/dLsAkKVVdRfPnsJR9Tu9OEfMcoILUNRkAjF8PN
fkDNdL5HHu00ReyHGu08ennxkapZ2v6O2HCRpgCv3DjKyPDU86WJ5kXZtWxxITU4
J8D7zH+StuDeB6vgw5XcGnF3u75z/Orx76hTlF8WMXR8Iftda1iFMm+99mSKGWnR
HYAmG+Entg68gwYbHDresZWievfE4rih0dvaXshOosd2rCcJYRjLXMR5ELibvqta
4oIqEFEBB3l05YrbM5nmziK5gxLInmTrifJRWIk1r7MKWGdCCEtNV0T7gpg2Pps5
IHO8XLPO9PsyNVzzcRTdXLOeZykqBqpe/I4hWgIg9SLYS+HbbGxmDRV5IwiQxs+9
OAzQqxXV2n6aoEe8fkhLHx+lltx2V+sk5ajVWUmpLtCkuhlYu13FBrGyGL36Uo26
DNprRt9BKyD5NE0sPZYR/OB2TdgxQ+HM0eIHZ3VpDZI01GbHDMeNsp3tZ5REhjal
mZaIln8RUgUxmb8/f/E+P58emMNnF4ofcRq7FT02CBlRZXMmeiNt6ReQaDRNTOZH
NY1XMa0DEylyhXEZgjGIEuiM/Op05JLtIR/fQ/jD8LDI5boOZ/k/qfutz/sOi3fA
RB+Fb8E54LUcGpGDTjJV/fxe6rBb69xVHIB0SwhpqEjH5rmg8xjKg36c2CcR41Yh
hnenF+bI/ntV6Nl+dx2qePwgnxwW6IhWldnTF/73uzpBHt+LkKTWAcisFCThVEWk
YNV68W4m9ZtsSj13KrJJGJdptZ2sxH7AAkuxrJAhzer3zkikLLqceXIzBsfCHyFU
8n6j9lTv8w7v4tBX/Rur1qCows6ndVifUnSq364C3K2T4XSWEOdRELcKm7KL9zgn
kKm7ss6r62ImNdDKjVh4VJvQZy+1aQL7usD6CWbpWkJLAasLKemc0FdIr5nP9l4t
yB71n5yKeufLgExNRvqU0GtSsNgtvfAakBPFBoGKlGWTeNd011VKF5g/vlBfIdx2
jHd1lQEFHfKKJG5IuGVq++1RFX7aNOHFUw/1peWPPpfmCW5LAa2a+rwoL80YvqBT
YsJRMF76/VtRBA4GfoTaDIqY/whcruTBlZo+Nius07S08CFrl6ugQI4HBNTnaBgb
HrEJtmhJAnCKx2+nScaelTLMPkZnxRBDw24138vRKdyUNFQ5YQo2uRFEZFeV2UzV
xdcnIOedeyWt3OSdSNVeBPbCV+Fs9L9IGhZMsXUruW19U5EFvDOfbPjTYw3oKBWg
Gw+n9VV3xUlfXFnfyVKfOBMlXlDnBWqZm0wdfOduydchzAH2nFtefMhMDJiUvZ++
ibWM354W4OLFK4SQxihr9IKtJ3iyPZExLUBTiypyy4979y37jv9QHDQO1SZtwG4r
hiC6W7fOsA+pSlaM885Hjoz0R/LgODT7bdD7cufWreVmXPCEY+mKcAG/dAx4uovB
/jrTnxj1UzLk71dO6SHMJ//1SpeyMFxqjeOZPHLxchx1ahVcsa1iiJ9oSJODAJQK
taAvTl2dKBT5fTGvw/gqe8E0V4WeDHV3naQh7jMq049Hl8Nbzl0jFEEKqDhP9g35
XCtS5V2bWvMkv68tT1iX1ryygkMpDh1HGnsm5fhsYj1w8umpp+kE13qun1icnMRN
k5DEc3+UYMJ6163r8iiMclUl8Cpq0UpMzvELoqvzKrJAhALiUwAvxtV2rdhgLYyW
TWc03lA61eTWNPqar62vZn0fupg62mTH2IEFeasUkKxQK8OD2Rh1ilKLWngOL6Ds
R4O6BT1KO4J1zcegznxEY8EVP3k4nZcJttt7kxZ3oKW0GdQfST8IqBBnu9Btw+q4
EY8q7xfpQ7BmIljwi+rFZSCMb8PoTOFsR8DLvMi2XsGHijlj8qlZCP/51QNc/w87
OhEQ7Ey6IOvaRhCj9T2LzfJeM/kR2BqR+Lylh9t5LBxhcqOkfqP9XDcRVUfFscLe
E0iMIae04tmW1PyleZVQGVYlfbls5lx3saKTDZ4ovipG++jBCwBb5ILSHb4VK5ox
hdm6XE362BxsK4dw5t2xYktVcae6TOdewyCuj0DQIBMNw7blGNWGCScafFWdzTgD
dYeHUnJVMQiEkhILcpRXyuks4NCN3QMVKDJZ/aNCN13H6etqFXNhipC2g4yfvHiR
zeBixN7BYEqAWPnsYCkKJqYxlrxAZmecgzow4MEPYS2wUbMdYG9DNulgfpu6mhZd
ZJ7ghFGD4sqSFfXqK39HSIx/7iWijSt+NDmFo01MaXGmT6t+IWbYtaODmaKtk6/w
d0CH5Oi0ylhVtTQ5OyHdaPHf6HzKv2WzI1Xx8lFb2G+G2C5q7ZREgGj3r/CZ1+mr
QVCUy0XTqOn1Ap8miuGHy2DTbsQQpesxTjivE1LuZMSkyaS9M+rAMW4bONZJyb7E
TCOurEOX1LWGaAC7Fmavrme9lMBJDElXzgtAdWeZCnGXbgneAFBDpqN6fUNV4wg0
c42IqyfyWHSlVwhP4jTjot/djlnrs5j7BgaWmxlDTn9kTwEjWq+7vtsVrROlQfSo
E9dFEQbpUPrWXEyu2QlSY+mXNAf05rapFE9VFDkSwyl8aZFv9CRTHhXmMCkzHk2+
xbqjHwQoVl00G+hyFo4JlnQmaQQMA+yJ1RKe0pWMJgGhA5s8wO7Mc9ht7FWHkm2a
hfaouszO9fTzlh82YjSKFGf4MaiT2ro4tzumT1LWMFOXzSH/711MR/IGqhyekKqY
dLBXFLXEJX7o8MhPtmaQBq8XyXgM3x/kCSqLZDDxLRlJvmXA8SKg6ZVCxNBhXEVD
6j2TU7BQtMNHgEcImUJD+HAQ6C6lCVIGw2S45FNlupy/p6mrpfIzf1xY1wgZKTpq
XkgrrbJxDUtqiRdtW5+BBm4vJGkhfyNfftJ5Rp9xGRsCehamxkZXbel7dCQTsxiV
n4IEP+PuSqfNL1+MccKkLViK9RTurOUVm3pVjV3JZJWYdTC/EDeVQ1vaZRSKLWc7
7w4nkHpg+Ooa6mLkYMx48vpGt+DGAbICbD7aTpoYaKSppck8EMHnl3kxqm18/uRJ
4Gax2w+nE/6ffJFFfjiad9W1hCf5k3qxOtGzITE5K2REVI5+lNWnhr2qD7vEyH83
mpQCzzt1bRQ3rpSTCwiHYLDSwuBDrU3W3qnNc0fW0xD7ja6liy9Om0a7bZYIw0r1
UY/viA5UWwWJnm2JhPAPSeEhn4VNYsAhh+U7VXpeTOd9f+Gbr9VGZjWmp4L7dQ9i
gMu+5teioNqy4txbOijouWR4V6DzgnHowt0Ky7caSlFNM10w6cQpkLnflVafI5Jq
UicrxKmde5JA5KTIcHX1TXo0MZrh9X9cfehnlJxuSpiUyFJl9v+iv04EydUPjxDy
uvU4h9tTjt79Go/pDY158sSXW5fVetz7PH7+h8gJICcyq2Tw1Uydp2TiAEjYGy5M
bh9XC39zNfgdPYZ9o/SXdBmAKTXUjIRmEnKQt02xxaY8duhM2NOU9N1LI7B/6ROm
brHsZRfALKpjNGKwea+kMeX4tyrEB5s3rhPDy3FcrmpZwgIGPxTtJl6FVGrx5V3g
5mDFkxyE5xiif+gHJ3z8g6Iz8iJUtgtmFwxu6e7+U2zJi65Yqw1hqOoZImAdj79z
PeYXW3dKdYAPBtE3mbnv7NobCEFtiWvbvpMr1FxxG/0nuXSQwi8QlltLFEmaVdx6
uObM4CQx1sf2E8igxvf2XqM0hyESBb55qrGoS9ijJUzIQAsZc5jAqJjfzp4RQInu
uE5kxencAHBVa9l3ozqRJeeCi5M0GY6Wm/cdlGvTXP/PaDjC4qTokj+WQXh3o9Ca
CGYCMFd+gcZq1gDi8o7ro4J8h97Zu3Q88GC5oY9KUtGpqc6EBLZM+Fy5ctEy9XfZ
hO29ZCJXWpYzVOPvkKuV20P0vWcMybsdgmkH8j7sREhj3y2LTM51qG2rlQ7aZxo3
MzlBAR+X5o43ga8zBBeo0uglVz9uW84SX9uueLVm8y+7cNvcz5BUD0NrYMT9Bb7t
RKLwckDwIC6CEBRZLgYJxhXeraioLb92BQt1oTdun78P3inN6k61bim1Yyx4YKgr
Gra3pzt74DqPZkhqdHdEJifn/lbOom8Lq3+ifyTNWy36bP2j1qfMXtFAsQoqophP
0DuZ6QTyZ9tvNtcw8YcyRQZQ4yqslQYXmu1csGpJUIy0zonqUmDUE3+9VRhW8c3w
FNNnkfJvk2DZG07cpEje8MWX8qrmmCDkk7rkPYYpVKKMyJ84mfh3mlX6nF2awGSf
u0u7UoacIbnQiCi36b/RtasUqXS00Q8/RKx6opZud1Z5GD6S/DNU4Lih26hGbONa
HZBtzaW3vxX3D4m5S7I7iVyIQR4tmxdF7KSxFda0uNk13CG6+WnbFxyMeBNL44rH
EDLrsSC30q2tVDa4Wwhlb8anLiTD21kY7x+6IT3pya5QcVge2hNc4Kkedh0H7Ing
88xlIXDXjJTAerR3D5+EqvaK8/RehB+Hyvs9wSyPsBc2UXi2CM5sK8jsKeB4HzMn
zLI4IdEAQdHwgLUxxxIVKMqF4pNQRuJYBSCD/bV7edOvLGPu7bP6lxa9bO7WolML
xxhWI3oIdDarH5GrIoGsCLNeAC+zYbee6bPDTRGwvTUMZ7NOQsPvFouYACnEjj20
W+yH7vyttJUbEQeM5HrWtNa836kO5sO+Snss8yLmIGA8YdCYBazlhoMIe0MqozzM
+Ruhx1cXQzCy/6VtWauafCTWcf1h2zAAmOHsDAJwT42jFUZ/jDQJ7qcbWEtyoJ5B
0LMxoZAFOjdWr2Q5ApZ9pdFl3YWVHm0m6RQhACaEieVlO0RIWA976+KUV8O34fUF
b3+hNUxWU87nX/JcffUEivQpScF7JNVaiM/yqHXVISfggYaF0aG0NRdd/Uy/uqMH
FmH8K9RKHj/KFnicCAlfgMNgb+qjIHB5mSDNDEnd35UxU992mr9t2roGCbmACfPU
uLyChVfgpRTKtChbECx8aOeqe/9Di627TL4tA+mClIe+N4g522CAdCQTVBp0UrO7
y+JZEwMRl/3Cn2eIykgfgVbViyGZsNqEJpfH+lYWRzt/vXDXtyuGwly85MOclpkK
2sH2am+CqPxBt2agSMmK7nXIOGvOcQrLNe3/NOIPrPyHJsiCKKY+IVmJ3937jOlB
3pXAXbgG7oN/RmGIt6vJ5kOFyua205JBhXNGvYzibbsfnPv0Hnn9TwzcMzbzyh1v
ZSvlDDOKPeELPOypROTsjw8qyWeD+Nk+mZdlCSPbF9hvsoFfITqo4mcbkeG4oTOD
KUKhBoVCxNV+eY0HYYcKOyq2D5Y/WoUtJRa9owP0MZVERQyKWt/WSO/zn8zp2gpC
TqG/rjeGsx1PgFYzWGpHEjoaxBSeR5yv7ffK0DjJPP9V1+bqL2oJOj9VyT3RFhjC
e1XDXVZ3jq3/1V3n+AKtvasKueEP/LlxOo7j/VT1yHwhc0+W3DY0fIk6xw+rF0g2
m65UlvuCBaHq4QjLsx9dW+FRx+zSyWHf0MLyAqDPPGG39IrBN1w8+HQtN+RNPfqC
zEGI/xKor5IDXUsK9q4zRDmB8f2bE//2GRocyCF15eIPwO3X+PiTu7gy14Z+ybqX
AwBavwtIIABJwiJZqUGLd+JFsmFEn6McHw4oyp1AzJfE94R9l99IdGgzDOxtW6pS
qOav7e3fXrtINFoZNI6b3+EzLFMgw82snxH2twmnAf1kMCEJXy6fd6rwP0vcVf1v
7ogHcUA+bz+2Ohmvf4lrhT6H43cEC5rHFFUUIPK7eWKOHQ3YTAheiBzp9fnZMaT4
IhVK7a27WMuaIZNfZ1pUwhPDDHbWwJbU5nN5wFnqwv/Sx+sH1SuFMxp8hbuI7Z9y
G81bJHAVc+aqPZ1FEYc5TV4FL/6UQCuBD+hm9/vqaMw52lXlhxXrjb/tCMG4igeJ
ybo2HNcVKi7jmwMHpOFIZGf3uaKa8IlOhcDqSPrZPJUzZRomqxZrA0eGT6q0nLeO
Z8sQckRkdOGqRZ3Nh1uqG9W43Z+E2h5FCbEVj7pJYJ0czBQSH9T9riNESXJszCDc
/ssr5yQksdZP7pjfQ2hc5eR8LXrc4TEp+OPkuT5bGx7c1pvE9KRYlczLM+1F3L6+
1BIkGnFzJsqKuSwKPR51dB2wzb+qMjvGVvSb0ncMqVsvZuA7xL6pA5CLlQLuaMTQ
bJw5Sx3XzT9oIvplbXHFSW6qjW3gHs6sh/fKLc2yDrMfIbBRKDr5MTAwfvp47yNT
aHT3UxrAU70q1ZJ2YUIn+mjKqyLYyu8XVa9RmJUgsxpxLnC5haHtDeeMJvFGEMW5
Z5marHdacXrCOGtg5/xfGKySMOu++5WHgPDRf8cYZsOH6iYwzDaOqzwiD39rt0tm
U4S9KYHidmFID+azDD/FmebdN9dvpPTK7WXC+YNS6FyPxs2v1M9ghtWpDneU77Yi
HZf4z79CmYYOs8sRo7Z/Hk14c8lhRtA381hMoI2nwD6lUFDbJ5zp01yPBYWptVDc
FJvTLOYR1q9McXNCLEDFb8FIAxbsxidh5eKiU7bCPzHHdiYr7p+xCBlwumEmOWaK
SfetVj8ZVhmKgS3FAKPXCcIjZHNMnBHIICnHp0Ev5yEo4DoLfA7T/SQ/g1Znkylb
PSoxRh2LJSv2cKTl7Dqpg0h49dJ3EUptqyIiK0rYzcafYxBEUfCESnzSf+T9bk6B
oUzyRF9R3pTvUOpsAbZXvNJ5eRfYFJUNvSQj62Dn12XkOB4w6PSEblVPSEVumeyo
IoG4du65qxtETsKsgIf4mQt8HGN/WsagokOpJ9rdV7kSsiFLHeWOyrV9TER+8wIn
GT3k9Uteix/vuAhI1ezi6lh+3qvkZDPiAJB+2aMrpJ6N+4rY6xVojkaTzVem8pKO
jEWga+PEU+oEfR+ZwNKR7CYG5ekTiOjOb17B/juJ7YuWmDFsiAQB7ep3DGj/oNFT
ifCaQB7hWhTHgC1umtju574jrIdVTScRw8Iu89sjxbv8SgUMP2NZIoPmuHcnIado
rpHBxL0jfX3F8G+LN/oJ9qvhQXHXjCxsCRWSgP0ITweWbSSwWkjAMMAiKXFEkyS3
eXaQH/IfsQ2uuuc/PCC5qmZUIekYgCyhF1WXcejO7vA5vw+Ca/obueZiZ5hdtk0k
3KiN1TLpBLThMiWT30oVnQhNscJGGYKXn5wZDza5sbG0EQKyLZ+zW8iUPYqncV+B
icJIvKbb/Llu76Gjm8Nu61o8t7yxsDAlDALL6XOQLZIIBD8pCYoINmn2fd7/Tkbs
6+1vOqZgpcHm5BHB9Flhad8qQA5KRbIj5NXgBf74RFal+O1UCkErUdFDJ28ykjA6
p2BkP4w+RivD0KYbonF4wd3YVjlbzi9DH1YdqQvU52P0pSTXJsGHhhnF3o7ZbUyA
dYjeU5aOOyiIhfjSMpB0NCYZS18xiuAObibj/5E2YwMI/IpRO+SWEtipMZK6/rdW
KwnHljJDINRfbuL5vIoaCspWKNt0c12uNeqM7Nv662U3w6+PqzoZhOHX+V+Ut9oF
zqVeFqmfSyBtsn8k5p9MYU1XaO2ylUYaPRxJr7FozzpuJD337mx4zZwXMPWQySv+
C1c7X7A3p4NBOJtYvSsuPrD+I1WX/fSqAHnEH6Y8bCrcS5px/fshsG+f+iLr00Gh
0VPL5+6M/vPtUbsUrPNfkWIo5ydsUvj8dFC3kP8DU7+B1U6fpmUbo0AXUFzvM/uf
VKYugN/37RvSscazo8OmxBudExVoWI2Pw0iFs3VSci2TCYvYKhyYvNQkKdCuo5Gr
+I/VoxUNaOoLd9H3R9x6ad6LTtNOo8DNN5ZjM2+MO9Id6zH2YGYGhaTw084Y8Upn
zBlyZahQy2RA9nAtVWZ7gySVQmwoyuddPewudyBTJd/jJQ7hmegEXlmQuRyIL6QU
Vb/PM3hmvzAFwTHf6MA2kpiwaLnG2Rhtq9VnOKMi/6NCk3c7EClWNaUhfYrqAtA+
hxCkHPrj4h2B33Lkd50uRx6Eu0+9bJp6bWe3pS5WOGX8nH8HnVBYudnThqP3fxie
MhI5Bp/FwM6JOYhWkEbW1QlIzC6BylYx1iIKWSFIrYH0r9eXucpfWA0ePgip+2Hv
MyKSX8W6JUAWRZO2k9V3dWO/jpXBWuWZoseWNg1cq8CNH7kkmD8tIYJRINJE/pbR
aOyKP0gByfs4DIjPlV7ogthTEAtsDBosHvLvwPbMZMLJf5/bNiH2XBtfuP4aQYwu
YzuB6ouuO18a3JDVN5E/om00rXkqezzEN3uaBG3VSms5rDEbMbbsqWp+iBE3Fzi9
TDnBpTJ9jx65oQxCI/rq4l3zmiS4gwtRbfbTXZJPvlJRAS9/Oyws4Rmhu3Svqwbb
T3RNnO4qIf3wJTUz60PisUtnkAHqOa5vgnyPeUJEushXE2OFYdaDrPcp+4wmAmh1
zz0DOz6pbORtMifTyAGTDUJn2uVBq2AZfsG49Yz0Wm1ujVOh/LmGZmnhFtHYn/zD
A6MH6nV2GH/peqLQO3oezE4vXV8qdKYNRSRup8jlry3plQJejVzXFy2p6ccTal6S
Kog7NMiTmhAPIlJ2fami7SQ6Y3hYEHBhs3XaUTjCgLOMDsjNZRQjtak6Ue2a9EER
5BJJBDZhpBrPjZHpdj7t20/330mniETJaKSL9W7mH7xDwOTjCxIor9jTzfq/sT/N
xP4uwFoum7bfhDM3p9nfj3n8ADDB7DXAM5skAEWNrRiQx8/VS/uXDe1omMB75214
4YijCtX+vIbbTxm5TPDhZi5mNxksj/Og4dc0pEUrPSwTjE608SmmweFTWEKpYyYQ
e6GbUpbSixe7VpsFWRRFu9RFkJgR3sM8rYZvdnNzfZJTZG92DXN11ormdTcOvvun
DCExk4jexf44YA6Duh/3ztSyo9pWkFvPxAajNtZwjcuFHnCRB9197SDigrPOx9/V
1yQJ7i5f5vmv/fcvnVD8mnZ3Ne93t/u8sdUpxgSHOF1k3AuXY+sLOafuPVRN3Aj3
f8koCT+PNeta85ZSTiUcZferWI7XBkLa6AQAI6qAFsG3DqDr55T0AVwqSzQgWlUW
AEqHCC1GIMr6wL4JqAClEHKCrFwrZfmKXvEiVyczKA70ces5orOWhSlntByfM548
FUsKWXBul50EVFas4hdfAL8jEnq0To9G61Xu2mpdMvs7trIMeFJl3gqPL00+kfZU
8lLtYA0hR2ZyVswlDbDqL78PQJMuo8b1cqb2Ku4Suj2/fZ7PbBHMkpVdjoVpEcC2
fsfbwv5nHO2mQ6hN/YkXSyh2k55tNd3skc0/iJZzGXQUXE+tuQOvIV0RJgYTdRvs
7riEroJ+D5vrqAGkAeoWmWL6eaJQIV8fjJLpjhmCa8v17v7B0ILnDX+60OMvqovw
LrUSSp01+22URDh+DwfwJ4mewTsp6XvOFZPB8x68J5f+c4hIhgQdzxbf5pbhYsKE
Ypqkkny4B5K+Lgc5/mmyTh+RIbMXJMuNMfSvt75T+CGtXpyt53t8IeW+edaX6xza
OqWEcvLFiAiMGHjD03xVm0CIUf2SlRZnk/k8wxFXZozFnrOLPdgFm0MFQJa1AYqE
SNlwaNkOY9wXDDaNjxslC/mELNPsQYHZarNE+C/AvIMPNdfwVKc+6xEXAN0tKTmr
MfoAUj2ZO089Dsq1Z5E/DvWDTpF8BJC1nbdYd9VPHBc1v3ejaAFsgJKP/798hBcT
Fe7yZkS3jt8jtBKe8wzDs6J/Yg4705n7/2nnAzaIeoO31g6I69mlQDPlTaN2bCFA
0lu1LBwnuVWz496dU8I1rv5Qa2m/fQn/IiueWZ8/KRvb2jEprtwzTiK16V4FBZiH
FleH4mynVoyd2eKMWxyaZmib68wWb/m8p2KEXovD3qKOsD42vxZqfa3LtaeVPyos
V6UA3YCF0w3+J1YXC8wu3M1d75KXQ45vYFnBQzZiXW3cuWvSwbmCYJH3FdoIvj02
dHpjowZH48/jYgZT35Sps3w4SMSRhB1qUj5MUpEosChZO7a1lQFSfgMkircVkCx1
98YGErD5opgALpA6psfVtUhwiUCYourOVE0VZDHLP4HXau3AJ6SV2iO+S3KMRflY
Qp39GTS78dG9+WpalX7RpPcBV7XqfnfxJRWL+MbjXSfmyiAtqgtAqKd35OBnadkf
tYKm+QbH/8cnbOm/v2feRALV/4UPLg923a//WehT+ee9dbdn5SwauX5JWL8hHZk3
jhFlMzCGCeXGQXJ1guLlEZ7YYMtOyVKa1rrdRjx0BM+fJQjBw+SpTlEefm9bCSjM
0rTKRkudQprDbXfa0xhaHghQGh6SkDPHJpLp9lkY+lzvCTCHlI3cOl31HVF40LHw
EuRnKA7RZNIpHulufDE4GJYbJ7Wx/r0/a/2/6V7kSap58fTDCKGgjhP+tRiFGF6N
sX7EouSFwrpnpln4/Wp/YV4+LeAjkuWGRCSuZnxA4GiYBJiNHlDa53Jh/+X8YhNF
ihyW1RKrcU3LsTrBy1gpGZRq1vuxmPF1M8qEYqB747upOu4L/fZeqeX8s0PMgdkv
0/BXrjjOgIzKTIG/BW0ChS2Gcv4/big+lBV/7xuQE6mVmBACrWHVHn6Iz2aSk9YQ
3NcL8www+u8m+BZauJbNanNMzpf7NjKh/WZLIj7I3is6kB2po5EljUKG6RCKsLFD
CwiDt1y7SY76M2DVP8cShjV5321xiHi9rQAWDTl126GRCl/4o2dEr1FdTU+GyMjw
qDOapSl2E1w+rTQzxObb7YY0FHYdHSG1AGVS2ZNQRdFcGjGY7EecRDWzcfOs3SQG
LMR0Dy5oSKV5EBkns712rJMD6DEE5QtS1/YT4xVt46AvwOga9o/hu2skgMlkR4cu
QUnET20gm/n/gPa7Vd6uM8wKWv2qkST3eRjEU0N3tvEVmnT/suj0xtqkzGLd8VIo
DU3cS/mvWOeUY4YNiEMV43cfLG2T3vxAp9jPo7XED0JGy9iZ47+PIX1DIy1ZITz7
IVZyY6zpE5MLAWM8tQvdDi7Gry63tmabB15M+7S/3VOdBIWXVxt458D7b5/XmoF8
WwJlgu8TuD85l0Rorbaw32WkvB3o/ju+5FweCqFqgFKA8c3psNMSPy1BofQlBNQK
+lRMElDF0En4B0kmnSvl5VJZiFth9Z9z0LCjTq6u1AxIkRScby93SayNc0mmhVg2
rdwcMFOS+BacnYy+HeYnBqyVcn677dKxGuL7+sRWdFJ8i3Yzzhfad6L1WZsTOwET
k4+HjiU+b8SU1IQzQREADvbsTm3zVrlLpGXs9WGFsW7AUKatH1gKjbax+IQtTTgc
vPs/UkwAXEDgL/SEaiHy8hpRz8laYeyxz7hRhw7Hg6F5c5xl7laWKqTEdwSIbjSl
6EKSQF4VxbK/vX3iQKlyPOpYnG0Xg5+4ys91gSTBAQT4V7aSfM2Hf40e73qpwRXr
8+iMrPidWE10n8JppPuQ/0yoDF67FP+baM/bvpi1VKmQF7+JzTQS4ZeEhve+QnmL
Q8NHxp4P6Ghgpq2Wvd/gm9VgDRjkzHQRpKL8UnSOmpN6RrYiub9n4Chz0Sbys9vu
AP1+dIJeRmdAbzGBC4E2k1hLRQacNTFsTh2iZNYylnSmplzmCamq4xLSfXzcybZu
0nKeCrvGCX/3s37eyeGgJYo7qH8jT9fZS0gdH8IWuYj923dWp4oA/uXk7H+d+Xhk
W2+ewnpdyfbPuCjCORGoO8fD/F9fal9Ktz2vNb7qfy/9PQCUFLXN26Oy7i22cX88
eFP2qk6Q+JkzLK00NWVhpWpIuI7EaEW0Y7i2l2PbDYnLPVj1Q59MKxc+uCyjgTH6
jvO8IlEZA8TkLhxcbUCTTMPw6u9CVq6Iwry02mkGp2lSCHcQ90ZAzJZWtDpkjmVO
cCKegspHpTkHDQG8yqU68uR6wIadwzh/DZne6sbaQ8f7J3d/lx2oJnsF+VhKSBgC
/03IZjvS6qxtVM8tI25mMXqcRRZNTEnRscR52qZNpAx0mBvh3Q9nKJl+977bPkuM
4v/TW3jVfLY7aLsxz1i6j0U53v42sKUe8pPK/BtvIUFGhQ3+G2PdnEPPve2xA+B6
NqLGR3G7C0DiAeZOoR3k9JJuHqlDfmPwbaw1q8N96Mu/NEDZ1udtuHtBatkK/kSC
STN5H3RLadyXVCt8iBsRoGfqwzfpNpcKhdeE+s9vRXjw4wZjSlTUTY1z69axnEcH
znmOPZj/2Mg0DbG/MbB12J/IhHNX9MCR1ducYb56mj0XsJaMo5OezB8YTNPijfQD
NapgtUk8KHKZDEBbZUlAYKTKzqQcXmdsrxhqxo9bsOUn6gxXo3zkw3BZYb2P7D5n
juvxrHXBHN9FOVqjcIzbcDCn5n40twbx8XgABf2fpegGY4B/LwGK6h4sq4rsgpy4
rDbW2Vbb7MN2cGmDhIBcVp2b/IC2kdyptOmzdZpRAB7kLsB6PrLpo84iqlz5qZXn
RYJAknO2vwkEbshd2c4pPE5RZkymR1wfCNL3CywTEkX8HPpiIl6YEKu6IskViw7+
HXsitUgswF+JQpmCNZnvaDeO44IGXbo12a69snRVF4T6PEzOLbHbh41jyYV8L5sp
SqfdbqYMlQ9DK8GFalkTHVnGMTmWn3GeeR3eWG87ucXckzJOOe6SGKsqCS/8b6Ne
lA8FTCdTABqUp4f2wihJ3H+AnAGl/Ncahl/mpWjjZJcequ0CCbc10F1Min3JYwaT
wnGT2jDnoJ5Vry/OrJOp9B4XBozdNKS8RnY4X6NNQWpwvqPx/pZqysunS1qFXPet
Mgji/ibOZKPJg7CxnxW0ls76XfWL3ke4/R31yl4SooLzE4+OSbXgHqcdalx+LWz/
rrZxYJSPM9qUs8aZuGLQHfIeDmeeJRCD5UuFAav2tL+evjhhlRKwAKB1Dm4L8/Q3
Q/kYLVuAOxx8Y4AjxsJZ1jW8pX5npOmrF1NtqTpBGy3cDItTdHigEzHARcJuscN3
QjKNFtGMM/wWySloI4bz1i0P5qFEYlljq7GLFiloYQirwqCUQS6qPkGDL1cvJKfc
3KbeaK0qrwuIllcwhbt3P4QnRZR2Egk4EJVE9rNJeLOlndRpRXXKK5jeY98W69a+
K3pmQWubz8nlCbUlaQl7qUsZrG2N94D+rxDsPKC9Te0blg5PhJFJjfQjgs4PY78+
o4dgNIgtLG6vd604Jlk1xgOIgD/vLGqGu+MND0vLzZb52aswv9FubSv5zESRZ4kj
TxgfM7OEwNzYB/iOAHhm1MRWLwrrI9ocZWpF04N9PC7VUDEeE/AT1lbMjDrsWRRu
SWjMWtD602RzV243SgfmbDsgHt782ZHOaQTBVswPFo4X4FMkdg7p1kO4uqzdVdEI
Gv1Lcumi3Ca6RYMi5iVu4YNtsGOGbBvfb//6K19b0Mj1quhtcqhAHK4BGpC9Woq5
HuOpyhHbzudMSGVJQIDN+mu4+KURiXVAvu+Q5kbdoTrYWVEyIgp5tucsyGDTWmcG
urmIJqBh40bmKz0WUs814jsCa7U5BE9ffQ7iVj6fCo+Oz7fARhfX7qqhC5nW5wdt
hODhV7BZHIRFdA7e+NzfuUf3JdiYRhHpjm4gBV7jEFFEJ/Lluz3304ZF4PPIUv/u
fh2Itn6xIhlgWB1OcFfNkNQsMBD0JJ/a5LbNca1RAdAo8qFevjbzFVERmJbZhlh8
fbmzLpxg6nJ0fp+hEz0oM78qwTN/V/tRubP6UlWXL3JNgXDE7KaF6+YW1r3r0teM
6jmhYMdPHOuqX0RUiKc00KTLp7uOA+YoqNdSLD8owAROupm0xkdDor3diA1IRC7e
C955IuZi1mhD9IbOqSBDhFBGmVhcgBjp43jSVPRjqaiwlrI9dUMa3bB5v3wOxVOz
2jACAP1laeVeWCuy99BilzHH3LE2sFXV9IdAQ2FHvjwoeiwHmnRktnEAKSwIlopq
dBgipWrTAONYYAUwyV4OLqwVbr2lRpuDMPoPBo7Z1wbsrWNRMwE4oP1O6a66a1Yf
W5rIt/ZilKoln71L+s5kkTCapZ55QVbTmeqbovN905uX6QQ/6Wc7IXeFHSRDGAXK
2ynC7+9vrGX11RO0eaeWF5aUNjavNFp1at80RH8NfFUgvtBLyNSIjRgmvvoiTRVH
JWy5FwiIuQ0yqYkXn7X237/FgMUHI2HaRhUs7WFaA2XvNIJb+HpfeDazqiWGGL5W
Lfn5LmCvZIZhcgs4JAF1l3EEU5++DB9SsVchVEuOGy2Sw479hMD7RGeAI4jCO6rE
YYoDLSsBZlMqEj5igDNeM4li37W4inusAPn526YhDjjVt0T0uaQ0h/Vi5xx4pwTO
BDJWpBHumb8SKParMK4wqcoUpymSCuAYdcEv3QIB260Zx8+VJPnm/Q/bn7LflVKn
YCqkopH9oDDtYkK3J5Fk9YctgLvQsjQ979MgUzXszI00NTwx1AOqzn83xtKK/2Jk
mt5hY6wAk6uTC2WdKYcDWpXKkCl6WMdUbWaIbNN6JOb8iti+4pKR9/CIsXeHchpX
Vl5VLQhvvAEhVxIG2u9Ga/FknMIqI/fMUish5IWI2gkyJVXsSG1okMRur3kpHwcA
x+ijgauCgEPbNIus/BZeJK3dXdbj6DIyrFsWZ5wM2cKcdnkeF17oH6AMUMO/einU
nyOQ8WWnJtrTbjKadYX7ucjLaFPuEsnaQXGXeun9jLZ/cta6sXlGg6uTJxUyyHLa
LmBDXA+zLWP81/Ax0sQwx388iJQocZRI07vn0t2C5/WN/KoM8wmaT8pOPCQ4iMna
sUqCXHoEboTm0EyESnNYNevwhdFKB0kBAGCcGFwmLv46+a+JkLRPPrOT4lKDIqUj
MP06Yu8lPp2HcIsycfCwNyV85Cr5dfqMRxlZCsPZCHOyQM6HXG2UqGTzjZOOtLtr
vKrau265hKlI0UVGYoaCea3qsReRb0kyY3ezave95MXaQqTcRGpLTHrLxmL4lfE+
`pragma protect end_protected
