`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NjSWDfEZ7CMCM0JEVKFsdN5tqF+vJkfFaE9XQh7GuqFTkPBLHkJVrVEUg2jcZivt
fG7GyphPz8W1ThWd3MXTLtETurKgumeGCFb15GZs7ClDf0LV+YL7wPceDafP/1GZ
Oa2rUAe9OJdqrIKbWwIXIAvYQc7eTkrr8syuudsw+Y4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8960)
xaeygDI6v9m1iySvMNyKcR/aEED9UlZtnZUeyxivFMrtfwEIlU3ayPgVaRTCzuvt
HmdZGgE3+FbsGXy2DV8HPUUPlNRz2R/weUXSPHg/ZgEn/zl2/IAQ9RYdVNJ5ga5v
0MZqhBPl3bi4bdWBZv68qXq2fs+UYaiT8tskCx3TtDyHOZIEA5HlEKEFgwZOj2+/
O1cXlfu/ht5bEo5yBEyWIyajffAPMgqphNNlBuDx71hqQXQvbssI4wcVgh2cgCs+
xLjyl2AazS12JY0STu/jfSDLEUgSHqy5t/FzF84lKyNAv0FIt8C5Nox8TmG1i9HC
uDSjbK8+nZN9C4RBSKXHwygrRptN4SEpv9NBK6Gf+vTbdLLA0zMae9WEuHer8wh+
HUEgf2gyo373rAfSvomFcHn0QRtSEO/vOZsVGKK1thY6X3yO/ly4M+G7m9dpwOlT
twFLjig9cjuaACqbyFpf3jSb6LrUpUXQL6qsrI+Fii1qrVaQhUAfL8STpHJZb5IF
Wude0ZGRCMYRc8N1o9DNFihbS4oRIC/6R+le+VXC+O27tmVs/hL0C4kpn6YTSceO
u/5CM1j3DHEm9qT21xbDIsUG3jCPbokyUX6leCdKQTj4HBmst2/gsxPbyfuVo/AA
RmqQHbUCJOQt4qnAdmEnRtKIdJFJscsTy0+3+wZWkPytwZuP8WwVf9h+ooPP4bkG
123WTYNiMAV/8HLna3SkmOfUQLthgkPVMYiDGteMePvnrR+jr0G4IzqnCKgKJOZo
GJorhHxswRd2fGoGP84H091lj1KqlIS1EkulGGfRpw1/YkIcuOjae1V/QMgR2bzn
ba4qVeOnfUYzvOnnFOYlvKxphsSrzWnxlf8RvIGMYFUClbvojPKQd/2sC45tX1Un
lcEFJ6WGSmv2AdRRqhtf2THICWxcZZ4dOVvE9ePaESdJ8SeleuggCb3y3ajPz9ax
GNNBtaCD2GA7S307AEAC1RvhUV1XhyNquEqVs4I+CeQ8GNGUu/jpPoNX2IDe8c3F
NCBCdQp7OcK1f4AlWdb8lLvCkJKmiIE6kUFgsnVoZC6cujOZymHvf8wBafcpMsPO
HbSCkxvPsXpivJmptRcG3hQyI7lT/lzMYPFyk/k2W8Cv3pWMZoWhwIRV9jzEOzcR
VwtfQzFgxeduJMz1qwCO83CQYn1D55uad7vo0u5gaFs9e1j1tl25MMEyedR4vu+O
nB4SrO2/nGHjxPf6n+V4zXIO/bSo7CKR3bXjYIzQwRoGivxHJVLHjHf8LYWNKuaP
Nk6VG1W/OXIUvihzIZ/dsFJjMrZypmoMPJDAAtSHkgV22Y0MeVfxFNY+ab40iQ3t
gaOy2ss4kDJVpQrEyRSdR99gKJOiSdFoSLRLR0/ibvaAb6jSAvUAJNnSGirV094U
3ID71qh4ODbTZQUjsc0zk0M0hyLXJSKEG7/rPx+RIn8ILt+iRSUEhqH7zOZqs/+z
VDX19zQ+DjgmNFVpLpaphoYLopAqw4/Sm65jIcCtCl22YaYbrg6TP+wA5hyysMwG
GcCyknIzs6QCV2+/7qwukIni6UktVLjdOOe3+0IzBKwWww3rdZhvSgo/roG0f8BF
XR5lZTopBbWQPpvNRLQnkG1C83L1uxhWMvOwZbDopKw5VMjZYACsJxLLfYDMS/ik
H2BSqPTyO0/dyjg4Tr/jDSJYTy5H7nK/Mkn3+tnl4xYHfa1B/+zityfdesuFyqAT
zQ3xTeOcdVe+TVH/XgJexcrhMRi/u7cy7bT5xjBvTbUQ4qThw/aFbOQjU35LH8C+
7Yf1VJ4PCUwIq+VC7O6i4cswZpC9qBWZX/hmB0r17LJbzPVh4bTJ3m04uSO5SWY2
390jnidFhIKl6VnU2tgAs8dFbgvqUkauPKIyXXpX6iZFgP0DCDNGgjYh3y3yY49P
+NFbQ4IkGa1GHtuWXqnYBmLUIVreRarVvoCnsT7e+z+0gw+yXgsxLrD734ITETZh
NFraGVzUr7dxEW35nnTIVOBjRXgdStsKbT9d4nvHjep0ZPty514FCzvVfXjOvmFr
EVxdiry+/2y6HdywqgCzUeK0ZxCRDEieIpPOtecY3PSlbOWigiXZTOgUYCJMrxVy
zFpgDXlNxl3SJOAYsGgdwMgX729Ybb3/+U80CwF1CI8wkSodZnZqwJHCjvdbi+HB
SMFj19vuQI1meLsgGsjvzji079x/yXzG2YOSFCYCTwyl3pXt2Ao2rBinGXObjuIk
sraMDPQQC0RyplHx5SDc0XaAG+ZX52aPiAg+yMTz2GpoxDYJ6B5DO9ybwakaLGMW
A4kexbcRhGnWtZXv2ELHI8Hat7r/wbzEFu7AYDlfytYEDYCCWnpxoRdDz3sxQ0Wp
f+fWditIuuqMYQqo2u1fj1cJyS3CeFboE0M1LJUCnREd00ern8ZHVfAbVrXF7KMG
qwME+cn6qpTcorBcs7l1SQLHLAP3nX7QrO3wLlRIS4ZCnroIr25jW43/Hn+cgXqV
yS297YBdgfJMs0YrzlYPvLgZcnhI3bpJktSdQD47zK29DvgOuH7nWSxDs+UIdpyu
hTbyFlprEvCoKbm7c25OL2QbLk0ZNvDu4xKw2gd0m9MeULiYy9cxv8urABE+x9a0
wGB9aS13uRoqyO6159HgmbOw744f0Q+WB9AkC0scK/S1GqwS6yluQyOXIKKL8WOa
JNNSyBYeIQpG8fsq9UIuOUjmxFdXS88wh2snKCqHlRraRRApnHDYs2CsgUkHtSmU
LeUQ2jsEeudcyA4WeXC3RD586EmtnRKoLGVAE4FMwWcnzcisBCgLIAsnkSc0e3St
n+jyOZSvrXjyLNnKtamspiJHHpLnX5Ibd547wy0yGqFh5P/X45xLa6aI/yOpYiKD
iMcu4/cL8ZGNGwojY+TUaUUBfg6kE9aFRH8amnDbyI+LlGoYVkmexd89NZXFS62b
Z7a6cW56yUIC2ZAv3IW+5ZMd3Q7XxFj4peZgeWw4NRJd+R3B0kc8B04/zbHpZAUU
h230UOMpRJ2TekveXyYleapsEp3keAIxlEkw8sxvBeOc2J5g23aUMe2z9y0mYcZr
nXyDvbCOlW5qilK6IsagQpzQsxkgClzUK5GO35kTQcxwJ4iQybrcM6jJBZt+eoYD
5bPeCpG4PRB444AdCeltxxls9f9FMBkqyv5FoyLGEpUOnRCYsfeeH7gqZg4ToWYx
wRnlqxs0xdV6VjGTB4lsmRN6k07LUcibTcXmtX7Kxdf6NbMtnM4sK0I+lSyc2j/C
6NHg4ycU+A7MqkgkcXCBoEzQAOiGtXIFYSsNydR5wygdjB+xJXzgh+xZnOJNlP+b
hFBA1rNLRu2/rRfIxM5CgJv56G3ewSm1WPJk+O3xv2xyssazNmrs2UMjcQTOy+c7
jcaQswvJHpO60upIcW1t0nw6StQgHmbG1owjy5HL2D9qPZJrrxX5XpnXEu+a9o1b
TY5g4J8AZc0eS52fUz+XtjqzotGDkXfwdxqwiswKRdssKd4vJPHTTA6EwnqXcL6e
X0vcJEbtKHg96IqdiN/f77L3cAT2CrrtPsn93u/Z2kFwNYha9KNMbUNYbVfwZ3SY
OLdIK2DYzkMqR4sziHRdoWFttqdOrIWjJLGlMDLA3o5xoNyTmQODd9jvMvjuwtxI
k9CgJ3VWbCabk1eKpPXOWnKtvxo7BX415U5WKVCVTA+saIUc2R8Ulr5nFnoNUiFZ
Gry+cnQqjyifE3K5dRbHG/9u/eYsDl+KYEFV+LeDNWOg3C6HrihYFuoiolJguaHd
ze38g4p2i9N/yqwdHUDw8tla6iPG6eZgK+RIYa3Niqq8a3BVS7MAM9zy2tg2Yx8X
d+yJS0t2QXsygBydbX4cEsYe3jgUlF/sVA0t9+pIuaKEa4jPROrhg+EVxdWZQxxH
7mv61MsHyp0YOIXSDxQX+9e9cC4hH9t20i9RGvpuApvORz8lMEwLYpNOBFDiVge6
xGjxV9+BdQEwGm2F+r4jWXG1OxDr8su89WOLcG2YhzOjHcO2+vYjkgRBIJVn8wy6
NgfAYx1L0Q8ggbPzfA1L9ALOPOBUzGmTniDCP7lSHrUAUqJtBiSCA5uNzxydQ6y8
QsbxAwolZVaCSmu2PRzRduuAr2nDuUYj8YehJBCiXT9Iy2kdm/IWfPRtXw6IdXxK
WNmYeQqTSaHUbOiYEnHNwxQ27HrP/22euYtDdn0tmaxzDmj9C2j/5xhoioiWxtpl
m8d2lMT4NBmFT6sKapS7FO0d3180eAkkkv+UWgyCFcGL/HvOSDRdWHRcZj7/mpMN
Lhnoz97MqeR8XQ7jHoR6HckFNvE2aJRahFbBakeDEklGGnCYOcbq9NHYoVa25CI/
920mR37/AeQBloMy1ueZ96V3Wyf8flKjo7f+0Jc8GugabCA8uxHtqvHHaBZMCwf2
59ZwvX70dzP8EDkG7DDayKyzQtOunrL/ud3p8DR1zDs/UPN7u2ro4NC8xonBZz9+
QgWIz3k9ls6XNvEczdWT81/ESOH797Zk/Cz/NkLdSreya3BVaW6Pe5pF2/tliO8a
20quu+B/BYV+ivo6PkUip0+yicptxyE3zpd3kJ3WcLRU8lzK/DdMkPnL+78qRN/c
5UnjGWLBxNL4wFgHSDuxM+jXxzVualKB6t1YPOcCwuV4EBGLYpeO+lJ+mpNeXTWd
49EtkyK18TlQLcGXgwPcXgfmfNTYE/esTpzdi3+BT6BY9lCg5BZytWQubZ5f0d3O
eyOLUpVkhi6q3ok1UfYc4iACAcm+q9Ulhrr8+2r1ZBuFwo8xo4xjM0wT+rHawkld
VMSUxTAHo8ouruyukFFumrTeu4fnkisxn/qN9OqjSKamX2QhNnlfR6k+APfwdULb
jmHg56sxt2jaUI4VTqbV/vXErXdyyawZpHz690+vd+HjXBKEpkuJTxsUrGWTU7I+
ORXJio9OTgNGwfJWDl4p2q8+mrEkFSTIAblIBMvOS3ZRnMIjo8MntQJa5HBP6Fx2
BfjoFkZSYW/5oRZXeoD2wvfdVnZVqkRGGo17lFtINZ3yySPjAtTa8uasTkHbHWH+
vFtGYDRKVglbvI9xBLOzFHVC1VPPSQWv9Z2C/rDp90HKJOmyDV2B3etBSJ84VJWJ
DQW1/sBaK5+C+0d5fRPEmJvguJMSE1HU22jv8VTBVFWYzBsJmS4F7Ze+cxn7cmnM
ekTn3/RG+h9lHfXj0Wq+fkFmvK9w/BjaYPW2xK2qVVbCKTIZuSuLtYoAAMsMaVMN
mawdvMzm9F3EOxhGFgYD9jnbMvCOavnVyVrvFCCny+23akq96rlThOKUev+ef1iY
BJ6HsYk8gOk+9bC2xfcSq9hFN5Uo0yp4qBdVKjkInPDFzic+rBlq3GesvawubF76
bgevgSkDKhvsS8vfBu/7+WiHYt+9VuJ5/b5SKObd+kxsgyeC4qg0LqhBtjgmLIgA
vrIqmOZ9bPAAI7Z5x0NgPiV9etl2DnEmrZQtYjOJJ5kaKRS86ZOyaer7/T3bfutz
FXfHAlhoMDAf2V5mzUCJ21pzB365cOF6kc2pym3LXTIzCipZWRfwom9RqeqvYo3Y
ZG+D4AvFcoZ0crwnR8iM/RrUuQdwyXi5PL9m7snmNvJwMyj8QazNrFR5wFtWq5Tg
xBsM6V5BDT3ElEckoDllSBo+09drzG9JfxNwysLta9hGPCbLRook9HsmJ9+lNe90
19dh3pdICCkvmVAUjFx7LD/RgSXS6RX7ldHOcblQj2NoA7/UlyrTij0fuUq6nEW2
Vv+vBOaJe/5vTVm/7wza8UHUxAJkDx5ZIO/Qc/zu9KGEKuhNOHzyysi6WxR93ibo
atNDvgperS8WZPEJwEqbNzauKwzU79o2tgN124Q+JK72FuWgPurnMqB3T+tkI1Kb
ZSxr8DSE8Ng7/CkjeHpD6KMm7B+pj3Qe4IDALsfNeZVsZTRkVqSacwcEcBs/beL8
ev8cncNOcJTVw9GyGYC5x2jxSJO5tlDpdyoSjpmA6cx6kI0qNLendpsdIdoj/swx
AZyBVxSOFd4DsmLnwEz7FIpAMKuUNTallNAcCC8g3LzYeBFV2nPOO6q7XYFBgfr5
JmL1RLj3lOsKSk4SkVFjQgDUdsMy9ncuobGmWuydf8lPRp+ahjRBWztiBS2GsSUn
756zXXjj7Q3uUjhP8UTWQlZbkcDDkvehUbk/yZt8ADpym2faGJkbCs8nUcOXz9s2
o7eHznrIjdKwBhSyKnfcMytyd0AiFWOjJhOI+NgPWln5DA5l3CTBsT6McUqqkHkS
l8PDiFrKiPtaUR8J36MpLmLSkXXL0VaHNVCAfeRJIw2mpwUfTfhHaHBBH/dOxgpi
CtgnxN1gwbI4e5w04ndJlqQHPSMnne1/lE6ClLwW+2FwPXnZ+A8quW+ffv0YHnWn
tcM13g9KDa8r5ObSkRECUolI3fTo7+rErC5686m2Gx8COxwDUKjLuICMWgybc0nz
ayj+bQa53N07Rc9T7Y3yi3315onpgHT18wYQnrcm+5YsQvij1ZFB7RmV02qlvX+I
3/tVXq1VVY3E1NO0a0AR0IgitxEhUsm018c/exjbKF2TyZWQif5+EkB6w8SIP66f
XMq8ZjC4OL1BfJK/QXLCCPQ6g0Amias91mWFOBlF6ONAsXJMlhRDKQY5Lasr5SE8
1E0PEU13qeLHqGbPZ+uRwrrmjEr2QHnrCUZXY+/05Obpx8iDhGlq5BFxkbx53xOq
Q0/DuaaLtHHefJ3Izr9JQrXsp1DfIWwXs5nG5WdZNUiUw0XVnlscPkXnxzHlq1BW
FUTQuN+ekePGBd4AqJnjsBJOIK5F9QXmg1uya0ufHGO66HC5drATi3GNzUuwvBQD
qWxjcJycJHo6d4eWq1vAsp3ynPfHhwRqkGHptXwcWgcvA+bJHvew6m+MkVhOgZF6
o92F3iOJ+cJhjtAWCKVzuset29N63m41y4xyR40MtENtqDYoEmnQu31mB7/8PzMt
YYt0tYLHIGVx5lNATRtc/WVVTHE44obLjL7fO8/M5Rquhrlk2T+x/OgLBlm8ncqv
3qetOYwz98ibqtLMp5r0Ga88mkYqu0c7tSUxF+o6O6vXl4QHqP0EC9ZgsnJFgQYT
i5CLpSsrSMvXpexbwFc82XaRSdOunLU+PRXacCdTwBha43KmfPMjUFojLzrP/3bg
LFQdwAjHgJP6SiVm2ryhYdezGrlW/5wEX5ev76W1HUhCejgDvsefeqy83Y7s0qkN
wtnzMZL7e79ffjTndTXS799ltcQZX3h+Q2+X+Vxo1N3q+Z7GhlEJmTXD/t3t50oZ
Mov2EtLRvhIbmk4YeNizkPImtMev3y0Ad3mP8slPfWxkCce/OV4+hnIXe+gCi6l7
/et14mxJczI2T39kNniaRWfsF+H7WleD0PBx10jKxjwvMFKoLEn03AMjFJd3nV8b
K12bQCQjMEyKLcCsk2feQb+y63N6QYxRJMjvufFdXcc0fG9Jly8aR5qI82gGgBbf
X7zoPWyyt+bPqSBYAZX1iYfz1E1uo+4Zbt/24H10mTHoGZs0CzBgKvmxfYqm4wvJ
svjJ8YrWcSxzV9RqL/3HRjOC+paL990UgJIQF5K2iMhbFJnEdg/VhWJ4UZNAydvh
J+lBS/fYd1RXh5DIA/peGhm/hSPAUgFBy+A+5wKg/kPGFtDqTWUTSBM2UsjRx4Wk
sE3nHQ1aLhSrCDDhRYHLU3MMgSJI7OhFH8UFDuoEw+tI8X+q0K3xAXfj2nl/FG20
mf83MOQyY/Pl9Zlv1Hm7MVJJS/aY58SY+snHRiWHJmtjKwG4KlrSnWtGg4zXq4da
CVC5lCd4mfzKJDWiOvAtvafbU4PfDyQLn4W8yWOm8hikd8FpVXSnorVxbPPiSsKT
jJePx8qU0i2WgWV/EGeJKVXSGAaspaeJrUOdnHvKlzDNgjz46xKhZbQUVw+hJ7jv
HizeufxBdSVdgBsljD2qqm/7xkpAwR8E89FXPJIWZ7tp0XyjprTYfCdpLThCU3gB
WfDsnqtrERVhGQlLyeWt3wvW1Sel/DI65ZgAJFu1p2LR5uIpUzN67sPjb396pXbe
tujAKtXqG3F5T1qXk2Lt8CEE0IaMVPguhez9HQQCdIq5gefWFHpm2QNBLgsGAqnG
wzNW4tfFCYgjEPUe9BFbK8qsL8UkZgrC8LXP7M/tayJcv+VQJVE1hwQ9ZkCrmHvP
Qgh+9/CWJdf0MTCCLl8uyT9ESoCUPm4IO/xZp6C4dtrEfIVCyvK3dwnWbud5V899
PDbPc2Jj3dWVrzS7eywiEzINDL8Uxb6UQ2WyhsETCu0NqJ77X5wKQtDmHvfUfkFd
tOnOcdSq6VLa/aYIzQAOv3Ae9nCdV6N62WyqGjXK7N3wz0pUptiSOFXVU9Y/oab+
oUYOk9pgg1aLzb5UnBqMOFSI2JyR0GxZE6rzkMQAm7Jw3eNh+nNJW8Hc9Rn7rtrk
Upg3bw76cdjhyCxXCdSu2i1UnPRarkS5w+kqC+Yk7iT7Ob4hqGkdiveqIcDa3mm/
ASndYboRMiq+aTz9Vbg4I7/++8J0kBzmAo/FymRsXim0muDZiBuqunVu6NwcaEcJ
X2xW1Dotay+6MFTGU5kAVYPxU50GDiTrzLOL+P674brPL6OvR9uKNYTYQp3LzkLI
ycMaybwGiaQC4t613hjJpy/aDaVtrV/mGQx1ZAa8OwS10wIeERKGQxXnTSCU5MwF
CET8I2633FOf2aK+q1TUTMR4eYLC63hUWHGnryn+9VcuQ+lti6EufxyLc0KAEqn7
qp/tq9j1TpGGDE5eCgXe+sYB1Fj4YEc84hiNpDzA0/1478h9J8aSmaRPYkcB0PCS
J+KXFGvsfiGgGx50cFoZ0QemACp5VGTk3o8GPbXP4Y8o9PrhXMA0i9WRsTZcnirA
dDMYlXsl4kq0I80OILhlehnyTzGGi+XqfiW+5qscBvHizCXbhQ/AUU7RXvPQ0Nf2
JYprQa++CvBoNfI80SFoqvWUbZTEp7CZ12zBbCiEkhK4OORlrU7MppyN1IWhy3MB
74o/jTdQiIA3ZIXnC5L/sMvCf5AcJL46OTbPkBYWHYbNJ2PDI6daxEGQPHXugSbW
tTlPD4AlNleW3kM8Fm9PiNY65Gi6bCFYZtoO5RoMqgrOQ0e+/DX0dPgcNgLIf5qq
+HzE5oDrKuOkVYg2C0zRVc+NzpV8t5B1oeJVS1ccLvhoG5J+mMzWTKHcD1LrUJ86
tZLvvSExv/NH91qhM5aXCwEOZVeTCu+rkCMYgXg61AE1ZqDXgieH4X+/vZDI12Gb
7CtddBpDv31ymXyFWlJ6dM+LQUeuc0gX2nZuSr3fnAkc3uZBjtcwTAlRxUdOABCg
eBpBUMKM29Hi96II3Rw+/ryjhol4gAilVQh/SqkzXRwcAbxUWzOn0iTuaEKkXa4f
FWRfw2HVCoRJSSzLnVm+0Kp2jNY8sJv3yAMaGQCNfKzZiqinfJjr/QWDw3Vh3w0y
/qjAS4/ZmLiK2Wro1QO4fLyW5DghKhs+0E7SOcRCNACrbOtmlZalnDQoDk5MAjx/
VXk0OshuI8jN0HeGEzmVRmCRgEGjs/v7WRumWekD62evs/sPCfH1QYjoYZjfnnZn
hCmYQzjf/Skl9lUWnaSGhOA+scqJ/pRcZYfUUOOGfQ4nztrklYADng5ZwBfGcj3I
vKYZmb52pRblOXz0jJhvJxxgqj81xUcKEA/r+q/wIUyEWWyik4masP9+9prDOUNE
j96nPn7NyQXDn/WFQdw3effFKq5Zh/iVH6Rk/Vnpxk+eBWlFTT0jwrkFJJYUgAjE
coYVEJ1w7NsK0dWqKyFtEjlvJ5rA8PK0LmfxagFFZFam9J0uH445Bhzi/sRp7S6U
Qf4za+UrLXXOZ7rbwokE1PyJSlMgZLVWGdjX4rN7pyppQPnvFrBuGQhFm6/7qGMQ
evO4AtrsLi5n2Em+A9lIWwh2naxJIkZep9GOxliD+iEgxe4U9EuOHqJK6+/TYA0u
2dhoWsNB9RsT9gDf3OY6BCzx1muFLuS18kziJ3Syh2c832ZN8hMwcNNQOgRO2vMV
vhvFGEpkj1NNlLTQC1wIGyYhUwl9rJ1uO15Yi2MKdmqtykAOXGPx1DKYm2dhGRBu
sqixswV6ftnkP8PNIVd5/pyEpBvDGzaeTcPaSfYGvejcaBd0NNz4jdGxmQ1uPZUD
86EjQEUI5pTwxKEzwtCEPEyx5AC5JFrheSrbXEeN5AxSXCcpCQgiiTklHJKv/Ox6
N5OfDJVlSuz4cez4FzJnBLx/LVTDMeCrnU79ejZNhaeLrhbHEJukTxZ+upEZrT59
D8Okm7RgFIkHFYriQJuIcbshLHI6wyxbYe09UVoEM7C9XpgGim7bDkP4rG3/Ro7f
plGYFOgVWrZ4ejbpQeS4EDiVQnJniU5/cMhAvyRNKO13XTZWLfWdnD5I/FNmbyHv
5d418k2l1JoviZ6PI657ozr2rbsoXjA4qLuI8ZJpS2FOyWKUZxIGcPeydZSQDXtA
Q1aULV5m3pwaxOp9yNI0nWi3p0JPSL6Vu3KmuFTeWDGA2RaH5rxAKWkp/Q7eo+ER
NEwH6og0TZ3G5JzjuCR7T5AdeJAc5GRSPYtSwjxUZB70AqUH88rZP7/gvJ+0CoBg
PY5bqi6HfzsVTI1+47xLnVjjYWhCqCCW6TpAgoWFmeU1J7BxXTp6zZAt+rn4E6MA
jhqSTs/zn8TG3dnbVKa7/+dyNRQnlF7DEuwxNV8BReqnKSsI1vT7auJihDDfJtdx
nJZmkXEjaKuWFrO9yFw8mVhkjQYZYsvrFhNggKJT0Qj3O9TWrDgEsidAGqUuxVcW
ClQgchGuykg762vAJNXKmnQF9/rg/4lCs1uAgUf2qTdiMKpRMxky3cFtxIl1QFWH
ELtdIYBk7j+H9ckV84x9/l8p6Q0FiboAf3Freq+rywZYaY7aToKoYZwKmgvrh9th
ZvA6KRG4EmedTjg03ki5MExLHvdRT5g7/5VY8pMKMeJGMhoMIHeAhsnDhwG/K8cY
FIOcOHFb3EkVoAa0HCMjBeanjGhVR3fV9Bnpg+1XhS5rDfvGy9wA65vlN11kKaPJ
u0FS+eAgEehcPJ4kxN4n6/bnXXZHv/9a1GX5DatPrqD8lXExUwc2qnCgIU26V/Y4
gqvyZfbc2/q6EhKdOq0j4Ulws851BrP8sfXdJfvsqsIcejU6vR0GNqB3ucSuUPs1
VmzSMdGQWCi95yxYfJlEhMEMcAO8UXzgrG033FPtJyRVKh6GUtDRmjwr4zUvxoGD
2A0aFFwGs4cZtNkAJ5FU5knB5kyS3WYio9O6MRz24fWY6O2V8n2RqGiJllyynO1j
u45hi4Oq8xYpnUyl3Nb5/EGDm9JnfVlvXfnT59ysEtus95e4Sa4jLJRWX0G35ZIr
W6ToEfGYxEByl5oXZahjNQyFGY8j3ZAPWYOHii1n6pOW2BeKc7Auwhoe2/4WPshS
Gkwrc/FuVYrrmY/6BfDHKH8JSdJyBvfy0c44luPMs7iaXP6XM85oEnBDB6WpD9kq
pCwNbvhc9WP17bK+lcXl5Cm4ncu+goHDGJYWrgjEfyc4kIHGNXM4XMCQBHcdtN1v
JBF/lvyD14EYfX/4du3jkRDJb4A8iwefMxxz1eEim80ebGzkXSXV1VesMSNenweO
2NlN/nbWI3so3QnTljx6GBfqdOevdLLeitWuBM9QqipNtpuAa4hUeWn1NdCuNJUI
/pnW6uAXFa/iycAJ9T72J783LprI+1fNEAK6Kx1Dzt5wvv6An80tMrs+G8iZXiXC
KOJpqxcZUaHlkn3EP9uxPwih7EN7oq0FwMgJkRbx8xSlfPd1zI5lBM0VQXH/fVNU
QMzJXjk37eBOx2dgxvV0LdYJV5njdPtnQpvdx/uXXGhOtCbi8++dbi5e1bHrMhm+
3VJOzQ7DYrafgfud1PjMwk5xblIIzjoTLjFNvCKcCfc=
`pragma protect end_protected
