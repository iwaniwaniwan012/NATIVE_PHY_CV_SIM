`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
t9DlFGyHneHX93ha2Z2Gd2kGji3Uu2eGuOG2t2MuZ5I10OokdxIRcmy5CbuDsIy5
LRQT73G+zPr1Nq9rmyETptjm1fGmgYBzm7K3Wkkxrl9OPBcL6TQF82QhX/BgjEoV
1kV8XAYJgWesIGTtFS9GQxFos3XF3aybec9lGRpD6zE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6944)
SQx147KK6YtT0nCq5SUn3V7XqCoEXgmuo4IAeayQ1JPnofyV8GR9bZVWm9HtNra6
NTuqUDwUjAjBLb1THT2tsVUgyZ2aZFFdByl1LGigvsoPuUY/ZzPdzB3LOWKAgK7e
UnQ2G2gAL5WxRXLxAAfipAsIo8xKZAIb8YtCD1TCI4OtLDxllHdrIE2ys/TuTHJ1
TKu5dpVovnAS0sePYj6SVuI74LX47xX1OtpPuU5VYt2oeDpesYpt66ySAvRxkBlE
E9Vn/NaUozuzT2JTJksF9ZhkxgWgDh995msJFB7GVufVGIYVGdeBchUF1J99nYkW
J3NxVVikfXkFWiSR2k7h9u9yi2e9WOh8EhqUeYyMZrmUqxqPjTZkEDrUtBY3KV5u
scaomKO7ojh/zs868vKHvXKfz8xAd6qTp+6PDKSkVgZX7CAoEQ9QCMmno2dIf7XH
Qp2NBF/Eu4HqypvIbrNgEaQecfODb1cqGzHpXVLE+m1Opsm6nC3UVk8b1VhnZCqB
SZ4JGjWSyxuxdSaUdbXKdbD63Tq8lEBZAZfxFWvn8hnuHgFTkEoqLAwNe9Jpaq0g
LyVxw7SZSvTv+k8iXp8ZPzHgPOnVgwIX7Hdy169kgdM50WJEvfMZQqJojPYsGmER
G+gBZxe+CFsAhxV0sR920jYFGOLQAp4AxumQn33E+PgNMzHo13VZgTZuzblxrv9Y
/iuP776PWHdMXY6V0mSSAYnew2eRq6AohKoHDC1NtE173IsucZeGrZBES3ih1GGX
WylqbPOQ9usaRRiEL+rZhqYZAqijaNqOa5twF7L+ETQ79lZYD9o2UUexr0owqlQU
ccFjx4nPxgg/xmNgcvsX4AgRE02twowBP7CvhLQCh5zpIb753NiAwVhUdDzNn1z5
RTPHMsvKytw3bdIDu/xut8PFNymRUa7eBcaU8WgXvfEeamZctWE/Xtdr01Z3HWFs
pHEJwqYWxieh/uWmyCCFbll1Te3TdZYkc9O78yAEDWjfl/4ztrjLeoHXjVxJcyJG
NmptIaSU5UI3qpSvzAE5WAAwzwqoY3A0DN456mVbMTVPi6mukZgkHVvQ3OkccDW+
OMVvpi904GD+d1CvXKeODMKBlNDofxyIk7V4wCmXcbO7FhQJmlQwhjgvzFo0Ml+O
aHoCo0e7Zh6vH5mc23WQJlGBo9dnEVHZnWBXNweW94usvIQY2T5zDJ41ZGZg5jEe
vmNMApAWP5IZZe0uHLzihPRskrVJaGUXxFyapeHAefkZNJBbJ00L3/CRhQnRRDPi
2yezuEbGJi12aEhHFm2MJEnhUjlE/wwrkT/NpWfiFoWp/o1qOsZDxX1q/k/WQCZX
HVJ6ZvZ6N2rf1l3ebsNOaJraBtmgxzU6s66XzTrHBj/Svqmel1oA8Hb9/Ud6PTQ9
6lYYgP5W57xBUAeYeI57YAMBI2D8YDt6QiliIUljZt2LewmjaTSmkqru8IcW2HaX
e2/V/ySXgh9fXwp1l9jnUk3tvZRm+GQJ6MEFGEmmvIDg+3arHda1B1awoNW1IX77
Lff2NIEvcmSjepT+2S/GvUI4zyMpmVv/tSkgbr5h2qbAECKpYWh9COo1tjDx/hp8
dGWqFgY/dy+rQwmK8kyFTE15Rux2YqEGREMSd+M+8fFeZLFXF8ED8RujPbL0Ixq/
D52TR4WwffeapPgluZe4aouJUSFdx3MS3S58pCLcolIBBKaQ8xYRGjeYVErO3S7o
9vxLpic3GW/fo2xVhD360/n2AKekp0PDNl7NVpsSPP6M0rk8bKTDNIuPZvo7aAMZ
TSHvxBW9QOm7Avap0CoJk4vUORWhiobIUqNTrtVA5o5vdkITY7P2ZrqP9kjnci2K
8CEMEiU0ZfTSxA0Ev2MekrX8GYdgQjnLSZI+J+6nhuFlWWyO4eVA3ZOpvnC7rgxr
0BnuazWqjqF+deU/SOYg/HesA2K0ET9YwVXUtIk1qKRoZsS7Pm4FX1i4tW0Ew2FD
ZGx0/iFzNq8COiXWKbm193kgBznfVs2DnBD7ean7A5FDPceqUK7oZ04GboxIJzVc
99ekKuDOHB2qzJfr94FOxvTkJdm6nc0LhMz4C55BtmAXLfULUC98TGkATTxjbV33
WYeCOKC+haZ5+ohYDM8JAIbnxYe44t48knuVc+TubdW38FWXjStb6sjgCCDdTaEg
GPPrv2l70EkcL5oo6rQFBvtH9hA+D8Mj6ty8kc/OfnLMHHi82AeuuuHcBpKEpEWk
esTDc04oUIOUE3DKuGS6toVUnp6iaEQrCS7VApjYWC5jD4TOJPwVLRWn+55Uz8/t
Dm/9nzGoV6kRo6pKa/9jaYyG8IwqAMrRbgkff0oIXTwhreWEHi1oBJDL7iNaKjq7
c/LpayPHL3dB6UV3fI3sEfJALeGGRR0FlunSONgto+SfggHDmJfHFD0bEAOYhXqy
dv2nUvTAFAFE39gzfl1ixyP+1U3c1PzKfFPwttS4aHQfE6M5aTmvL8WnJVcmMaF2
FZ7p3DiVUQbmM5V5cHZUItqrdgnz3ChQE/HPn7cz/iMo0TK6OVRVHZ8Iy23uCeNB
Ju+SHw3Lf+QLsEAO3xjo4cyEWXaWcTzn+XoB2xGEgErjmNSqzCxhyJzqsBM2KnGi
uMs2exUaTvu9DbEi771UAwn/uJQDatDt5x7l7mqJgPFUBpjyq90VgVURGdxm+sK6
AjTQuzROATonyWrceFfzCLgnX7ZxUyAibu6no7M0dXAYOYvf02Wba/FWrIdir71i
Ie+Tw53hf2BSq5Rb0I6cA5NApVVDS3q9wpdBNWuuQeny6Trdrlfxx9m96/s+KfNa
PSzgmarOwHnLAsC437WYAC8YL2CJAMLE5KcgEVkEGMFI7MHEUTjSuXfCpGhmllnk
aBfBSJv93Fxbqpfkrv1JC81CWf316vJHqRj4Tr2Q0jw+OdZcIWeG/tQNkfHTOASr
Gp9eth6rS+PkiFqIPsbjlVE0i77MHIpq45iOGs3DKTu9FqRcVoiZcOI88Z5Qybpu
wkU7WsNnuTfbTWDh+g01sxwSip1O39R40w1oQx3KICsma1VhSPsRFlLd32DEKdkT
C0sf3C+nmD9NHEKHX+qJEsJDsloy+IpZXflLNSu3ixT13eeoXqZh6WBqE8EuM0W8
+1dc/bcf6kmvj/dyIjehOGq8U8e2vdojt5fMvCQaXPu7lzXFBZ65escm9I1jOEDT
JcCX/8xhHJ1H8iS3ynybqZObDwjm7qs21IZHx5xgU8J7hfk9oXRzvYPLTQu9HGeI
JsIA5+HhFbveTbuMxPFV+BP7oZ1rsAOgHWIu25c/pHUG7JM9zq4TpCT0Ew+Uu/OL
AGzG7PRibNzfWSqN1ONnevRyWHGtJB5RAUgZ7AIpyiK6zRQQqoqe7pWecQjqP7rg
h36/p5hZx2gjFhqKIOE5EqruuhTm28mKDAfS1txb3ViZ40FJOC5bTBXnG04Nltfb
aqZLdMdzraTz087d7gQia2CJLQAs3AWyF8KOOU6TvsnGxKHOGRMIw0N4efqz5ACO
z/xEGOL4HAQlWrKcc2XFuXFidJ1PzmycVXtC1oxMuncJlzLiJnfRX2E3xDDriie1
TWyqvUboLr8O2h0aTM551ussQH7ztnnNNDioosURJtregKIXyqZUTGiWng8BoNaP
Q5/D0eyJitesnpRXemo956XLdlWZfNO61sA/u8C+xGqTKvDglT7Eeue94toW0ayk
xAQ0lOXcBCWMCtbSg3vHFl/S1s6v3UF+dEWHAB5VsJZN5xdpoB/tdLIyvAKw8OJ8
UsOx5xvZ6IeNDC2ep4ysF75sjKmcoOoHSFsVk6Kj+7R3FD9hAQf7B8zmrRfr6qfG
9+49NK5RDUNlP67pOhm/HT6vf1WPugkBhtaSYWBiPRCxkDjnt7Yjb9LyuYIdZuJY
7xE7omnp9XIhK3Qs+Ghx97Y6Id1yeJejrsO0qFMNRKRymC0eLRr3pIQfxz1RBDAC
IAdtKobATsC2yf6NFgKi8jD1an6Sw8+rf1SsNP+kI3ig9NQxxNgkAoZqECITxjGU
Ej8jNXwoXwcEvySqaPFhwTJNsz8K2wQ/qIk2OzD+464rBcRgb8mUr74aSkjcURp1
NEaK0xIQWL9j7Ijzq2cujtHcQSMDCg5L1/wGf1TBpLNjLEje/sNFDYkIfxuxg6z2
+vztXnCBgeusk2gA6OPmzQsd/ikjODUvvJIPk6sYKBG250cxtuUrTdb1l5lZVJc9
16IwSGfg28vLGn0Wma+j98aZuxM24UvNzOxz56k43a/pjfRvKvoXJKxZa3os1oVS
pW7sGGYYFJtacAnt3CHqshcbIMf/1T7XWBijofybQmcsFiNHlY3V9oQQn+XtlhTe
JSQ9bokD3zvTRF3z9xkB42m9s7HmU0PqMqtwcGTxkvBsw78L6aqA09f0y3nCpaGY
GyT8kYzi6bbHOJ/XzeEB11kvjZ8L4Bq8ekZtF1el18BIWnfCTjLOVpX/+LtckD8m
vGv8Lh6Kv57DrWLEUBCUMwk4tsx1OiuhV1GTcct9Z8Z1Wjlem3Mo7T8aIhKam5OJ
n1/wZ1MqN0/FhVwQsB+u6eDGH77WeQvda4mv4dfugvWeE1SboMABIAn2umrNyzGX
nyIni+jcFLvoukCCj3sK9wr/oYcOe9AFo62aBSSWDn5c46s7Gjdt8j6MiFwbp/Wk
dej8AThSo7wrL1VYv+Q8Cu7majHMm9B050SbMHME0iCRYY2w/NpVFyq0NP2z3xAn
GbZUE1DdutuYbmPhpr3BwvijNXydfwdQaKi2ZWVuL6ApYT8jBHVwvkcg7tOWxz5K
tcArW/LDtZpHpvVS36cn3+EAd/7qJlXWRsxH74glm/HrFp9ILN4hlAPNI1dErfv/
V2h6k0AdCvnH2bwLhwas5M4BSMofzV6e5NTNYJ2MDjKkyAzwD2/TmyHOSthFC52K
XMjqflXaaT72cx7FV32G+OSdsxuq2gikY5pu0AFTamOjfNAuopWOmXY9u87dhRw3
2TCMYgaGvBL0cB608zLAn+Ys/ooXKDDyRiwgKoAkWiQYz9laPevI1Fc3TjFS+hn1
to2adKoDl83tNo6NrqATOh3Mt55zjMBwv+mAXAw6y9hrXTSKakky5uADjlZv/UH5
dNM1qsj55hmPe2+rPVkVUGJa1Jb/2sEipfOOPAYas+cO/0RIlvJ+U4In0cUXs5cm
G8+x+BogTqkbbWFxIMMJKEc7ywaBvvwqvj2L6rwTEP+MCAk1btjaGyv7Amn1NGdS
n5qq5NYp+GU1R3PQX49Scmh2ExV15+GbdLBS30K3a354TMZQmiq7K2FPKiFt9C+B
Ws/Sb6DOXoeGvrXNMPqDX+b1oV5nfA2BEfFx/ihCOZgQVYLrG7JzAuh1/FBozfe7
Q57WxER6vOdaM5cQfv07mKHCm0O+pdWetwIRgCgK5s1pBK+sVpRfqTwvt77xRsJK
BNLNAbLO+e+2WHINHbAPVp56PVnOAIHdPtvcqJyWYCIwubIJvxYHhX39QQi+31pQ
Nd6qwzyp7s8YPCp61rrvsv66X81FcPOwnwKdnjIlVxm+hAb7Z4FCCxTzkDSdrwOU
12iAnbC2W4Zo2aupi4RZBYdTu4wGag8kWCC/fjZEeNyJwAeVbsu1pDPXIL2OEAEj
rkITpZ5KMKV0iTkS3PUhnZJa0pgVTxrArWrXna7XpcFSmQaGNhJM2SRytCKU0fl2
LyxOHgYaSmLyfJ9Tds6BRruHdsE1dNcVDGDQ3mbpCau2yv6+W9RCK0Ui7v4iLRi7
aDhucPH7ljv75WF8IwkyQ9bIKDPxGle4MPakBxxWpgAODbo2n/vBYEEU4KPrdKx4
hUz4h07eWnNhbrbhgeGV5IE5F8EM3Kw0QHwoatRF941Y1ydyi89fJqZs3LdsAMVe
NL+p/iWvfLJQdYCYZtqjh76Lgv9Ks49B7+0tRup+cgmAgfcdS86uk+p+GTOgrTCc
bYVAksXu7L7msAnkrKp9qpg0NQnush4OZBobC2A0TfdWkuley7I76uRJkwYa3omX
U5BW5chSnAIUKj4skTGLZDrVrbGNvFQCFTITLCMhzWvngqSkcq2wZ8zmT0AUlBJM
Uxi/g1UhNn+SAVXZVTrWHhSX+upRRscnHGHCWIqfxKMNPW5sIn/uf3zu/hvXR1ww
MRXeB2sUnl1/URO4vimOnbE7IYzsMvO1xDyf3hL1uqfHKXsfRb5NUJcdLf9+uLtg
IMCAMfSxDG1aJa7OG6OTCNVgzPXmIAtFtxNJS0EhHtI2U6cXU8Zag0W2wXTi7L0i
AfRJClxY7zYDZMv1lkZy/gE4IBovbooXhw2NxzsjOHyMFFPZOiPCLOiBAayYTERM
drJSGQuneJSrddyTXg0EAj4t3mi8UW2dhZm6daCweqGTONcSH/BK5WSgG1uScdqP
kxFKCfNHiveaggQ61D7d0QqNdt293Y5TbK8kVohGi0MpC6m6H2OcIpxH8IC1rgt/
/n3bxa6Cdht/fPHbxbGfBufz2rfGrLr7uewLxRl5RZttB8J42uVYh4Yj0kl1vaOj
NnQeNx5fJtap4PjiwDFp19zAymIrP0uNxNM0KG52n1GLqJeI7POx8ucXSPN7LQn3
Y1omuy9YE4td6Gi0wRGP3SJsfW4oChT51mvB3RkIpV+LEY6R4xMnxjGHQ8+RHMAr
aB9EuuoJATFCtdBmAuFZTUN2FtnTOKaDyBO5vVPwPlkvr1dUBVUIUlXMZ+j97+cV
lqFA21mpbo9V2E0xs9zgY+YmPxcR6b/gBQYxzTueBlVLcjBl1e8rwQuzK0/xyLzw
bYT/Qu6fmPRsOHUnTU2mB0TQ02TF2BuTXMRqAPsyWs0f+tzO2c4HPLj1eRhwcVxs
oDa2YYp+9G55doH55/TEhBLTiYhTYry5frRaakUHzqIhCDXPVh2NbxGjgkG2OXqG
C6ZCj7fxridgr36IIMFEGghOBX9+FLZegzrX/LfjXVEKemOB/xRLQhmea7aCTw6k
VNOMoLu35RrtdCE80zplsdVa89tJQy3ZVvwypd46bFwmuvnSonvZDMDdmQYUxpXQ
Qus1ZJCCY2B9j5zo6TDCmaf+QVppHkmpfis3ZzYZ1fbCehYYj0YLjLjtM44JnCna
YXWaRlRxXpIfwTlLKWeHO4KpJMGjuuEuRuBhferSC7ZDKsMsS36G8gcPBuSxgE2F
RjsJoMB/D6xOSlaDsE8OXDgVI9y5pt0Na9D0neyzjYS9PTzsfL/MNdIXy1/LP6jh
15EGm5a4nYm30dGicC+yKmpg/2ihBi5f+gY5+s28Lwau+l3yD27s/BseiKSYlEsj
F5MXD1Jtadf5GlSE8Aq6j3tELCKR9X0ZU80N7KN8BR/nrDVKOzOK4abtQvUWvuiK
NfZ8Frkwni5glm6YO/uxT6h7RXXi01Qp7bhE5FFX5aX8SFK7iTsV8asS6Z1vPPfK
wti+f/qavA0MDl00bBjPOGgpztnagsBuIpHTNUHc5eIEB99zRl8VpVucHHzKB0an
v760AC9eZzkuCnQZ+dqOnIwW0tGY1vgz257z+QanQrqjBQFxrXT6J5PrG92MZdG9
9cdIADjngTUoeJzpaFZ+iG4fEMucTiJf5lyMKwHDFk4sbfc3LXCh5bybJ7NVbgqs
e6R5Kuwmk3RFMnTbal+DHm5EBgC+OjaH1kaHKBZ0WRWrqU8JCfub/CZm8EEgBmri
EloWljRVnPqNOVCai+lTr+NTCVVyCBxMGuW1vh4Eyo2h17rCvMJqwahbu12phYs+
5zAqjQPeQiZ39YC4SN88IMAZ0g7yTiruOiDjFYmKD+3oKo0UF+HV/Vq1lgC4HsY3
s7F7MCc3sVJ1nMjN328HwTYxBA8WHV2VpJKHCTBW99IbzyGsDvH2bcsnIE01JJlr
H7zBDw3NKf+MobCipK1tNBXq6aQUbnZ9ZA2N+0nSa17L9Gi6tapBWKgoO1khASk0
Nwapgabx/OF4x4T7haHt0ol+ocbO/DweGJjsIKYZSxGYWfRxcIOI41Wy4tqq+wnf
f7K/CUhrgJVjf6NQADl9yyjv/umEl2mEX3WaS5iTXTM8nHhuAeeaO/Xadn9+R1Wd
mGYLmZNF3SK4p+QF1mNT8spTf8wX0LrCAC112R2A5jJofKPa6nA1EOqkBqF4El+E
NFze8gnZ7fyd+PvfBigWWu73kj4gegC7jQ+JJycjejy43AruxW/iKDrhmJBmy+Gb
TXInVgUwz80plwSkHdbKeoO8ypmyOnHxQ/mjg09NCT8zMu2kERh14lSZHv8WM333
o5nDZ/kYbzLvUMWcjj111fOfUfjRSyNKyGhpZAkG859xSLvxGshbPY5Itug88VNh
YtruzP0iuRqk/gcnr66/Ll5rJrPl691ZJjufiQa9NB8uPL1EXz9w7D+aOZ1UA16s
6+JjqJPo93fPCdPIrF6QAgkG8aI1hwQC7IQ9FvJAO2gmve8qXfEElbB7EH2YaSRg
EDRpO3v9I58Ixs1mRRB/ucegKoHYlBk1DolMZh+VBsOUBvVTZI8W4rAXWjhW2kM1
xyDQmOTtjRvuPFVwvB4uIo2199mm3sVAmuYu/WcxZkIOEcWKMzZk0Ptx8Egcg92S
Z9lqTJkqvF3xOBN+ibYkftLLstaGS+cImWi8OTiU2JxjPGfLeVRTppsDPhW26FrO
Z/YnycH0q8DIFPYG0eNjPD6vd0zdhbhYqEKBMxB0To/xwH1cqtFpHpH7F5Xh5Xyq
d7RVl8ZUt6eNMqrLTwHNUJUWfWQdkK03KFqAdM3XnylPNtEgKfwYt0rlR6sZavMj
h7sQdihSK0lAeSffCsBWf1Y6FF9/DLHZ5oUgETDu+3PKgZgi9vfsAY2UUG6obn66
7+3D1y2K6ZcQzIHR2foN+KCRY9CzSJRXXbiskzqqXQ0hIzotDt0wdNOO5ByHmC6B
wWDF33a9Kc2M/H0U/AJouBz7LuBG16entA4nC+Av5tAgUV5BlH1XwPo+VbaIdmM2
JCnfHYIqjudzwngObT5PNT6+wf7dk59PTmJbrxv4uA78NHTdherPDNovDUTLDSqK
O0ZFlyq+eou0SK1Ad7j+K8AHDioSE+tY0Lfzxbr+6BU4xZu65y985aEMTXpNNaK4
h5PHsgYnNtHuzw8yi3oLxpfXqAtlaWl8fFHYoynqSROK1FkOB+jfl2iCKjdPuJ22
AkjtKdjMzQnYgDF5+/hOCludXq4xLkfgCXZChXDGsw3PK8spqMBrkCAQu9fHqiIj
eRW5qvG8hkIpZbGPSFhc0K1TkFPbgjFm9KdhCnPjwH8=
`pragma protect end_protected
