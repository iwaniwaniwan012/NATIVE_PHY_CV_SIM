`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
B4Rmh0XUXseqCdSCRGG7lWJMBzP9u4awowNpTqZDpE9KjnqnfSbCmPqjOxqKqspi
MfGwTIaWXdD5YfQLD0DfpypR8cGHHsV/1GIajE8aGUiPtuTVfKORlc62nW0O3vEx
pe9HyC6E3GQnHMEX2FJbfdRVWdW0hu6gGU1GkPBylNU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5488)
2mKCk8Iyc0XOpBN6aRzmv18fwmxjkGkRePz09qrCfay60pfFun1Y5jDZtiDF8bcb
L0AOMkAlhl2zXevp0MtNStd5YhHfFSdddMzwTAPXrZNsRxF2fbAU2UUqmxA5MNKl
foVdTvDVw7gYcfzIAbjhe9qHU30JX1McLHTd/PLq0kMPFaxNZdvzWlzRvi1HIA4M
722yLpzJxa0h7rjXqcoqc9nR9/tHsoH6NISQwsNhULvFYBbDnppmC9Ghdjl/2qvK
tGMbu7jHt3TpHFIZeqtQfOETBC1omRor6IEePI4R6RC5nCwUIcAhaKNfDjjcXdJu
cO2HZA1LG+QMjOICIxz1PD4jgefMyCHzRJPxV0eyWscRTz/kvHhfsyGUUv5mE7Io
WKGa4WI6/h6o1gfc7UfP/DZsKhzvY/byLbrXRJepAHq1hJIOFZomEX1pLL5reF+6
qpLbA5jDVqgN7wXCdXDmrq75HFWJ0I8IB5P/YpbL+Gu1DzQQIaX8mq/eezMdubdu
SUyn0n6oLVKHPEFDoC0o7LSZSFlmcpsHx2ef43M0m9HIFV5B2ljLPOYd81oFTB6o
hORh6IU/Udcr70OAZ8SxUEj09XXp+0/19iJf7AWAUFYNFKKt7nF4275uHB6/pJ12
24TM4cLyhLldHD2DM2c1OW99z0rzVpBB9Qmdf0XQpR21uHyIW3/n+r9m6Jafhe0M
z2MiQRb1Y+br0zX2+v9q8nTOQIdH1RSPFkIyzlu36t2soXkd13UIBy2mbAyVOUbb
oo1YSBCCA2hhy/AtPRjBRhV6dIeAZTtRy395q8Ho+1SVp0hqcUMsHKiPFfvVlJus
DVEl9EHPLg0vbeiZL+N/0jSnzC99tDPWSZCmbFMCfDzZZcMvD2aN6qwYVqbVjwF2
BBJw15Lt/5ftDGSHheTy8MomoadkGFmfIqlJJzUyswyqtKSlB9Hl8WjRm5Jr3n6M
h10wduooemRlTA7k1CgqBhALHR8RxEJSj4VTBm5suc7w+VJzrdnoSnMFPMQB8ExF
QY7UnqYrHGJJI+WnvyqziJ8mDDEcFnliSvNydrCknaSfm3aNGHmkmce27K2dNue+
7hE5UQc7rdeefarFdPi6yC40wWUhWkmph8LiDjwzbfrGHqvSX4YEiKgsgIzFaA9J
AatCIqWpBzcNE+qLO2amAhBe+wK6jkZwpKhQzXzQRPTSYHQUmALRyRBz1lmuMve9
fVS2UbZh/Yxr9xh6uXCeWsqu3NfZkZV7lWHRVDFJwI5yK8WxrrYB/vzULgvNRYbb
OOoQ8cVMsDF/PzvA3/WeHOzWrjEQG4z9V9OVceaItsXtRbpR01sgnmqh6oMJSqhm
iTXhnzc8ESRsVm/Qb3hKLlqc6NitYcEVg1y5dj2EvW9BCtsZcwK7vJEMZCouOmRv
1wLbp213bJVPJaBNCX49u8Kn5uYrQPxgx+owPRbGL8ROJ9MDjJBfxllAXSxYN7BH
mjZC9UHo+r+tf8/6hpVPhGH7bOIxZ+U4Ie+xRwjmuTjrU1Z1l94UBjkLUIYviwaz
S+OcI2uUA4+XC6NG62rmIik4YYkfPmJY8GrwvRKzrR9fROGWAy3/ps6fRvmEFxMn
UGh2AXEK/B6K4YlwitlzCRnq2WkhULr1Z6kVSeJuaCDHuEKtaYIKDSAm6IXvSG5P
Xvqh2bUGHXCxBKSxJygdw1X+M6BHMg6hD/aEFJevcQ85PLJhY14X5pdbB33sfh/P
LBgv//fS52H8G0qjAkohF6NCOIhRO0FbaMc3H5CNZtFJarS6IvPPLCorw4d8Dqyj
N60GY11MuDO6f4jP6d5Pm7LLlf1aSoXQh5cYJOrH4t6Yk0DFOdtmpo8Obw4LcBEx
8SXyX6VY9OBVLQGCOs9TGsjU5BHiugYx/jS0fgJ3Ht+H7NmT7z8Hp33jqvfIWJof
ladD1HRLN0sdwyWnGNWi9qQzTwDTXSjbo59qu2OJPNoFz2S91QnMPZc3d4rRMZ31
VcFqVJz21jBWAWBaWvuSkXPxn1KNkSaiga4Ljxu9npY8yzf/dSwAa4D81IIAu3F5
fXXpDVLi8uZwSIhpYi5nzztWPzXjW0+2TiKIW/1GemEwv2T5jYJrvSU0rfaUeO03
b5Fz90RL8PdxMeZ1f/a64rdGsd7uabYmmJ8HX3FDmUWGGguro0uPpK33rk1af7EK
5hf2i8EIGsze1MNcoSakyrdaESjWzC8DXsm235qLrJsYZV8hAPcBpSo5kNTRohM/
tquo6AkuhIlFViteJxq4I/tgYqXtT14wjXFlUb7lunmoms5wUEo/5k+dYU8Alt6P
0TblnLveh0HsN4qjA3MomHesbF2uXAhsiHjw9hmvrO8F/2z3L2nUipr4tiLkWqnO
4BZesxreMv3JwWx0jK6ea+nSO7VbQmvP/Ab5KPqxzl7B80cLW8UVfQFitSsnvJ2T
IbTMWKXN17a+Vbc+eJuKfBOr75PJHSvxopFrn6yuH3WfYUAmXvVIXVX7Ue2dKGE1
ny705yUgDq6Ta2aAJt0UQ0sDTzvWXjj9VahlDExVX8C8NYqW3s0UDr+h20gHgItg
bne13bf9QqfjRSiKsm5GW7gJAy4drilxUVwJYZw8Gv83P7xC8lbm3PP0w2NL/KaZ
pknlpwp5qJsiRCEVLx5q11Gp6CKNdOaUL9JydOdjZ70aDua2rwTD6RGESnUBrDYs
1liQWWqVj3JG5f2ktJ9zZW9fvb/M5E1ZKNmQ+0h4Hbl3UB9KUQANW0IjnOCKpw+t
A0Kk6iv/95YexrvEtD2tyTEHT6dP5Sa2tLFucxykDoj8HASCtF5A7ErBxrZeGapT
XHFoDW/5cv50PoJLvLBTB2odKEewN/uLlz+73DoBS26Agf8C+dqLA3xTOomQ4b3D
+BR6MoEesZjI4enBZGgqE0e2ajonduzfwFRSvqwwV5f50dkj7lQnTY9EcR0oN7xw
CkCNyq4eQ4aR9u7W5B3AMka8JGBQkpW1U8mgHJHZkvmCR8p0DLrGeO1/ThviY+cG
UTe7a6nZXT/Eb5oir1ia+MILnKuDp/cp9Fu3NJpKSjSPz/B/Ga17pYNWtvhxGWnY
7+MnBOyqBwY39R/kOcFIYdLPlLy7YYlzwNdicF2b2oeL0Z4JQzbq4UE3XoA3mLSq
z9/KC+/HintaXuPZ7HNnjPo2yiXdmYagQ/QsD21kgMg19YyW7txNYMNxalfPNqax
65Hy2BdqVSJ+j6KZOJajbSoksXIuHzQp+QRyVedD+X5B1ErnLEbXfXYOQCl/XhcY
FICwryF/Qs4sLo1aFAaIyMK3T1wwkgEvMKO4UeylgtK28hyGxo6nAORvKKFpo7jy
plvACWteD5+hFtuN2G2jBN6JU6W+pqYYrpKwf4kUbXqWbH86oFLI8sLeDwQrhNCm
z1Dq/mk1Dkg1Jx1aD91bHtLjBnn8cPsx2O8o6z80eKjqJiowt8vrfO8Zp+LLfcMd
vI1R/F/UUetwU8PIXj9f+rE7HA77zMydUz7GAko8SbfiQ3KRbMpDZAZ2jgr7VetN
gBXa9ByNDoCtYpDJtGaTJCj625kz7cMqFS5QNY05mtWapxGvIgdIFv3NIjQUqiXJ
mjOPko/d/JBNNTIvtGDvy6hMJJFkLSehuM1BsmqwdDf4pi9EbSH3MI2cKjisXpTn
/CG+wuxRRWOm4b2uO/pF8FXAZfGBIAUw9EJalerDVlVo7xbJBJU0vW0GtGQojzkd
/VreIzfiD3vn1H/XYmRXiYSjnq0OL6r3rvUoYBMoDU90mq0KxYACm9/3cEdX1WkE
LNEkBuAjJ/e8mhk5BNwXJSk/bUiW8ra1uMy/9kXj4iF+WpDr1aWuNJGeW+9n2AVy
6K95zjp5a2cnb2ue7ve+2vrHKT0AThorsytq0IKXJ4D4YC9K7LaREExv+/o9mHgG
ylSLelqWBpcxYchBAHnsNGJAXlohhpFXLvk0TfaCkdx9WSqWPY8zqLrt5xvefnF/
2YVAyNv9VOl9eI230T6A6aFto3DmnrBDA2AUii5k0qrVQZz1lSAFjzNlG/rKvmUT
qiCAArINOM5m69yK5wefRZGzN0MWmgvBxi6Vh6JfJK8asKUbUmhCj+99y2vShgCa
CU5x6ZJzTtmhNxKl6v848n8ntrHF7hIVXQH58z0Qx8ti/WPYnv25oFSaHSQfOOH9
IzkhA2mUnLXN9sKAOMQAddA4VQH0w1MG/60HstFac0A41jovKF3Yn70BCUufYwfX
qFDq1VbsxbnsqybP5PYnarFEgn44T69vDhRoHuUTOHKMJl0E8wILfrgTNDAkILMJ
7qWMKDXErgkp0sruQDGxwNztIwcvW5Y1At6H7IQPYq6xn1NT4P5jnIvopgq58ePm
HEKEn637cbNQhaJaYa6Nw5wrhO4D2fOhFAAqKcx9aD++EBMAAx4Vg5Sy4IadWFua
y4LiBVt2lTX9qsI6EAdgnNWTFyVdogJDfy+ch/eTdYKJ82mQKODu71DsCL4oUIIM
aXuoKJDaEhs4HKzeOaOZI+Ih0UgzlXiqwg3ksy+hqxIuT/hHa78pMKDMEUY6Zm+Z
c9Gs8tiD8E07tZ8/Gb7uTWqDWVQWpRXKxkivU1tqnu9JrSc+IXaYT4wzg4ZWd/gn
66dKC7uiTJZIF0wbx7IzTv2WHmc59WP6kG0HXuBRSsr++2LykXoE//TAtZO8s+xb
ZinPD7ZhieCxlYwW8TsS9MUwBDWgp9nc1l/79MrJD/Qg8PDsjWWQiwJckc7au7Z0
g4pruEcBQPMbw5M5zb+n86T2En8DMjWkhJRSs1Mp0ppU2sIfe3YpkiQw33dOFJdD
AQI9wHVef8ekxpmRGOdKChexR8JHx1/Rl6Gt7lSKg4TYQDCcmj+ORehGJkNhgf1C
vj3ba16eD6wVoxwNj27Qe0flxjXH9AF7Tt8ZDb83plIwN8jm3/I5QZ+rvCcARa17
UJ03fKrnv+W6vTIGV63v3LWzr7L8ueSFNnKokiM4SjWf6pvXfWVQoSw2iNJUOiyM
j3oeL1kPMzY8rKc0cwZrQ24034AKIgkPsDT+f9b5fllHw9HsT6JEeqcCDZ7HQaiB
bWIkkh7OoTzJ6RUUYuavSs4DVKPXpAUHCZ4UYWXz5J/NBs7sl8c/XGAz44CP854M
3RnspMoOgyvOH/aWP3zwKt3MXLQozbPzYAo0qFiQvihcO+Y/QNcmswNRM8UNLJBQ
huwL5Jmfm90HcxTjtGAdvfbQ/In9mbCLGtE/+YExnQb0OeAU5O0/Rx9b6mmbsNMA
tbj+KdlpjhK0KS9nNmD9plXlVLaAcWzIeJOjue+d4X9Qo305QdwT+Shx4ZhhAFtq
Lb+TYZURmxF0L8BaBEgLFBNb/zzgZ4DTQM8osZw4VVovFB3lVEVRyevjEfphj19s
r2s81BbrFA11WIjcNr5aq5Mv+E1ZFBmC5jqecWPSwsBYmCsif1E4ZNdVZZg3Ar9h
/NVr0V76kEUHOVXN0L9lgDw1gagD0sXo/i73DIlsmD3GuD8ERYx9qZyJvsIs1Sup
Sub77Boad8UQb3BhcGGFzLI+VYCnjG1d3Hne3TJQpOs1CANTZJkpFa7tW4ofc90Y
M9+0s2ucQ1xiv9n02QmPi0Pnqrysbxskf18LhzGVtNGCSC7+PkBf5oD/fJwgmEB7
aYvuBfwPXL3ibMFPhv+2buRi3QQHCdj2l6Ref9NHskZjt6+s5atFRjIdKc1qJ6Hs
7sqhJHC7WRYYI8HTwPjtyPYjnX0xNC7578klJLe2yjaiMU0ZXK3UcK03yCdAhgLe
kscV0OV9+efL4Xidv6dHZJZZrplgSudeeSX2mWgezvqe/flgOniBMZ09TZvqa4g7
IIOQGh68JUyV2JKeVgMYL+kZBYgbwWqrzOteDTGzb/D3UClNV5ZkcdvCZ7bI+gc4
ac209IFp5MAepqMwjNCgKptr/KI72FIv5O0HrcGZJQYh7CvvuYvSRKVj1cJ4grvB
YOzfWudj8E3mxqdQGNF4kIwOFmYbFKwKfm5JCsJ2MJWdGU5eUzWi4s6Y7wWVmM9z
zrN6q8wlA4tWGN6+5pCLmPuf5JlTJ2Ja4awAX+XR4jCJAtNE9OrZyapVE6KLp/Rk
wk6iFePq9QYXryiYsYelJJ9wOu4K2QQqZrVjEYeVddNWfSf7htSIxapEj2Tw0Tzz
lYnbEKFtJ4OoIDr+UnCMT+1qCufOiP52xuVbsvcvTDORgKuOdIohpYowaYd9Quh3
u0ZkrJLkNHtXWFmYsCSMZiAiReEN69iJre4aeTFZqd1I+HLXuvTRByOEzAQw1q/4
VN3LTVp3+5JusGFotNWwmowvDjEB8Ceor6EbpdCzrX2Q+ukWzIeJ6V7JRTAyiOzP
AOQAaLcalMwDJ9aFQuogHNWD/GeHjaoo7BdZCOgovbsEEh2jmJIfac5WR2R8rb2/
PBRhPGYeCZq0cinqz3dO2Xxdx0EWNRrAdwuhUOMGTfjXF3SxWP49VTGihqn2wF4f
nYHr9VLx60vf5Lc0nobZeqLl4+82OI/EbCrl8X/SxAcIilCjBkntyBeFE48n6VXY
JR4wIchu0ttho+Z+PC32j0ddRKbDAXH6ZmO4ApSLQD1ixHiWK4NuLrFibARzNqG+
geyLnR/NySbc+CUXO1BgEvpFTGypt0rFptrxMAHiyoSupHghMSl7/VZscGXNZ/1t
3qOznkQN2BNisWH2DFiuFMqxx3lPLqeJLKPt0QyPC8asIm71UYFrTOzadT+oFtpg
cdcgtUrwIBGlhg+StL6hqeFAA42kTGfwcYAt28lxUaS8KmOO6dXVclIvnsAGwp3R
mjphsUSdUCsm2DhgDms5SOFKG2BKp43En+cHWxZhBN0SJq6NS9o5p+QaULAoy9sZ
Bf8TltE2ApzZw1c3VxY1c7Tly4Yl7imVDTZLNxFzMkDrtLWpIFdniLo0SWcdcAPl
WzJYKsm0mU8qqM3T3bF+l9lvjJ7YugqYVN3WzZJLVjkql9/Yyu6mgvD3noiQ0peA
Dv8B9rXNRUSpaXRvt3XZdcagYaXjbZFY5sAhid0ZDwIqT+cZYmqZtL5GP5Y6Ks5e
cZRpSQNzut8aEBT8GjTpKE6/GJv9uh/FiquIGHgkKW+NhaFF4P3sNlcZdyhuRNN2
rJszZqlqdG1DS0lXDI7/UKCb1XBT/1ANKCeZWhmVNOgOAMYkJsl3zGIutZtf0P5U
MLAHpbyYRURLFiok61N+GjCqtwO/92UsV3pdaXY65V8g8AIg7OQoBRqs20qPAvzJ
I2mqnNgfQSv8+nHkDQtyXfzZbKWTnYInwggoBavUakEy1qttpqdecL8YFaG8522u
fVqJVVXVVREKwVifRkf85w==
`pragma protect end_protected
