`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BhCiusdJba/2vDNrFecd+Gtsz/cqtlq6mMk2PANSgiPvJ7CkWP3phNFDIacEHlS4
PzVHK1sitpZeZe6UBdQ4wxOoaMZqwEENZGl8cv5gh5hKvRnCG2+1ULmExxzECneD
u/BTQSHUSmYi/cDMEL4RwMnBlZsm+SqltdL9z6IcSaI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17968)
URcQRH7yo0clx+D+SuYFJwQq08bhUz+JG9cnlGgKDT3JCkRhL6GdeijWKAw9PFKk
9qhzv31bPXXjBkzIreyTxrylZWKU+4M6YRlxONAm5lIYT8Mt8kntjhSv+ezMg0Wt
HDUvhUOAskHFUFLaHoyTH8zX/5zjJnduhAr5dOicctM0aTsIaqczeQRQkkdY/2cy
UGa96edhcXCH2mfCbLI7ZWCcKBzDGu7DPj+tFTtKUzCEUHKktvY0OCKZRr6Rlr3F
fTpJDZs7VD2jUC4iotNxftDTtYgQBDL0BIBiVvTAHeEdq3jeTJfpmQKpcHF7TRPM
RwBc4TNSoKXNGs/IgaKScPJoY/NgAM2O7BGS2i/d1SDpY7mN8sph3+NKo4LCcDqj
1avBBoj86TmSkOZPaX4AsOPO8eDpmjdWJvwKWOLHmDCypnDeqZ/GxFBeitBWbZlD
JnjqDxqdJFzsoRno0gNEH2n8Zz/Z2Mmk8wwirh8bAYnmJGWBU7gTTeeHgbBbvURl
tqM1yrDwwmyiZR8cwapOg0VtLYsE9iZMbvHyIgY0D2ZK8CBeOn4egWpb/J9hTFXk
IaOFudeoiLJiR/g6ctpLzh6Q4Uys4UXGkn4CgtxLWGFbmEc2Qevjty0tdn45Vf2s
sNyBQwZ7751gFHFTYfllyoeWEiA6c2SPMRF4fX0y9ZlZ8DLF3WkD8iGMAdF2s/TC
mLmTYlQBkiHhViC3KQj5v/8uWXhUvy6wOIc6QlY0uoKy3oR+9+SmLZNOHoxeYGo+
GD8w5GgX52akf+mD3RNTPkzSvh+CWq8fuGlOnQCIHpUZzuZ79ZcVhYlOeM68kmx5
Qi+cgj3RwK0fGbCAb1XiJQae51pei201i9tgVE36pawsgrqF8N4eXX3wG0NYD7sw
vZ9VGdxltb52Y13YaSz9OJLX2i1nPNNUynwO5XxblpfCBcIrSszERzuQ1ltfWVq0
PyP1y2VF7T4Fxt/sduvg28/ZVxXHe72M44KujPEyq/aN1lZCv3+7+bpXQo/Ktgb3
fOVlQRYsE2/gwXKTtOECe7Ky0voZ6lCDK1NQs2f9Wx5rbEecYhrXJ0ciw5G6q7LL
HDVycMAw65glqxSAM98qbtmcGrI20wgA4J92FgjBE9R9wU6JzvOFwcZRmESbloOJ
2GFDBcXWt3ZuBoilIrKGTnD6b+cuyuUE02+GIdgWxKwdAUIsAjWPvbx9amATlcFX
QuISye44Cj9AVNLosULbxJc7azUWDjMud9/D2UFS0RlB1hzHYelSsNlxLUTcXgKo
aJ/O6LMGvzTgug0BjDfkKckSu3qWOw4c0yTA9Hyh8rDCzDTBDgYTVN4/iqXQgIcM
I4c5mNjjkzGK+Jodggm1SuQEu+PI7w2c6xq4TaAUnPNVpyBZKmxcZFrHHBqN5dcI
e+unlS0U1BLqybqfmEm74LfIJb0hx+bz67R6A5VI8mShu3hPnl0sAI64n3g50fY2
yg/kFy/O0ft6nfbyEiHlE2l1Qxn4R3UN+p3C+UykiGUzmaxxDndUQxxeilPuPLhW
wviYFjr+LF2BACWe5Ok8jFc0HijskZK/E8GKEZbwbiC4rHjGMtmsGiKa/3MR0vMj
xzSIODi2WmWpOeKtGWL6eeeJvSJ2MuSsHzeUDN46SJatwZEx4yWJujgrdRuCiXhl
3MBLbx/EwSnkSh8plWXrvpakOiIVUHwtJR76J80V3EhbTJ8pCraWQO+I34Gtf9zl
d+8wF/myYs8GULsJu5/Xo3ZSbipkXvfUuKmlQF4zWPquAfEcn+vL1aLUs5+CEoO6
Utw82ZyjBamkkDlX10TiyUPiIpyRwCXqD9Cx3V9mExkAxAaBsoAQLG1a/3qSOcT7
tuKoi4phqaljtmq8/BvRNfpLhy04IMbk70MoAay5MVUMeU6AlmzDAMwpcLjTglV3
k5pNzyDgguebu1ECxYrcLYi1fvJ03msAEdLz4JeyHLLETAwruiAU3BEfTGpA61++
5dMyFyAJ/ifoNlZhxU+n5GfOwYovi9H2JiAlLsUx+ZLpBqOk1z00ISgT+NcGocqD
I9f9K+ERPPZRuO4zcarhzw0vkHKZ4HRAKqu8tzZ7nukg47jNoK4TJVE09ubFcC5Y
CctHGweI7wHkZB422Ud4WD966822o1ZLXTHoEaevyhGiZ+6ieu3MuOOBFVIyWjuW
GYyo9Vz4wVCknl3cV1Do6THC2i+Uew380io4XaN/4SjFZiebZUT/3oWq1CwFyynI
pX/Sg1n6i88GE++DHqW16+Iw1npRXfF3SuteFeJjSHMzrkm97IHlRNE63EOv1DK0
g+x23+P6IeAgOyHgUO+QCvEBh/+YtC9aqHodRuzCySV4N0q2FjL/6qILPraudtx7
EUt8KeXwN7+u/AcEwww7vAV9KhPwCe5CZQGOgfm07oPFQ5wjpMpR+FLdSMWIa6+B
surLdLZ2vj9ZPDYLXclqxKigDiuqXwcSYQIJrmO50QWcE7YzihP7IW4H3lht8wwg
4uRRfVbGQvO4H/f2+LuQ6G1ahzOxCKpSYP6TlFoPib4Y3zIhZ5nxmUxiuev9ZOY7
omDD6yqF48JT738g7AWwY7f/RBjq0x9vg9/ey6Oe7YbllFT3+PYEsZyU7MzFzUu9
HftI9nIQhOfjzcHpgTClcGaAUtLzuVQ6nYc6tRfDRlwhDQRM+5ehJNzn4SEqYGHR
9J6JWoBcJSSQD4GCyDZwux4c6R5DQvVdOVUcIh49OuKQy7nCSMQuRXoG/n6VDnBr
O03Q2LyUcn7uZDif1aHCIwAxs6vFAQ36VFRTZXNkVyEbKdRJ2ond33PbdXhz/yC7
Jaormng5VWTBpo150uiFekmFQUmx+jqdYtNYmxa5p/Lig4MRM5wW3NVJT6Ysgobo
Jih8GZbl5hXzk7JLDzrRf0nDgwsgFjwj2rEZIROfY6aLndHkehwzXblQHZ2utyKf
rJlUAdwwnr1EniYMPzlgE5AT51ipa0f2TXRHiUTvoaq16/jlRg294cf76DPf8cJD
t2IGrPnIQCNVFA2CsGrsibJfCBFNysDX6AikWtObzBNQkj6qz70hInA44SyUsmvC
nBH2vcFo/A54BUT/He8dZ6+dKlB+sja6vOuEv2f3wloduWT8mhUefUcDyxs5h/UY
plRXiZ9zp8/3OFtdYV6CfSCa8h2Q9H0i9Iv3H+sjY8r4lXa8AIQm6oalV7Pl0umc
zEXX16PVwoHk2DU8Ey4QGFcVxMJnlTIn9eITfP7DvS0JRSXSr76MhTYV11K8H2Xa
SKtfrRC3aR//iMWjesXbMay8KV06/FXwlurm1yNIU93TJWbjKL7fm3MlO6rfn1B+
yCtaE0/G75dFx/CVMiwpiS4c8YHvVR78veWyzBAeUHTA3Q8phEyLQJY0EUshLEnx
NliIG6JNGfD9ixeeP5yoHdYO+S25Wu4SjLj7APxi32xiShk+pIyfYLfjESpWhDpc
d52sH2qfid+7Mk8QdaBLZOfbB04Ovn6SpzptC8lc1HGiEY1m6Sib2vEA6stOOqIq
bsBfzxf5CXE5KJZtH4wasY8nNe13B/IMgc0ATnAWAo0MtZ8IiG7w8CHRLuAeyvdN
xIzinsZQAduMO3lM+cHOUpYx6QP20IhxIAAKELICpToAKsYN2uFs8/J9pBgRX059
QwX2zyoQWq2CnFRTI2H81OIM8XZomDmu31xy635xN+mBuarggKz78dgeggTkt/9z
vEXFhXOwCjhaBH9+vrClNIXYE8x7hlFOuDwFRHLxAS60pVNQCVWD3cCCE4DXLo3O
8M/U+oVwGWGQIzKgtpMo6HH6NUvdE5l2k32fOjBD3euNA0rrZr89MBL0tdB0rN4o
P7V/BUBlxYt6uhtFWZrlaahHXtyRdN53MK2VV+PqxWiKMNxeJw5zyxdsBsXz3vVp
UJt3zreGk/G6AwsE6U7bCR46pj0PH2aHZFkbGgV0voepRfYFL7UiPbYY6pfjrwKe
qPRhavJ1eZLW0D/JcBxedokYbz+g7nXMoHf81rfjlso0vKZlGn+a2MXxhSQG1vwx
fi9RhyxGpzzMNrqbzL96eN86Okxe3lDcQUFE3MGsJOEFcuVNl2NphoUug4oHLV91
gmwREq09trLYWAgtfqg77eZ/C50w0fu30bqm4C8wgQtRWU96u8Wc+gjCC2G+g8sG
iexAJM61UfeWNLSXmbogkSAI+8anNYB/SK6QpJWHEVcXCHi9TIbPVxe2okaKTWVu
r7mGbW9cXDfJXK1kCUgHQhTmBXCSDXo23Zxcnw23vPGXnYavr9nLA+I54x3Pgmo9
NPkd+i1N1d9pwu8B7cb64ct7XqFoiIZdTPqV0NjUEIrWt9AV0ibVcAhMuow1uzlj
b7QGcTWzA97Zu1vQGNdJF4SDpuwKFgnIJrl08HPG7t62wiTxDb8LOrLREoO+vQ/Y
Nbji/4AEAW/iSXXbyR5umcK/eYzTajCTPdgh74zBeH6QDY7NFP+rvg1XdWUV+mNn
gyNxpyyxLNB084WLeyCbedKGRtMsmJvdSIkeoPMQ4ey6zQPSyyfhtNOQGcuvCZKJ
4d3lEkgw9E7dYBBm1mN1wgFyjOMQMWYVrpYHBawSLgz2HkxVZ5cPXaUWpZ4h1Zqp
MAeMVPsF8alx2Zk9AD3myphNjjfRDi4459nlyfn+4Dz/tp0PdzX0MJtoyDubNMG9
oZgRGANu4NloJbMrQqnOH0ZSKjxKgepb7o9k6dV0/wLGZWCI/gGLbFGWDbreArJ0
+XV+xNr00C86QvD2fkVK7osyVWYsX3T3x+2XSp4sXPHvx94Dvy5ONp5TkSLtSTK0
qAZ09VrgSsoNtww3th+gOwon+bqP6LMy4Tai19eoSQrpsQNfhM+ew+c4PCtodSTj
gcnub6i4IBceFvb7jybPLULO8HKeJE58ehscfcN+rykDfVrM/U266NVPhfyE5itM
GIPUqzP5q1FSSoqM3w5G/o2JbuniSQ/G+1vBD0TYdjwC5yP93yDibvXWtXyghxTa
QlrMLTBoheFFGx9e3vZALeIs+cuNdQH4GwGae4ObUAnhwlncAC7ztyO8L1/2YZwI
fg5CQ+SYKLhi6Rtcbz/2z8dXDrq4MjTA4ueScY1667GR27kfp9PxNtwlU+TG56vD
7Z8quEQ2/5unGOamxFNTWZFmksXebOW6//4JOiaavWPmJZWSZXRmR/vzfRAbg+tC
p1uUi90JPN0zS+qKW/3yH2gdFL/0x+12Kf25LCdQszN9bpRPZleBrzFXJuRtNwoc
43jrbCLF71m/qVSCdL8SQkI3/KVdBHuuvixtan5JMXEFwHg/VkTYm2SML8OIqASl
YWZK37vK1swc7WKVC3opsiTQOdEhM891ERiGgw1luLm89rOtit2hPp4BItVdkVWr
Gn4upIoHHJ8uVV0y5GKJ0QyXEihWGgAG8qLcrWiCxlSxJFfER/+QrO1yH91Vzi5v
vDMxPf1lH5k7IxIAgIuok6FYAij/cMPbq++q/ZxBfw0ppUqS0T5pNGmEq71NoVeM
DsoKEAuNbRkm+TQX6a119vCaI3WkiExPOh6YKuyQwSw+P8O2weKFt3avXlW/bl37
VOKJ5OpondPbj7mqJhzzOnfsqLk0KQgGW1yJNdW2QLr6OrnIPdoSzuzmdks8eJIY
/6HOXrVPxOgTStcLmaOPd/kpRiu/GiMCTFPrCIH7W92Rp+dbIeiLrF8YsFmM03w8
spjqdMkkESHA1l8sikQZUm4D8XOfoaJyTpKGolTpwKYP87Qb/tlUuFZ2dJ9GvxiB
WVNQ9pvXjpmTC8E+jofQUHbwNdltpq+NMJ+xTzj0vrF8UPnTy5CK2FIh1UOvPScb
Pao3HJyqAC9sHJD7rAySx+VeK53ceOz5XpsCAHKHQwBUUuBTve9de+RUrEol0ur2
W8hL9WvmYoCBUpWIhTvU94VakQBCMpnmAgCbf0Mc8JEgnTt7RpxQNau+FKMJP8Tz
DrTWBXmoh/oMYZmdSM2bLsDHTAvUW1sPm/tyfizuphZKcUqUBR3Ubza2YMqwN+W5
Lw+E9Eo1JxwwczU5cUw3F92cSRh36UXCqjMbWPWCdOqpQJUj2cz4cldEjOuo+unC
J9vHT2Rc9Zas9lyvG9RJCx6s8MgTZ2VOeWMI36ezdWG/E216U7oQ+ODVDHPYGnrk
7dBSIG6jZPlEweUp/bXYQFXa175Y3B6UIeJxi8XCGxR3xqzzbNNnPFfrECc9F1+x
rvcrNCYHr1MImO2t005cqXjkrwfKhGG0N2Rjqlxakc1lZ2tfPHcwXS4J8wkM29Wf
R26YBz1b56u3BJxfUq1ubJ/VRgFOmDxtNXeUpWE6qodb8mzmQHk8ChYSqNr0kqwM
9C9GcCEQ4O2YfCf6Qup9VIDbdnbUSFpj0Feryrgpt9xCWcF/eQCVuwtAsc45i79T
MCTlPaCADG7dRI9rJPfZKGT+84ChrRdDpkJrogNo5tZHAVtE527R9vZel33FSPOn
eBAhzrwWt7RjJHQ5Hj8usAofh6XuDweqyd1Ok1BdTB3EymKIG8PNwPp0TgG/EFQa
V5VrRJLwYxuUWBB/wU7IcKzSzwC6AF9oqMaDDsCSUxfivYSWW9aitqzEaqSYiWqC
52rdtCktTqujUMT8P+OiCWHHfEuBgnBVXev5wjOn8ooAJzKAmDNmzFXubcdmxePf
LbQNfs/gUvpur48VvIZEtHKcPt1vvDIjNYzgioNh8kV6RZn371vD65h7EndCwzDC
pH06cJzi9BMuQB3y6FW/mlqbTIBTxvUEiYmK7HIfdLJflTAFhpbcitLsvJVju4/Q
+YT85ew1BzTl2OTGmci9K2SP+PjfMGgJ34R/kDg/DA6Gryf6f+mpUmuU1BxnISg1
k4bdIumE7yy/p3liuI0pg40U54I5ucA0G9ZfLLIilSto1kuDnvtGYN4e02rzDvwl
OdDuWINlx8xmJDbrYYhKEN+vol+Gk32mwO5BWnAGj8iz150q+RgtWy/yQOvOwsPK
YZ1be67LAvRf13JUuWfBWiHh2BufuLvKIKYy6d4pRwEEJTREzf/wZAp6Mv2gE9M4
+Ku3iPciiwhkwndXaf0m90aKu8c/8EWkD9Eq2Fa5A81nQDZ9jbBB7BLLQ8Zwv12X
evaqIZ8J4mevItpAslqnSblJ9fAc7S660jULvXlXMSHhgmQwKQ47CLoHhI/6rdAM
JK4dbygnUC5iM/QrfkYyLKulzLW9J2Y2ZC3IAXD16/wMqYwrJ024S303EpDgYcVW
CQnwqk64U0WHM1Owt82w3USBxLFWdvVPh3tY0JpUBY+42MZ8G1cBEfKWCi6uOoC8
+t+7zdc0wo/qjii/+Le0Q+twf37yPq4Xz0a3z7xy/H1SvQTTvweDnChkK3Q5hEO2
uQM+3JD2gO+HcOvcxdeMFl1vr4WopOzUrkjDo46S6wjCm3cQkF68kdJXEl1DtmHX
AtGTzjgG1oXMBZhva05o0nP2Cc6QnFNgB7zhk8roT5/fx120R+i0Rp/dG4w6a/uX
CbahzRzPBvoOqjGAzwFlj2NxCUcutJSJ3Vpaa60F0nd7l3wUVUfQltk1FNvXnJWM
QkFQ0TAgfTqQL8QnJ9XFdoyicwNhLbkRQyp5TO8d1hOomsGJc4LDS6D/ny8VS/uM
Ap9n7SOEXGyTewwdfPjDdpjUeyLEoqltS53J29iaXBqGpWxVxyhccMALN612loZT
PGc3I88NkcLsvB1DEitmdKSpl6CS58hHpbkDCIjgl1ilcFudNrT63F71TPvAX7E9
lz7lLipwiLEklOAAdAVbZB0l4eR9erg+5PwAPhMX6wl/PwPH3TgeaNJdGH76J5WT
gBU6tqO27GmxQgfJt37VxA09TWtVCvwgUCGoz5Wm3opQKIk7wh+r3E8vLY7lVOYq
nIojttm0n/099L12SFJuoYDdnxBVSYYfGDVtqs8gYD8jMFdiA8+FGLLjJS1EoQOI
5A5Ki9ZnNM0aS0HDeUL44aKX6Vl+CF04ctrFpIbA/FsYBWiB7xkheqU5KGqnGyCY
ZiFxyyX+byXAjm6UxmhqcbeB/QwgS5qpFjaVKDANsALxQmmxie7ED7e9ZZvtKoIy
nQ71uBSp/ax4US8OGHFNo7+Cy7lwBrRUKE976PVYrYvaYALyk5m/XUWqEqoY42ph
cRVPQp8ze6mFFs/E8DwtlHgRWcknMiQdxsbtKnOghXpelDFT7siXrffadpu29br+
g4F7VjgP8phZs2MNHlPL5Sw6JZU39nlq+ctI/jLiHNttwduaI5hDAu3ZpykRJqMj
sdwFWEPyPF0T7a6UYaIQAlQWlT29zr+kiGrsY8OIzGT0+m/no5hDKUF1x0Q8a7bb
u/HV3zhTFF+bZ/z9vVloQAw8n/jb63XTbaAWdALsRlG/QrvjqIqpCM57gilR59cA
cYU+iPI4xlyXFc/rzJEuN9QSH9vTS3y1yFvqMXypHPTwFoh37VpB+hZF8ieJO8Yv
0N8GFIqHfeo12dgeWvSwylPW1HrASJlMLqAkY7kmOGnN4QwZR0deuG9EvxfRY+P/
DMTU6YKm8iuHd/e3Yi9/zXZcvmwLeIxJSMqy0YsvXmViJH81o1HaUQW6wg4T4d6X
DzBDguGCJuDEn2+Terx7RcI/BeJX8AO6G9ZWe0ka+1kbDr48NdAs3NyIljIbUT2m
gDVKktWNnR1yIrEH3l6vSa77BENMIt3E+xNTaUm34tVE4PHueKYzH5Wt/MAIuMyU
oVhjLoFqyyDO+KfbMxvqhUWe/nfp0V4ZmnD8q+NU7J9dwIvIkwcBD14vBSeQDroX
xKnSCUSwrTogQiDxBG1iuFIEUPF55UPJPmsm/syX843xYVqwsWI8Eta0nK3AUWgP
Qex+K/0veWCEqzDnJMMxpQDWFYiLu03dNyoElD2QgpOEC8A7bz0Tb/ovKCqrc2/E
C3nw4AcSEoZPUiCiZAj77EzjH4i6meY3c9XqQf7Y/7kmO8pQ/PHrUCZtFJk3K1bI
C+Yt/6CwFcqhaVsvB2RFtzzSnqGr/GWm58mdBkFnU55aXWnr2BzaOvgMoqAnqbc0
hyHv78VjFrqG2PFFox2OyZUlOiyURG74Eer4C6fETAzJYtJfPMCUVdsPsf5cz7Ir
lVUAlRWQW4eSj0HRUMIqkZ+jHybnw77GHGwfce8SuSvicMExPqPU/Jrn33xDCQ5N
MCG9Pv80lQOiIC6+o0lQph+QdLwf+uVsb5u1GBwBE3m8CX5G/mxqUCVSwxevxjkR
2EPaRJWcw7Yeatkg5dZ2PZIajDMAlPpJFn66w6+nlhlFKtzzyavBF/ahD4wngRcV
OBW8yHC2EJEIDiQxyhH2mXp7iXB1Bd8jkE1bDivPNzYkCnmI5BubCMs4TCV3+ElN
Zv4SELo7olCvN6GfSR1AS90Zxb6QW+ahUEsKfWl5Jnopv2cfYxM3Cg6Pr7bXLScE
ut0YVVBHeEhKiAUHAIBSfNSdT9rXGnrR/0AczbOIQnuWSKOcL/GEKSRaL+rsjV67
W4KC7bNtrx3KC/KUkSXt2PmA2fDvnDaekB7Fsii+0XrWNNqzCzc3JUdClTHmP8XU
OnjhTS6aKyFhbRQviWBB5gfoEgcy5fg72amZGbp9qy04RL98suWLxeDSUyXKzCf6
YL++WcuUG1ap1Mrr6cPheCSnzZfx1YDBxVMam3Y8rLEJBWDzIVt+4i4i2fhfeIqj
EscG64PHr4nirheQD540IqSMf/g65S0IJc2FPvFZ+5xQN+Q6MoaZnfCdGBdFi7lC
gxdHUzvGQLEezZgiIwklpdU4FgI1ZxWUT1ryEL2v874ciZ4PLC21V0192l+P0qor
vNCUIY6iheWCtbwbtaVE2mWAyNJDpwdEDOjWEkQnH91IcztNETCzRRCB2A0iNmQn
838jY0nlgnpGIXK/TadeAyOwtwP5rb/ffa0cEeuOhdUsPR6QEfaPSeDFT32qzUE0
7HPtplUf5xnIpQN2yrU+0N2kIMuOqoT4/vTOo81f/KhpWpqEsn+BXAFcwa6+Gh69
p7eW48HVd7qqKz96h95pQPye5UrJXlmeYTLAuNGy9dNIaRn9zDCSLIsyxNeY9pZ9
eD+RN03My9/eN+sJTz+qKe4XwFnrBHf8X3tJ2LXtelb5SaKauOkxOz4DM/wqogJB
yimbLD4NrUQIEIcrjGvwZkJpPXhCEv7lHXwtpOaWPJJmTcWds76TyOzs6kcSXeCF
TzpczxbUtpRGW4NAXfu/bDveDom0vif3TlWew1qIJU5DTvdp5nvyPBcmD0Mabw/A
HtdDt2c7OssO3IxYSqQtay/h/HOPOgfGax1A/tQhv6cTSDIctrJgV5eDSFFiKKrD
hggvX9rG6kIZL5wTTsGsHD+N9vlhAdI8dAEOtsnRAuy0M/Jqnmyi2CQktM1Weywy
/IyiGl0RwetshOiUiBjNAwACVR38sEfBDR2HEWJyQa1ro4dbzwAiEe8W2iK0vW7L
LACAGz1OiK5Ik6NjwpYmXkhZ452mvOOxPcdf3mawO8veDGR9SmLT+rqANgf1u6z0
TMkjzSpmo4Z35+VBiDl0FAeJKhujMyEh2bSRW+0EskqEkE6PDgmShRIWG7P/zSq+
eHNOvnPg2l1O5erpwkpWOOeHSO7WB0h088zd50SX6iUo/4cdm9PEXItK6ftP7zfI
KiMgVmHAK6KzQd83CBWdpxQzUUDbYdGVBdJO3MaHmLy9+rhL+BRk9T3ZqnRBlQp+
EZ+hVWDzwS8e4ax30m7Ex6KTi2IW7o7yZDsp+8lf0XQvix6zMmtWyJ/6e27uFRfq
3wJDZsi0zcmlsejfEsNLlyWpMrcjQel6tpSOTAHFUiQThWn4QWhx7YlQFpFYLsW7
flFrfZm7l9pmnm1F3TUn0tuRGjIZJvt155Afz394PtmcIYjG+jrsIcHogtoz8B31
0vQ+dg+AN8yJJ8J0bCkxCE4PTS3Bzu7nRB0xvcrxal2NShYQSNHl8vBDJmlId2Wd
VYcPH47o3T5N+LMnHlaGqP8gYBi8pwhOTjGkAp4tEjb44GX6t3rHk7AxzKk7k2Bo
bNhv+NrskQavu2oZTAm/iINv0w1hrXzpoxZZUGucohfkinZZlcuFp4ER2Cynyq28
XKkQfzcYN91k4IvKKhNGvtJBI9Q9jWr5pgx/FLZd2zcPTi5A1XpsfnoXZkIDOFvD
U5zfrpuY2qDcJPhy4UFeUJHZcvcooTsZPIwipzLFntDqISmkm6TPpekihinwad6+
xpdcJJajhtQ3qK1mtR897aWC31S8ulxP4FOm1jvNoVBrZZk66yu9u/KyPBCsJXx7
t8sSOJuKfgzU/LcRZo8zU7nTA6suR2T8M206N6g3D6T7/t2T5H1duSNXJODjQ6By
IQbeEH0LTLACkQRUGqGfCHFwv0JTQwyZYbLX2H9jjgBzSMOjbFINYFwpsEr/AzgC
nDkrQweRAfoRtA8fqNTdATIPnUtmPhpT0shQbs0wXaUDN1wiRonvNjIqDl1knsk3
29JLl8EcHFsG+bAxKHTDECbPKvM8fw54llEVGCI7rkPR204FUTzTJr5Wuebgf5Gc
Y+8v/wAuQZJyShuEJG/9nmDcMihxFs+ICWklS54pm+gaiBgcCaXsgZs4yOtm0uPB
JzooYLgGQtmnxXrb51h07tGxzYLRokEWQwq9OqAQI2eekAhKJ9Ln9QTV3exAlldD
IpJTT65B8DkEmiU+dDJC6xCQzqu/R6vJCk0EnmDfuN0lfTgumiluSjlTnPXx8RSU
rHG95cPynwmWJSA3w4I+gwl3s+DtwGCzdtljP6YiwJceLQCOpRKIvzU4Z+pnwMI4
x0SSqJ0JHPrJinlvYIt7ro8qfvz9jagpeCPbtbAheJ5ARSLaV1EPAun1b7Ph1HBr
scSsS2TLXpWsHmpGvrAILJo+HUzkwhzp/1VgtMk7NUzg88vV6KRQi6B3u9Fi5nvi
9T97AENqjBkKuR+q0nJX+HBfurihAV1RqhMEPw5/fbFJVmznh3QCpXW79C7OY9tS
gI7QXvNBece/ZIxfJD0XN7drjfeQEzUcgRUt7vRy7g9OFAFXLmeOeqiA8ZdITvL9
tPPFzeXPqtOlHXtG/RLW3Yke0S6OLFBkORoDH6ntttLrfROHKOWRBv+juDNxAZuY
FAPkBeGPUHgWcX5B30nGY7yx6z4n4MWvvPzKjv1Q9lci7c9ZBhQVSpsUarcrMb//
/Cwb1mWaxFQf/zy/nu4GhM3bBMdKi4um3gMMOTAQYCmOuuQrBK1jgn/eQCct14zv
SxGxPRE2EA4N20mKrF4E/hZUe33RP66SPzcI6sSXvljCxnBH1WL/pYjNtZxkA9f+
ucMRgzPSvDekp/fGvXHhMnmEsOfFaLxbwOf5PjgP6y+sljtjFBlCpRYTJAsDxZfS
d5kbLibw/QSQkyktjOZAZUz+NlJS2wDQyb05JHaV3XTyt9ByXRqM32K5UVmvdDi7
ndZW1XH5mXyv5P9G19WQwaBe1F6ZKf1EYR7/dbC+W1XuC8x6QoUf4DSM3qKLzTTe
hABHW9d4J5PvoTJVqAoKSExAL68AQGC1slypo6oBPK9oMrwuzLePibIOS01Zh6+T
8r9EEUEeC4n6SmgXWm32adLHhFMcsvZzWZbbjfChbNRu9MqTTEKkMRT8A9KbywWu
y2G07WFEGTfgZc51YNkujpO0M3NSqfSK4vGa8Av1Onu/Xsc6M/apK3WF4UF0oeyq
VhiNw26LU5BGb5Ay3UImHJ4DntmqAuZjkCVEjvI6hsfGYvOE8vS/HTpd3kpwNxtS
pTUUaRM79gAGIcbn2eAQ2Jj1S6WGRe7ETsLLMXCRDsQyFVqq6pVJfhatt4BrPiTe
zIKaQB87BP4qi5Q/Q8V+ExHm8qVBm0ZAHs9wSoq3acjjZfKiwRYhsWQGzlMgD3qR
Z4PrlHkJqPq/qC9gfgZq5lF2BG+pt+NgzCIL95LDdZIUwx4RJMaWFy1UJDTW3oVk
jC8AcMMPXB0vgx7wLxORn8/9wS4vz6XT9vbM0UQo3f/3rPqdZWYYtCtNphj6g/ro
Qk7kwOoEgf2T5fI08ehm/pAG4SQltnO/d+MhZZNteIqHO8TzHDElaiN3ENL3TCCp
1a9h5Fnd5h6zP1tes50rVjka4Rjjn4RJwPqd4sJ3fc9PFaF6pyGoAEl78s4oKY4o
fD8CqPEQoF0KDf3zuH/fyS4Ajnoa6V7PFaRhaEtb9jp0cIzdOfIzBjODI7sOzMIM
7RjiRG8HDiCE7UJIAZmS2HSlYnxhQ+PkYwxs+wPua8VU+SrnsSF+0lABCzVRYPcF
vK90yzIYu7pQ70T/LEfZ3tPSwihkTp7FqaEfmXdGT+GXDWUSuKUIXlUTGnh3hJIO
7iP9gcK4jCDV48lC2aAC9+o6rNMnyDiZdvFMwUzT3fGgFjcPJpM5rTQ0hiCFs69Q
KF8vdat8znpAkEw+gmNuwoo+N03VH0J4bYWjw16nAchLKATDKctQ+67NTD8to1hO
slSHqX0fKXe1iha7uqZ2LWH4JdbY4cOX6MuYyIUNwS+QN+UfW2FyMvsM9IQbiArH
g+DYYS/JbXEkNcsPIBtNsw1PqN2GqMLk61OgIElUaunwPFV0/uIaTF8xbdCc5M9s
zr9HUe6aMgMEcyv9G74yANKQkFSGxplDfVaZHJtSuUaiR16CKrb9kOuvQNRd3Ncw
2ZhdZfTXm4J4bTyeUh++3h2zLe0HXYfbrAqnktDiN86P/UvtJQNN+hfCI8xPwnp3
+foSWd9J/06VAbGXjQlYYJXdWtN89WYKaeE210sxa0G1KmrA6SJPF+EPzXKJ7ndx
dqbdRydwZultCSrJWQYMxI5VwGzw913BrxG0TVBD8O8H5LMKb3DWFKF/Y16nu/Tp
N+w5zgcVMb2KL8RMjoEojSSEnwUjaOlK50yG/5almIUn9oUFhajI/1A/zR9xB8ns
B/l2Z9O7bCZQeNBBm30Z0ByF+4vH8a0wiYRxQNz3Ie9w8ZN4xsaaifRWP37QUnml
q+7mwTYMz19Il5WQ48FwASP0mhLZy6ZWMZnqO8dirTAyohSN9tSaVTbLgGt8WkrO
MyxeGM9hy60kb0FcJVQlmNIDVB7CHaRCLLHfZ1Med5VirhliLGhKtYuTYhjC/M8e
cQtXxtNpSlLCDrj7h0vclehuyXL+wRo5fUSDa0dkZmxe3+lvke4Xfks+8KijNuKe
bHKgAuGeE8DeFlmJSDFaVUgAD/3qbh88xO6m3x9jaQkUEeGuSDCPmIDSB74shrAb
gb0hbj/HFskg5Gc9cpzlEACJNKewzp2cjU+yjTQ3e8ve/qhkASIp25/Pki25cy/P
NomT+lizny5FZJx2jEYHvJWhsBMFypxfoaIoZp72D4Le9hAr9YSrVSfSM78D/ocB
ray+7H2hSfTWSdDbaJb3yQQbdlHci+zdjW4tpDchdf1pjIgNn1A9yv2EbhSAuNdT
Do/2Vn+c80XWiczWogrd0sWVrJyKlWwfLLtNY3ELmF73SNS6STXLFBPMaNcoJGCt
z6i+j4MhAbVyxER8lBL/5+frnXY3p/GXafFEm6WGL0XU/unGPxs1nnm8cP/pIc59
DYRJK3IfJCou8hoCUvjWI4o+1xR0+TOyNZ8zXUbNjFR2VNIb/nuRH5TT3mg0TBKd
YIT9RGNE3isoc8ueC+KQnoZzSQzZHECIz0PyR9g1yy/bSTBF1oFVfVKx/kBmjH1v
410cibac0yzN4ZuQL0CH5tnP5dOKP8bfRt/BQGhLfwiVnmHqb/oda7QS1Js/Xbc1
yUtZZf5yVLdrACek47/Vs4Z5xI0qnSPTjfdzSoeFO3O0XcehYDJlKNmiyLz9Eakp
+PM+wBLdA1GpouURTRZq+M7RbxXYrhX5g23GLwInHFj6bvkOINPLAy2AmVUTMlaQ
1QaJ+oSL7Nxj6oux52kJkUmoO+ZwXecmkZp0h4Q/wJOyS5zOkYT5ofIizHihw8Gd
oT3sP51AnmCiK6wRRDZeU/gT/zG7flSWc+FzfwAZQq1R1BQUKVPNZEkSrGHWtAhK
FhQeHdHGhdXVxw7VO0SHtN2S2QxqMt2eJ7M0Xzkr3eqGmXoBHPW/sbz6iTk5bIZB
XNK/kKkh445Dzcxj97v21tSJAZAd9qqGIu4O/XmAEv8rvZK6Ney4q0MrtQFisgMI
yKwixTKsBUPeVZZHNRUP61eC4lkQiZkuusVbzNP3HfLTpIGiVu5ZyULxjjacMRkK
wkyRmj0XcNTxKCjFk9UtjaK3VFBoGMAneo8/UTKZg/wVLAwMYXjgpmYNL7+9xKhi
1+a/uZIrey49NwHnGhmWZVUQXJZjsEMcq5Zq+/t9iD9azrKnxdHUo1YZjwbh4X/a
gjN2Zu5/xGZcG+xAqhk5gL0uTulWKBAQSCNIJWFgtSoQR8u6JNzeKWz7ulZpb1vr
hb6yS94rj7Az/p/HUap0akakcHABFEwB8HQYUdqjhPyExYTEVTSPtEdZ+M0MDrTg
j37oU3AKb17BWjBGmBrdZ6TH7SVXpOf2/d/ig/HahHRwSt7NSH53vQgoA0sowVEJ
H0mcnCZY81LygLMvxw7ftVmRSkTRydPMothTaBlrJHtSlS/H9xbT8vIeGY0FsZza
8k0eZpt5sRbupnKKlOUEJdrjqr/hej0bvHc+Xtxg5m8us6dlPRyB5v9YYd1sOzoh
fKPXtnujs0jy/nCGt8orPFPV+AiWK3d6+xNY3jp7X0XttsFb2eum2sdZCKWFllDZ
TV2C9tqK5qzCLxijknb5MXDfpnvK1Uu6lHJvTabIC6+F5TRVejx65rIF4ZrNItUA
36BQGj9b3rmYPIrAnhvqdkOVTo1NZBBcrb7lcT/JaG40d2VeUOMz3T7evvqhGBgp
azpw80N9UBqv/sarnRbyxO0Hl0xYyjfLIB9CMLc7uUppGamraOW4DC13DsJeLhnk
KZ5qRGaL0Ns/du+enC5RFg5++Fka8DS5BnGA/9RERXntSFbSQHStvMBnoHVli9Oq
fzeFZlVCVQ8NaggFZDuDzgnCOyTw74oigNYMG5+NqkphzeFLLUWyv4IHC85At+Lg
JMu0oNUU36xGQyKiCOyhryRGENQeLeQ5vDuSGNtla7sBTSyr+NXhlmyJ7u/mr5tk
HjisJhrU33cxUVyFihRGLt1DSycxNzcW7ouGvjjlQvxUc+7jf+CwP3BTQS9grLK3
ZFK6ZiVcJfdKZNa79THX0fGNT0IwTT5gS0ZDAWT1mzh1PAAJezm8rx3pDmAS7Wyv
A0SD2P/Alg/j3Pm2aI7thCk5pdiMUGjwynSs3zn5aCaJxLc3qJTALx/LDkTjQ3qV
SHFVHIdwT9myW5yn62DTY5/GYZnYlfhmKbQyg1CgGaWtjHSHZg1vYfLqlBQPbPEI
Or7bGBrMKU9qWXOQ6zk1PhfLAxIPcou7jOJblvc5n3AhUhXNeezqMkghJ6Juw0Tj
nd2P/PkR5tofL0I4ErFPAZcHSM84FlSBI08J09wD16/axmjDkld4KnjrKR5KGhNl
hZa9xY3akLGTSeggk2re7sUkg/V/6eqmNS9Hb1zQqBi34+LnBPWOAluG76hOdrUP
gAXYWQT068jUUxnsFcddkFfL3LXAxsZpcYA6FFYaEOhwRlA/NE+7qIAngPjEcSJJ
88mOvboe1iVGQMZVAf3XadyekWPQV8ScfRQHTa9FiJJFqJL0HONyB0ADwxfKiVBU
LY9qd6cvio2BBKtRxZrc2FXfaF+i2CRHQ/hV39rUiSNbA66rjTe2jfMJHgkcw5l7
X1Ii/TeeTphGb1be3WXFsJfWeK332xUgwjkoCrkB37QOAmQUpl2WCHH69lgBEwlK
TMvuL65tdclds+x6vuHjbZKTu/ViuAZMPdyL/hTab+2Gzjk/grJ0yVgg7E0Igb3o
qL9FKJwHgk4b41lMSDR6m/yPXQbm27dHOBU4VsCixlV603Iycb+8DqgsPA/Eqdfe
C8Mr8j9NvzJ6105lgpvWPCT+2/JlG7DBAD3jBRnco37FamPM5DRgewq1P+Fhdbfn
shdHII2nXfZy0+/8NmlzjhFjvmK757N752UZgO3OZya6l0DP2EOusBJqJZ0qpNOd
q27TWdSV33uKB0ynFN0OGgwS5iGjphZf7Ml/8WGwDlUhn+QR/67zxLrxJ6AFj843
B3oaCc+rRgvuFmGRJpqgl/77AwLr12fUawFycTk0enfov5pw/9FQXfpG+2+dw1hw
ad5i/uFG9DJLA0HrsnvzK8JwGyzOlVqURBJ67xnMLpGNxxcGmvVEwp6D9kYEMl19
wiBmp5j86lEDLK3JeFmpcqE2x4kfP8o3nhw0Do45Q293zHCVC2x89R2fo+xqfO9K
1hPCM+RPgaZbB5RTjYuOEqqvil/cxIjjPOF/HFA+aILY0quS8QVblX/eeJElSFCO
b1/VYYoY2MtdJOb/Jbiw5jN4g84DoZyINjJG2Q2vZOPsMJzJb2GQevcpTuw4U59a
Bc6a+jKnyHKWUyOzdE3vSCcMJJ3d8txD9pycaI6FNaEwM1OglWJpdy7/Qy0UXMvB
o3EBSKEtK9k3Q8OyILG3LB6dEPqstHiQVD8j6QkmPwMhoxBLiFltoEm/R538KxW+
JP+bwlNTm0o/lWAS5CnF2nWgk57A/J376c8wLEYWp6c5RotKFdvsmg560p4wVPdu
9+3dvjCuXpM4bptmyyEWezcgWJ9Gvb6V1kk5SXesA2S/N4WnIEo9T8cREI2LL77Q
bfKjRGd+BCLt3R3ASKOkD8cMQsGWAnHOFDZZ3nOb6pfH9w0jLas4D8p4ez1X6Zh5
ImkFBw6wmZNTDENVPliJLfcJqfqxY33/cMwQ+o0kZI/96oltK7zl6SL6eg9F2U/E
+rPPU5mmXn9IRh4amaI4RtmQZI9XLb1JiJuo+DUBi0pzFgsC4vWtOzxNSEd0tbVP
bUFvNih4WFJ8fePe5wD7pxUgIs+UMe9PuFBstxWqMoyq1RL5zeFojDFRAkTyW7Rf
f05vF4cn9rSmuXduTz/a7YZFUlH9uBRxW/rd2OtnDaVgPuUP6ANJjuGGrThHw5sV
fFfMZcS78gehu3H1aIfgdcGdgF1SEP9wMgyl00axdbMcNh+o+WLXhUHF90j+VO83
jTclPe5dnk/x1MkFg33x+di/8SL09llValWWSsedJ9wrwQt8npw0ZzWwDFFN/54u
rKQUyR7jbznrauX4ortVCiwgC1+mo9gKY+yBv8zTpLZTJX2qn/5o11uBCzFnd1Xk
SVPUKoDUu5ad+KWufbWATVuqcqhsKFSglu/4fcELXD4iaM+8nORWV/XMospcXvvu
8k620S4BMhOQPjr/DHLHdbnfNY0fy0QL3pQD5/a7NxBKAY+X5n1EL6OWpb/ZXALw
RsusIncnFEa6BZlIWBn0DGZeR56xanCx0N16uC54MFYXmThcOAH4p5LJRVu8rmaq
y3Cj8VrJ3Qc6yRYSC/8VWdRWzeAX2vKImwsPQxUNOUK1YbTXnQjlRNn3o8X2Z3ou
OQz6KEWU5KdVxVY1rDWcJdBRCsDXMXjBzQDSZGoTjCVhbMMHhHQ2iDFydPfsa6s7
6BC2xFXYeL6qonA1hOBexzYi3yGADr5pBCDRGXK+1nAHT9nTRtu99ykrVJMjHpl5
3Ztv440V/el6WD2kyd/R3x7TC2rqrsz1aSmAznM0en/4yc5bipuFZsQd5fO2E/9D
4BoYAH9KMN8TC8di0aMdfRpDW0Z6bxMnS6T5k+7IpVVdPssPRh0KLecBwCke2kxj
U+W43qKZUjbawldsos54AP1qzdGkeNakiJs6Rp2O1xXC+RnGidSfZhFkSsam3/4R
FUNd86iWrJ+ANZUn3FddkiCrel0tjeETRpfP1hj7kKrL3lBVqYLw05bnMzj6aCfJ
2l1wdAraXEc8gOzMGhdhtNaEB8x8UbErj9n9j7iLNNm5NIf+Mu6drl8VoaUf1tmI
Aw4spRHoQId+fPtQ6be5eQXfu9uqYMpUeljgX/cgiRpSVNktLn3BXeOgcOYtsuOx
uudHGAzWBFUq18H/qdwGmKZM9fiIalE3NbTLP+2kA5hgy/Sgf4hwBw8FCIA4h4Te
50qqVR/AvF9/leRsW5+Pgdcx+NVd4WYdeV8RbQiLCb9tFK5JE/07wgp2JZ3DFlSc
M6LsrLzTrCe+jvgV8ytztUcWQuM3ClBwL0MAcXIm/Btk/vdgEXCtMWuRinqab3tz
2lr2OqLV1tEEtYfnycg1cRhum+ZQ0hD4MArHuekVME/FtJGZpQhkqG7lCY2130QK
KTGqulFRLxbQZUbYUcY1iE5hsRJfj4e2lUSkCd7tCfTF6LifIuUJ53CeihYK6dcq
PB7iK6huLt00cRqVuIj2G5yDRyyTVwy85sRFvCLLOxGBgyYw/qzeGoJCmCAO1vpI
YhCAzNvw3U13qmesA49yPrvtQ/o/bSaPrTGc6KMIHp/UxKf3deL30kv+b8HsArsH
Z4TjnZUQC5Pvl0usyCVamiGP+z0Dl4GrMyEGkQu3DfriGkGFiWGm3b7yF+LfSEJ/
70o0FUeqQYhnggh7VFVHe8TEkRxtrDK3/YpveQ5nlpdyJkZ2p+zrW3yrwB3UAKZc
Ot3tESPh46rVw1QAAHCpcJwEs4SNmLFVa3dIWtiYMCMXeXXn/0t/5R+nwZTdFxYA
aM4EvXdD6boUdxzKVrz2XbqPlOIZtfmgIlmD5b3MJcshtN5vcqyhVZryKUOFFnNW
9um6RlTgaQuhU+HiFsuSy1yr0Mf7FL5w4XJPBsilvhpUqofh+R07MuIHsnBACyP5
9+EuL5XEOF1JN8azVWGVi8icjD7eJ6593EymqkW+y5Sh6oLWMzORlBkx+CFybQE8
4frZvDA51VFFbLN/ukJDT8SzJ4ghKngb5esiKeR3vi3mzy7FJv1eKG9B4k/Sx10z
RdrbvqRQuLBvwrCTYxlNnNE2D6xSCqf1MnZhYEx4kLmcFRUTmlhe5h1XcnwMlXe2
8w4FZk+CCO9xmNt5sPyDUShie8v+VARpxUQ8DkYrSApSj2qABk6Fi4T5TTkFs2pU
iOecp8sQYcdg+uLgREmTyLv4FqgJoSeA9+a92RN88vpAXQ7nNtDu195On6cpZ/5I
yKdcQYVl67+KnH8masTT6lofukZJrTyGLhpSUnQUivReYYLav/DOaaCXDKNlHOqx
G+W3/Y3ctbElMzPCKYw/du7HpgyjNVmQbPWr+R79wWyAi2xg+HuVNDAg9eR7QyNI
kxx6NlpgckHoLYHA/rpXjr97QqP94bV7egUOz7QO2GU0OzG6kWnHPAARc8vo+zCb
SPqhG8Ulsqdrzqp8xATkEflYirCmyTG8QtqR/N6gUC7SQt4Bc22RL1sqOXXL5UZQ
Sptc/nbg0GdqmcQNDZ0IOFyPBgoLGq4o6vmMOG4mrErDS0Bn5Z8p16l1Aw57FJjO
rUzDYUv2T4lSni1BdwFkaz4JTD2fCM8ogqZmn84AqQPRhcTV62yjA4YiOkguHLoE
JGtKuhESR9PoECWHkNfw7BAQOScHV7fpF0mXG9dd1MF+RsuuIWlRA2qvbckDmO0d
oUccDsY2FnmDlbRy0ShkoqHucHO8cx4/PDMfiES+/WJJ5C8xYwu1dms7tSykpeYt
OJxTcIaA6Iimz/7MUPJW/avQVzUgaMfrSde3iqSnQLehz3Ld04Wf0/XhmV2dorDr
Kjlk4BfK5NFHmKz8FYKEh8273FFs1kBQqFmnyaq0K+s2gFwFATCq5uUg7h+FEKy2
ETEXosiQR1n9MoyAo+r4oI7L+0+/li0SArtBfEHCnv/3eCSP+YPEl+l7pSdPUvji
phzX+GpkSeHaPBsvtBeq2jw343z+M2EVixJuowIjBuBz2OOmCJuwSEX6M6as+sqS
8QE+9tB5ShEKFpDpJ5t+dZy1qtccIL4O9Nw79ovkdtlRQdtnzUlf0LajYk3dkE10
by2AnwH46XpDhaCILgzJvP7nOZZtAY2PuVQE5rz4xVFH3C6/FkYXbTCDxfeqt1K8
H915olr/5wTfL1FXDlktd8LsgXJlKvZlqfcBUZmtxIy1tAV/ZI1Uw/vBMJ7znhwp
GFuWf+j/M/vBoHyhU1nJckbh3AOK6mEqDmttswpklxKYKiQIhQP1+lcyPPk4O6mk
Ye0oSEVKzpfMgEzU2QHKNxMWCww8ZnK+pXzoN6G7GY+0Dgw0i0C2e70/b0ykN+1y
obfv43SbwdpXV/Z3p5BTRW68tQlQGx/lxqH1cHwkkTNWru3By5bMxYGab3a7SqBc
svNkGwww1WID0UqhiwmW5mb8Yz11hr4zh2idCPiI7meyL6MBZmBaSG6I61yyheIx
BCw+yRNzeDXtQbwGHTImeGmpQH7et7RMtDwBfwBdRpAB1lwi99vopnO8tn/gpe6A
e4Cxc58yihcQP1/cigXZCALPxdRpIfbuzqmJi3Z3ljoxXbJ6qCJ9LFKm3z4m/T34
/eCogaoeTWZc169jJsAdGJswL4MFdWbzPY7raxQxGExdhhSdByDEhq02D7FK8Wg7
AJm/oJw9feYjjiNvopp2lZb1s8bkcwp/0t1KkmnhDJZqd5d1vEsDPXz+p6Ms6Jly
s9iOUGuwEIMhDuLH53G+t6xdE8qyDpZILD9f/6e0CeVn+ppNl4VkTBuMR2jm65g3
4Yy1Gz1yI5QC83NeghgvrwNi0IECjb7RZxkOzVRaKUgBDI+7r2YIKO46/bw8/EOy
T4L1+Ay4wwDnzM/QL6FE2zEorQTNQq22MBYvOo6Ku8VtyLrT68lfCBQOCGGVMjIZ
T81DvThrPVjJFWaGl1Z4ia5OHNwHlo0UAMVH3cswjBR3f0e0EQbMNbTztdOXRwJu
JehsQ7XfLmhwTohaHd0VMGMi+IqPTp/LuTUCqZMTcCj/r5NR/tRcV40lPurPLk1Y
tn6KPeyQRNOEG21OmMeA8pItWZVwtMopq1wvqmRvs2SJtRb9/faHD6yrbY6mwwLj
bAT9iwOheKRtHuyn0VIi8gGRAKYBqQGKIFP5hX8LG2bmFrnppRGZykaMij/+wNxf
TkY+UDUmbYzFfoYw5lB9reexerhTYGeiCqtQsD4XDJLlchPSMTYuJZYFWUMiqytg
zhIMN66HeGWpKFXeRVO5CozHrqlIbyWezurf4qpFSFg/C+96+UkInGele8v6AdVZ
2PVGmEbFh4IBnW0FarMYnvIWfCiZrh0nmrhPH+rwLel5I0TvVSp+OGFKrVFcxrjh
XqFiBatjKy0vpZsZhi80gZsaim6XsF3DEkIXVPxGVnYk295gfRM9v8s4MXDoU9Dy
l8fIod7dcC0gKPi6hTLQ8waOxt1ewbw481Krl35ZMUy64TyYw1ewgWrWDXas7TDB
Qc29AXmfDgybDAoNxeMbenIgP2s2yd/duAG4eOUjQWws6Ajy36ho03517NdFDHS1
lOPaI3jJAavgl6nk3sDEKGbvHhVRpGe/oP8fHAv+FiEeVGY2HZcTcTxjQCnQCKkn
4yTOIxsu8hkYFjzRyr4VbNDi+3XEtDcGP7yvRMvOCcVMMOEoJbQm5HVgUuj4rlf3
aCsP4izAeHQR5o8yCDmO5fgWk4c2hNaeX8nKQRMCvRISJxXWTAy1Ua06vWLjszmk
wZpqqWpAbI777sPv/6/tsjO1XHPds/GDr5L4kcm7w+IUZAxOFnnOyefDfHX2dYGo
cWlb+553UVc5ytB9m7InOKxoi9ZDdyAUtqupB5rdfYmxbJgqAAW5MLGpTILcJ8RX
k2FStMndBc4ViQzs20pQX2FO8dsCKWj6XV0PppePgnCTL9gwpjn82qL/TfDMxRsb
L1aMMarfQ06cmgrLOx//IG0Bi6Fe7nrncMOFV0SG/hJ9LBd+mpM16BYrf9QDXYZk
wQthhfTwJGUYDK7du2HtleWhNCt6DxO+pWdyZgvo2qwxdWJLao0vk9EqGN143/bA
YnjqnVhAcFGODcSdvVVnFCYP4GWzO3omMl3vMJanliAfBQ7zOAcKSCLTe2uuGFnK
knhStOXhCj8P15XBaQYVPZ+WusP6jAH/OhF9tnXAllxNJTZD5qKEVVJZgtEPXZZj
6HTpVLy+2rvvl2/LeM2KJmj2EoYpDarNQT10u98gNoTU3yb2DSnNZQBudxaJ8rqa
LLPVV/9O2OIWR84AueStyVoci57jOqMu+q0pKJUD9EpjTdMglAoYIvONr/fgG8q/
UkgWSc9OBvqqESMN1alY8rdtKUwJbaua0Oznw5cswaGdwld/GrAGgaZUZqZI5uoV
GK2c72sHIPLEeoc58YzZz7xLd9Lsmc8rToAn1m6pKfDCLyWzDqrnAM5u7uJVaqqZ
w6RmAcvRRkgi3orjvvStB17vV9hLnDylBAwmCSlMJNP/VDY8k0DRgb0HWxHKCrXD
eTv9So8EYanlhd3NTLtujemGYiWwRwZ0z/uDY0Ea7NZy6u9gWnCsgpAr9GZH/rgo
Axf+mbV95tlslhUEozZ1bi3bykC6xPDtDJFLVsYIfU2flEdY3g63YSwVnRfoQbHw
jghNf3V1gxf131p9YXJY4TPJ2Sc3mMku3ebpJjUWkU5iUS8mFvvJ5URYo079LtHY
/ZSF2prGIoTaGNvSKZ+WBp0+xktj01DPiD55lmAM6lPODwdPu157Jxyk6xBIuY1M
yt0L14znuBgaPQcd7bMyTaFhRDYwoBEv5fg/v+ScBtUz5JPK7LSjAM6UdOAgHbvx
EbZ3o66tANT+76hjJujjYlMr17bjpne3hjjTINQmHuMtyB6QNnDE+T9Gy84G/jIn
36Eq9WU5I3Jqj+4lOcZBvItqi1v87dVzHeB/u5KWoOz4CYvIE53xhjAYtj2QwbjV
9d52Y4vxB9HfC+EK0hyFNO/y+TCLB2FcgXMNXPFV5/BMbz99YSXwZ10m9MNL8nMp
+8mYatVkWctuMqo8TwmUehMDZZUpD2CX7G9altGsFcDanekfhNs+rH9ySzWUFY9Y
bkrxacTT4ukCslPjZ1vdIGKZCJWH5KiH5dk32xDB7R1ON5GuwnKWpVGvqvg7TkzI
meD9O3NcHSKTRAnQZuM+/w==
`pragma protect end_protected
