`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
V2mTsho8Y9fARR3b1VmIQ69RpfAwaReMH4yAVRaSsXUZJDYV1OnQYA7pwcG4Laz1
NMGZ5gJwXXccE45VqpexI6Fp0wUWhbU0r61UO13a16dFp29CZV9w17q32nQYx3Wj
+Ll7Bgbt+DJcchYbczrmnHmiN4lB3YjBU7zdrY/XkcY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10704)
YPIdj3XjP+nFzR9jSsbeaAQB/6TTA6yUWIWgSfOo9PTLzlNutfiOa+FGt0iPSP+/
/8N7dwTbRMxKDClAoSx+6eF6frugWRA9e9VBo9OIP42JwHxFnRQ5+OtrPYBDWCqy
Xirgdr0mSnH0DDGbGt8fAvdzjuGBJ7uDmYjMiNnRAOIGk6n9aUaFmByXt8SQjd+E
JYrqwPrksYRfMuw0mkaR0W0LxEO9Yt+FL+ZhRBN8BHj2ihMGE9Q4ZxEG7AoqQQ0Z
5P0IhPm2H3bnetb53KAxMH5fTgcLhGX/Pnn/B2XmH1G+CmOnxfkV9H+Db1l3TNOy
I2kWvpOsSxnUaUtjywosYEdAEUUtgDE2NDCdZAiLHWct3FP/r/LzNhEk9EZ2BWOt
ACfU8TAXUJ8rc8P1k2OPaGwZR3VcwJwwDugAB29Guj/iU3h5FLBkuGPrSda2zOx+
honKq6Ipu7EZs0Cyi2VwBcD/dOJXiWGkkhlRc9ZrEyc2KICR0zVKcX6WdgMbYbl5
krkCUJzbp/ktrKtGl4q/9imQRVlpbv5hm32wOoqR+vnRLZA/yIUbJmlBrdjTnz9N
8KPUX53WvMmbRO/mf3OqN6NImRmANH9v0jcbsGC2b/zUUQwh2yP60H61da5jfJbq
wRe9bnxbGK+i88x01CBXQ4qqHVveXShvlPO3RMqkf23TSAZi/rn5HSK9JvAyf5n/
OGHVxMFeDWbVa3xXwA7dHApLgRiNYHWPkEY14WH1wTFADsVTGY/1oqcsie+218hR
ChpbSAx9JNSgBG5D8i0u6JIkFZyr3RKLCLXsyqEoLdYwj3SDr8a/CWq429Al5dvy
cYscjGKVwvQiv4VDrCkYy9j9yBtejq07W/jKoAAKDbRFQoLgOReJQa8tJfugWsJt
XUv8fcIgZd8/uxhHnFDYVfuRtSI3EYI/1iXtVX9kUrD29w/v/yZ+WoMdNqJwXgHI
ZHUf1sxhL3EnulRwRvGFB6WAiiusTCp8bTAQXYnUOkSRXR7s7ivwi+plKDOcDtd5
dVr1Yl2+U3o+FQKS2HvpjhcCeS4ni8aJmsZGE3dte9Efgz4vjaa1gBh6NHhu52Wu
O2LyJ1pKJ7Ak3S0oj6pK/QLjguf+eOHFWOZv51PbLqmsROguZIR14SWxqBLOqO2V
52vBQPq0fo9BNXdWDKpt3iZkCY/Lgma9v9a70IF3Afb7JkIthvupgOPX2hIqBgmz
n16bGattPJO4kVJ9rj0d8/5/tg1D1xrE1QOsdQ2VLuAQp33gwI1XU4u+bNFvctKN
KEO2wxCBaXR7bYGIJQtA1Gttfry6fF9d3OQuU9w/HktNbV7zOFjJMmAmpKhx8kgR
uypHFIGK0jOUjG+iSjUPymzAo0KhK0HVtdKVQ305E47nGq4wl7amjzhrC7fsOlYf
5uhc2hEYN65PSkGJiXBWTjj5n1151ZitTkkR1OrWeOaS0ZQryTSlTNIoQ4+Vtycn
LANlDwbQ38G+y/mNoXU7o7WbnQxw1f6TbEkPr18nyzJ2WMq1cISKN+KqT51kijnj
e93LFsBRNiR7nEKSe9MQNZMpGidveedJE9zKuZW4KVfho2rUqeN05lo8W04hY+FH
w/yrre0LnCYqfTNEW6qlamyxJ6B3XHhfdjBM7AYiID46JvqY9BjpN3LZmidcQGvd
pOa0sB12Pc1yIJIEyUtMF7zHopeM4rqdJ1w6hbZ51BzmPOMFmLpxa9Ay5UYwrT2E
AcbrYm5sFFeziSi5K3FE1j0UW23b6u4xNDmIjqsyD9MkOiN80x3VrneGAHe+t1dd
miE+hhXEq57r5dtXTPyK0qHcfm2iOasc55mphuV4NgBFQWu1tjfG184GaNz0D8Sx
c7c+o9cAMEehYMtr2Wakjc94Gi3RNZrynBQNpHyJdK/ifCMUNJ7BDCKaKtr5XT/o
wQ+pb3qmNYRiTESzRfJ7A//Swg8d3XxUfhDBgDIp6lGm9y0jTTOvjMnGgyzuh+aF
2PqVdih8gXZHUSrJfpeu0kGDjjfHrEFu1G6L1b8cF0EWy/LwlwzkYC2j950b3D0u
syM1qpWMdBIgb39xWwrBSJIFY5Uj+2PzBKs30dzo8DySR4c5uCmIwoERZDYm7zGn
MYJTULndW+bV1jNWsekiNryb9lKW6LkJ61KhO134T9Zhi1sQqrtz7+7tlzC6jU9d
lIdFcr9VoLi7bZ/TZjqAKDeX3xrS6I9oumtUtQg2MXnJADlYfKLXMvhI6HUEYIOR
sCUGSJyuiqxOaVx7UzjuOX7w+0Ws9PRCqt4La6qEGvQ4iIjXdAcK6eALjcqosIOo
X5/C1zK5uF6cyUm1Qu9RgvvoLB5tGu9wWK5TJ/X10FOtLGEB0TbB56PVsMmrDBM1
hNQ+wWLsLkj5Ri8Bp/YDd3XYB1STN3YAq3NMgmqGVeuEZ4p1aRRzMDFfvx7IizmQ
e5RQykVH9Lxn+FcLTeo5J4+S8/z/zgyIo0fPerab1FQx6VW4stqsVzPHWoGNQpmi
rdR3relUQ/aC4tIPu4EhEzuFNJMyqLy12ms6NwD+C3xteOQmHw3PyxvSCOpWzZ9h
GWD+UoKTd37dx6kycrIKlFDYf5qr8XA5jsNSoa3uyrOzmSC5Yr74TZeyFBbv5Gy8
zEBHBe0vStUSJkCN3vCFUv3U7r8uMOZD+VDrAUd9+gSEXesjcDnfXsoTOmv9jufU
8ClhEGkVffwnARsaNvXjV1W5uGdGRaaFgEh9/LV9Ga8fBK6PMLNJ2zuShJggBnPK
xzITkdt0z4YyR5b5B7F+4o2xOiqsQbOyIYQcz4VoTeEc8iOeJLVKDU3RYMCGEFwq
3wbEoCJoYIdbNCOd74sfQmY+aixeJyIk3khX1FoyX6mgVi2uzayxetk7dguS4F/E
LZgKeIPO2HDC9HzQve86jjiwzyBJfAUVDYVdoUGCCpidgPOKjw1947jOgh1WL+v9
S8j9wxF5zWpNAL7w6Lyw9vXFUhGDOc0jsi3NUuvFBD68NfLdhsVDYNg3ty9mzrMy
bBmQnPE/v7FW9dtQWE63nTiqa1O+JODuAOrHa5usde2Vxc4nObL1QKjhIaw+l2RS
sUFdryQ2cdN0iSO6lHgPN5cVe/tzNq9I15fO6Ms2eTKpQD287nZ19HL/I51nN5M4
raL8nj1vmXzxVldAVGb0f48D5c441jEnLqIvody3I7qqVBtwabkaB/MpijY9h3I2
+i5jZWsEABdPZnuZPHb2y+8arUzj0uPnG37GJD9qJu9Jlo03dFyWZAtUeTwVmsGq
IdELh6ZqEi+eKyoBCe6gJvYnCVRdXPkI71pkpMKY0vhOQDWzjmy3xPMSAZSGarzQ
vsQmsDUovNOFjO8PolQdrZGXltkAmkUhMOJ48sM4QvxAJT0AIwOoDScGwYTmmCXD
U5yuli+pPLg+wmF8dfsienxCu5qeYYkEi+KoPIJbxXKmOBY1P+rS+SMvO6BiTOgn
Sww6GExzR65ibX6aWgmQA80/auHCbD37hbICp9EWVVHVmK+YAxbuSyhNOhxjjSAx
HYmEnxyn2UxpixS4GUtPDW0Ch1WJw7O0kznJK6hmUKc6LkwQPAncUvZvKkkzR/Zh
8vnw2+9OLwngB3BPZtTYxBBP+c9g7PzDnCchECgnC4+kUhRP6/YRfUGUGD2mzBi8
o+TA9Vq/hzkHpcfyD7gAy4YNyXqrYqaBiHL+e0jJXXOKeLYZRA8XdHADKdHzGpxt
88nnBbqjOYL9Y4CEvaJzHsQtOSoDhIEkL0fYpHtgFVF/R/NXPXDi0FJpFSBjaSu7
Uka/8I4v/a1MNkNZOHu61XQxQH9XZOt5mSR7BTsmjpo8TkNHaA3O0IShfSUt6R/U
bv0jRKlAj78wJD+qOkxL0pLPZP4xYRnSuwbQuddJRHLNB++Uxc9AzjTRthjltEQK
kMQpUUfL1jKEv6IrgTLfCzsQ6/lXRGSapnYSsa8qRO3O0UKjXiJ3f8fDYHYs+Mog
J74/1MsENYvCAi8TfMCwh3U6xG4fn/rmdenK6utC8J+wLNHBAj+oxGO11y2Zl4q4
7KU3bu5+ckhBRGJtvpyY4jOzxPrxXnAFwAIaXOmgase/gq+5LgquLb8lycX+3LZw
OjmovKphOrVBZfP94TGSIDYwYXMRuQaY/GsUh0UB5PFuImyfgYi2tbv0p7DLW7aN
cG1Cm2xzznHYWYJvJOqd0gdbNgpu+jnrlDE4ZU4QyU3BIqkiJdJD4TTyv+FLMv/I
HNOWKddC8vGIsCVoZQKpU1QUX1rEqiY0zBtSekpNSFJ/obyfMDBjEMrbzxjOeA0P
szvbdl+EUaVGN/sZBKzSyBpoS+9bWxa5k5vZpz6d3Ec76WQI39dRoRqrGkY9TQQw
sLFSMCYbbIQep0f6GuxAHvn5wZ5UInXnc8aeytFsMv/krXXN/33AssXP1l90wB16
PGIXhjtvVth3Bc/c9WwuBNnSF5ui/hh37W7CIhZiILcYkUEvRYbqJfqRssnBrSh/
EQl2igjBZUcHtzkTHN1jAMvdGNweplkOyJeC7KdcmUhY5Y5OSWAoaubCxOjXJXbY
RJ0/mahqVThUx/19rvJxCVSnIBoRwP5z/WdpQsn7xmxKzAzeic+3vM6dcGGnlkL2
DHpRv2HpMqvdx+tyH/nOvmxXsDzH8n+S5uSxTFCKCjLAOVDNN5ZQx8RuiVf86VeD
AvNDjTbRJmcmy9dLbwdsRVdIWHPaewGwUwiC+JoCNsYwWb6I6c0lLc1q0F6iY51W
toGF1MeaRqnkgOOu41MmguecSLFfGOW9PtWDmyOPzFy2bjdVZjnG4hvLKVJp7SM4
iwe2EzIgs+OsdApnvoBjTYQHb7Yu+TNLAWxfdBHVMuUMT59A4Wja7T/Eb//00G8A
B0cQl5mwdajhHa8DLvJAifwYuKsIf17opmVT2VHCpOuKL4cNIqArBEiFNZXFZufz
fKzlaLSYtP9pO7fuVhNDFMtbjP0GPYQ7tsq79cHjDoZpJYvFboZXMvc0of/2h6Xe
e8m4vrINdWvLOYVYr0ShUhvDXZWrsXlPg0mxacY5M/BStgw9XUBAQPjdyEqKh7ky
U8cATy1bCCTPbmoST3JrUBdlpC1pCt+VZcWHJzidUPiltYRzI9/dy3ps+LrsxXL2
m83su5yxZm9NNoIeiTp6uy8GkOytDIOPyowfD4I2QikBw4YH/qj/YhdOvduWbtFH
00LdRdcXEflxGTplSoQyAWoXGm1mRWZ1XdwP8bbnNKVwHLTXlmgVorVowIYq8ApR
/mtCkvqp2rLUn8lkvXyNctlJ4OqQw5qbp6nFDdMFYvtrSBZASO2oNQ5HTpIt5Z4w
rqdD0CyHtaV1KK2hgxzrLN3ppQ2tMFAC9fwSy93r5QPdVZDokX3jnqdNnHkz99Zy
Al84QSeDSIDMQxGjyftuhHxJ/dEp4Qoi6XqVJVcTNwx2K2FayLP6L5tYlHbZfkfK
LGl1OzkrqqvL8G8uRTB+58jZH+wsNZdK+PfpmupbsY8MyhSodVo3J0D9wk4Jteir
Ye/MrxC7xjCavL/vwO+orSKz6Y71khW9XgDoeVeeFbJMLiNcucJl8KmFECIglPlH
w5ZmCESNI0X7ePqxG48LkXhhgbgD6gCHBB43rKtdUS5YLKHn4YXTD45sThBr9uNw
+i3mmYRmLX2sLLsqnb7i+wfQ3aTVfnhvp9LP0yG4GbSY8fSbfs13fXSO2Aqn7fFJ
TE5PPrh3JOU6AeiYABepE1O+IIT9ZphGY1QpnS6b3cCzCw7J4YKdykp7IJuwmQrV
d3mGa6ILp9pP+w5hrW12lsL7WaeuCFyR5zK5EqKfZzixZgIGNDDHc7SrmdI4rorb
UfXk/h4MRsSC+szIAn68GKI6OdrtMsrduq5rDAtIsdllKfSduug0rIsjopKECfvs
Gnmm9qYOJ3hiK/oJztcpKELbvGIZDjL9/ZeAdwKR5sYD00c9jVeOgoRRjSDliZAR
QzEwO6MNqS4u+S4exGCoxApzPSsJOlgNssoRqU5hnu+VWEh+SdFvcQWlCJHPh7gp
wIiz5n4SNrOndjJUiXOJoUm/2xxfvVi/l56rvSh0mw/RFGzzkLYdaNx9VA7BjqrA
sFFjXLGfkPPTVpnTbF5YY+999inT1GMA2I+//H8dVNyy2d0kwR/Vo14LRkwuAgK3
FVROFrxq2j+WrihqwIIN/+d/qklOcJnvQNNQ/gUQ18LgrsHzYiz6E1f73LmSIdI5
YYACJ4Ieg3Y2gc9aQQmhDyULfE+unp8hlwBrBnAZofVDwDGgxqZEz0WALBemc1BW
Te1Sdy67qntRRoLeYmf5ZMHYUWu67V/JXtxH8o9vonKdDtEQZlAXAckQ8xDxEcdt
Otpm835fzcYeCNRH/ciunWWujQvb2vDRYs5+57MXgnj4405Gy4BdL0o2cyGGdA8k
hohR58prvmzCJq1wzrRpBI/isVkgVVbhPVmUOKT/YpXU3eVPYMuwx0PMP2Bz6wel
Qa8KDtCYOWknBzPUXljjH/equX7eMq3LuKsSdVo0Ml63MNYg2z5+3Wym5Shti3dY
iZqX/jyvZtnXql0ChEUnsLgxaDul+37RbTynePItcgZbDIZnu49ONWmJFd5i1wZu
DH1B9id01svWL4nGVbjx8qlkhXv+NPk7sPlkyZ/Wlia1jHiFDnP1I2JPHiJ8yEfG
nwDU+kirZKe8a8G5rbx+JT7ef89tuYqSUN9wO+IU4su6ddndra+z4cZrPi4MoEia
tTt2XmZ/6hxFKz3wNV77LxJtQVvbyPBScwaxzO1764Kh4+ICi5foC2NvuxujeTc/
35esOY7RfWJad743/QH+ewYupDQ7yEL6RA8kgbJmeALArlMlLFsmXQf2iB8rYuuH
147qcB2+M2pKDrKpQJOMv2ZCEKK84ke63Ka7ts887se0DuJl4pyivd20q9JuqKHC
vos1P6il9UeY2ZNUVAvPWdoL7iSBSO95yNWfo5V3Fat/kVXh0fy9Fphdb8IhiKBr
lwClAAAZslRVpZcQ1En5wLSaKV7bc4iEyzKH4iJ9yHf3I1rTCihPCmUCbVk0rtE2
nA34DIb/YbMFMwfUr/ZQ+hgzBvZGHIvWwuP65dqjPGEXUtJ092jlgduYkHUJocz/
FhYdjMx8k+RpUBOkk0uLrHW3Jsmc7UI51WiDlK2FYKF+c5CuKRO0REAVf3MZKmRR
IH2WSjWG76vvT9OXUeKgEk2G/Ll+NOtMDkpbTGUKVNifu/1erMzSpDDHsKvWTTOT
AhRQkP/oejOTRQG0RMyPkUeQDPAKs3Y+dLVCHGwt8YvxuX30J73YQKFPoMKvyTd3
Zw/Au0Xz4LJJO1jTdMEw7uR+9dOt3uayyutG/l+ybnZCej+9U6Dpzo8akMyjlTgL
Zae21puDIGwo31JW2SbZVyIrJDBMdB6yW+4xljnNKepv5Vyv/MLL/mJxc3KM+Lwu
YU2WU5AOGYfzCeT1uvkcbDpHQoykR6UXb/1D3QZ/FpxQMQJdVssvSQVg12Dgben0
LoE9DL6/SvQp6fDLwCs/aQreu6nYxFoJekGzWY4OP7qv+zleEAebJWGimRUS6Tk4
w+QtD/xjzkVyNIyQzAPgxHExfsKxty8ZjNLW7oG23rkyiaVoRUNUM+APwE5KE2r7
W8888pz2EQNQNAsm8Q2OyZWMrfaJVV7O31NkbzHFzaPiD0qXMbsYCjdWewXNFt1n
46CkjhYZITGGUJLbqWiDrz38xrKDedD/Fd3Cn/1KbKajfUR81TEMN9ldvKsE2mzS
rVN2Ls0lnJ2rOgeyM0yjVOBeyTegmvpIjOOfHa6KsZ7TeU1u+dqTZWM0EOzlIxl+
teP1MlPQmR+bmhADBTcy/apSvef7nvtWo8KnNsxtnOwOyrfBDOBxe1pZeMaw0NQq
nlvwn2wC657gVxYcgGtdgAQPf0iPE7EBdMdQoheRBWPyNeKdu1ZyDzSfaCkcu30p
t3qBUdRxZ6ZJNNlBEExPeAuaTQ2VYckcSGz/0K9qlIH2xHsj6h+fJzIyIwlaEjlv
Mb3Kdm9q1oOfBLsC9mHOlMxo9s/gbpwj/kUgOLJpuI0bAdOqCSDPHyqMgrCdtdK6
ZIZvf56WRdjadUNPfjlKAQBxym/w777ALBe5GHdFV0QD2eAZLRqv/5982f0P+rWZ
GI9dMJBiwEak4eoMmvgDT4q8UkNHEsz1vKhq/AfS2JQ83tMzFCx8GVb0g0rku14E
50z0B785wS9Cs1QHup/vzYuu/Zs8IS087zLEkoxq9i3AM84OfvdqAteVWYP3v2oS
Oe+0cMKd5y0/VGfZRWZvSAOZRljuzAyHzcEVtp/LOGBDzMJD1QzZ523fHjnpErNX
/k3H4S4vb4SZxwYnzYHn3QAeXVYPgFTvgfWJwBtZ32pRwGz/6rnumiRB+/syik7q
cUB46ll4EquDGooH9WBvy01gyBiiImXkFABtNXlZSkBvvMX7xwTL9R8P1n0cGkw4
yBMgjnySUQwdeO69w4+xp0oCWfrJRMM5+RAzRbC3VpyTYGDL6SGQI1pMIpCwvp3J
0KJPLOhekxGt4loAdo04exukVWKDCxF/Bs5hNFdIvxTWEsiwealazekFPubfkGGs
ZyfPrZtL3oWFFqNKbEMopx+rOpsHD63FsMNe8AC4E6cMpCj+xweX2GvSh/3Qe7s9
dNrqfnD/jzSTcIPxZCcebvD9FikgOdOk9bgw/0rYkrCCPNLO2+btLLa4UZWkmKRa
4XnTUX7suR9GeCxwWLcfA5O/811sebx/nMbb67NwaSIUU8rnZZ6OtRtND4cbkxeY
KwASiKDOa2KCYxECXlSIKRy2K/2IZm5HZ26pgB3m6FCkncApXA/I4Qn6KU+RmiFk
PwlPIfqpQQ9zTs7vTMdIT8hMADImHuO7cY1eyPjNg7ffovApryiVBaZCp7NERUvG
c/OAlLHivQ347lHREkhHF0V/LP96m3S+nc9hx/3c+igZ/Khguj/XhzP+hAocVUO9
AXB7OfR0IQechEJwLuPptwUZBJd0BroPPoth8qmayAh+AZVZA3tYbSR8jyfVYhct
I71bYq7JSfvjvKl6N7pw9VBL97ISZKlduP030cSPazALy7CJLhVsA+yK7Zt12JLv
FtshIWgA+nVIVTKlgSubGFfvKjMOnkXp+OlbpdLMpmlSCmtruX0B7++R/vuBKTS1
l2zF59leJAPWfncacSoPe95TUvfyByDTapwOpPnJFf15EgPK+B/6M1ysMeqt+6HS
Fl8kWXbx7QFLGab+lQjik8qvmZHDb13vExNcLKCGB2mY4stIa/Oq4lVOsP0h+W/L
k69E5MnWmteDCuFDVfkQYjItJDETicCxt10jc1ChpsWXi84GsB6WKyxJUovLATCI
Da9Xg6FYgcIA8zULGPP6GiN3jyY/IFnfiNLaVgKM3rFgcLFZFKn5I+rttfpQT2M7
B49GDJCH3/P8Y+3mfmvxQ8IKAyecnzxIlAMIvIAfl99Tjak9N9RlfWfAQYXrUQXV
19GmILF/saNEYqTSJb/ZbbshCzfUvZ3Jhl7ERRdA9cGrXAylSzwKBP0o6tWdE1+j
qYVoSJ8VBeNQeB/+DtFOnEPeC+LB7oK8VGOHqucfzumb75TUtDcvPsVWwjY6iwQH
yV8GZ5aLExrmI478l1+bOwYxAPxL80D5TvmJXzaII5VMrjJZM7qJrzRTHGrhBnjc
c87Q0NwmL92z9p+2hQ/NSDXfbrQ1Nnw356nNFxhfn4poSXaiNwSQyCKK/z2AVjQO
Buy48GXTnhOIYkgj9l6FqbIZceW0al0bac4JO3kQRwuRpIcDUGFn9xwYkj8V2KOJ
z0ZpkapGbnhFDTVzYvXpcQNKXWUdPJifPX9Ni76W5CBR7OBJmQjfUUX+16H2YmNi
n+FWAyq1F1dEKSnpA1+GkKI6n11FGKaAYjQGHeqAc26q9eQ3BLuTx8//RXZKUgra
QcG+TthVsSxHgMWzTm4ZZxvlPWxw1eeJHy4pjm595rRYqpLeahkGDlWUEB4dNWX0
Up/AWflgx7jPEME47Fj9RJxrA1m5jIeju7VdcRXx1ZQTilhOA8R85SBnQeMdIBlS
tcnxItno3HT5oAwU1CkjMHxkw2KrdSJ8EiNXdImQ74WnYKP/wlTgFIyUGMrLWCjV
eY91C08j2Ux+G3Ylau+77sQak7ZCANjgApeu3uJIIZlJwRzRd+7TQYpqN/t2dN4L
Mx0Nq0Jnpg9mq/+Eqy770wb7kBsIFY9u+r2dfyfvySCpN2f9GRqIvar5wj4zQVy8
++TrB0e9LvbSiUj1ATaL+XzxXe6BCwCdLnH9VNi6M6iG5IG6/rsW3v7Za4eLAk37
gL6RadOJqnqueFSdZkGA7ETnPnyyqteJH5pBOkSit6kcx8h5fg1RJMwFo1JxRAQM
706NaO6kkexrbovKtGBNSWvFiIDnBfNBo7uu/ErSno10T/O8IVs+wKsbCAta3fvz
XHCfR/d7FPpTipcVM+Gk6+2k+8SaZY0ytnIpquUSif8RKd5COdw64RAoP6iuUKZL
jUL4cmBRtqpfRZxmpCRkUZ7VIqDd2xCzUoRdEpTWI/eBStY6tdtcs8BuIeUGLu7t
gaFaH9ckiHDvXZQsM/YLHBloh3uQpDvQx57CbGh5V6G2LjNQKuauTbiBW+MoLa9K
QSDwaZLq2/itYjPmHwADrqOhLA4RqyWRG1EiZkmdlSfdXHJ8YNLfUDsKAxNDsb/B
Z11MW4Cx2hohoS0XZHLFvTFWnvOCwiijkXE/R8MPQ1T0QSQKMceBTie8eiI0s3EL
FtzRsoV0ylb+NsZFybFRmjX3N0l7zKE6R7SyIPTbK8b27sHfwHxLG70gzGqspHF6
TJy0vpSWieoAikUypIbGTKre+emcxO7uO6qqrP3x4JwQTP5ib5YMarpfe7cn4Yra
WzQXFFPKM3wCmDGuiLhMQi+H64n8/wLqY4cvb5zstZpxP2X02ndN6P5Md0ZriKKk
nhu27YsyNSq4P35nwc5J6b8kzmHTEVdOiLKudmPGLs06E130N0RZGq4yPawDbPFB
kl87ESCJDF+5jWYVs0OQENKypxC5rxPwTrBMtqk+xqmGpcxAblqZZQLBtF/hTcYS
Xns67/PdCnRJEuEqPAjLWYa4vwgAUssHlKx7LNDlVa4vp1iZypC7KcQJxwbGMWCB
5RgfPtpMVm56lh7PMyn8FagpVos5cm7SO+hvdYptn4QmuLc5WygWbluWDIURy9tN
lZRF2cUv06ALHwKs4W7AIv29Z4Qd6kSwwlBMiXtw7MRlZc7bFOecTx0hNOCxWKMA
fow4EIvpQx/SkwDTfT4rqWyuyZEFxPKGhh55r6bnIQWCG4+uSrSx5NIyMvxLOFtr
xvOizROJUo6UkPLjvmOKt+fpCPF0TbSj4rK1T2lKtNzDX13rZSGMP7ug51JTZwYu
notNHKoWd0ONSeVkc4HAjbMDz+sw794Rl1lxhf72uQIpJ+/UivgS4CBANMo2vYD+
9L/UIgBtCIbgItPrvMZrTr6IhB4csLh9qCqQCcysRpWgj03x6gt5rBh51LTPhtUR
kZ53qXDRuv2tEGzTq8XbvcZdzkO/3KbzgfkgztcOq0W0/a6fO2HwNJ9O7eZ5BjDn
Na+ry2Sp9YLJ3ttrnKrnElILDqum3r1Q2xDLHl6vXdCT3+/hrPF0lNGPomC9vPKO
5EePuu5BVRSNpiJGL3HoP2eocqUln6LisFZFpmnnQGcxBM1ZqFnevaz4F6QlSfNc
EpunqLjLZJDMYdzCpcWJ9nGkyCuDiDXZfb/CgVwOqca2l22xEvhzTRyYp6qCzQna
Lp1HDvm9KofF+AJ+pYBlmo7CgG8DwYYZTYLBLGNYHV9ingUSuFO0+cTlrrNzEZgO
Y+UH/8XQx0+1s7bZjedZawJ2j/3bbomSPaGKNQJGgmbpFX/jRzcLRw4qUFzIj5hC
NPrVmzrFb45Iu+W0Db8O3CZTPZw5jXCAy+ZNmHxC6OxBiAsuP58N1UT23/PHRlF8
IMDMhIXTgSPBiLoOJ4WwskgABrrkepXYYE/4FV+Lvhu/EMZ+/cNvrpBfLPJjKnhx
zqW1V5kl1cMYlVclocFPPKHxos0GxxO74g+g5R7Dcl2hk2aYvXlAV+9pVJ9cNKp4
1vgoRqPc+f26ErjirD/1M6zgx88X6fI9D2g3F5veMH6S5tXETwEnZueJkq2pzkQy
5pzTmkTSWjiXzI5K7S55OlEv32YCHcBQKTNJarIMtCCGJ5P201HnIARU2Wz9LeGK
O3EtEqfrEWnfMkknkACSHR5cdhiyAh7BODZr+wMMmCqs+Dr97o2fh0owiR2yjgHB
8g/RY2X7BtT0R85qP5LKYSKMlSC+pmCUdodwU9PCl/r59pDExF0bSpATl2ENPlfQ
2nmVyqiVDVk0gxBUQfZWN8gCXY0M4+O/+iPl1RimAJqdZbFNzQwn8VKQHk19HAJH
UKpzkL48AeYwHAzF87SD34YSX0xdhgOJsP5p1yLiY47f/n4QOqnl6gfIeFd8pSL7
jbnrWBkn++Udo0Q1ExfIhtu09y7KX9xS+xJH8HaTs1eDYU4xa7oNa+JXoGSl5Ijo
xBs0VLQi6AxjQ7dw2xa/2Ydq6pkRSY6wHb5HmPTKcnX7mQnzaKooTE60uICMEbcr
+yf6EfAHUG6cbXqiX71Iwal9hs/Khz4KNFdswJuN90yD94J31Km+GG8rCC3OrSXd
FYtQnaq7gS8NicVWUPjb66So31ZHs4blbcad278Whr1W3JJB2oHUfU4hkQXvmFVF
9iGAnXjJlzJIr/xx1yq83FLa7WnJrP2Qk1Wn8CO6rF6y/Eb1gvqm2wefItmo1yFJ
xhmzsaQcLJH/T+ic6I+D/7iqiQI95CINFox+FYi+kMV6VpVCU1qw4Vxhbo5dxr0X
rvG6x5lzQoqClDTmRQ3iR4uvLduy4zNmMfTg304C2pRd0Bwz2vhIRwdZXeLhMC0M
udmuIx9Cs00H4VXxJBIFxWb1TbqK01Up4V8zbYgGgy3pzuK6pTHu4wdHzQf43rl3
Lf21J9t/USjyD59EVt6K1eHMfcR2IstGv1JILJU6MblDgCYrNyCuYNlf4i+agC9a
yuHPtZe0/19y79ZDwrsZOuUw1KJKpX/BGDhYEBtU2trIf/yOlDi0l92hg+XliYZO
KUKow/fXnGL4oIWfiU8DWg29Y9qzSlhUZa/ln6RxHKAPe6t7lP3ay6wG04z7zUZb
ShRWZAiJ6h4xhZY3mUI2llfHvxYONruOYlEFQ+sn7KzAXwyUnO/naXX25rBDszF8
UHzflkg/02YDuHpjr8zwBk9sxaVYbjT/Tl7qstqn23KSasqap/wYMOPyRCRIh2VA
rPGgMW8F5mQdjxri9PW4X7QfD0THRi9uZDZWdOU0DkTrJbzbvnEDeW4PoTCKh0EI
X/heQOH9lbKLyGVkchqUYFGQ+WdTCaeqT6h5gYF9U4lzHPrRrVwO3VHeTs5z0MH3
gOi+KgI5zKYdt6hkjmlHSTTNBfcMJjsIM5UoNBhEAkE2vos3i70OuT70LHFAddgg
lOYfBlbWQwAdVel6E+tYwPcdgGobzFmG4sxwAoydFe0qyBwlJLe8814qwMM/zlty
eAovFd1c0PfImWiART7STQfaoVNzqC/dvNXIhsZWfh80hpBzg0a/3P+Ekf5gVQgD
Iz9uKO0CunayGDetH+sFsCqu1uxorGri3RiqdrQVXoqmt2a2J+S7je9K2B0hV97n
LrYm7YhXdFBs313+Xb5y54TfAcZq2ucBnpEN9ldwk+7o+b3RUK538RQJiDCIbUq4
4KA4pN9S4ymVszeZDjd+ziel4EQjIftdw5xm/pOdMA962Qvm3Ia1DR2o62DJv7TO
8N+pgbu4peAE1UOFAydc2HIi2thdjYBdRgE2g12Z6wow7GvdCT5c5cjsw0RqV4yF
g1NCoL2/+d3X7V3tFTNwocQ53ybKAPhj4Q9QN8zyAZKNn82rlwtQBl2wFxalgin7
cFtuQR4oOsA5a5Mx5gyvLqPislU75EwJt9Ij00QZNpxvedkkIz/OlS61UfByvDAh
SHk6A29ZJX0v8bpshdxhkzY62YR3ErrsUZCpFpFLXKVkuW+wSN9FZof8PktuTx0+
HQsiZew++wpH5aY2jko0S6E/XZfByV78N2PfLAFoJuhZMK4Mo23GOyEQEbCp+tjz
N+fGGlW20NDB+TQ4jXVjqkR+9ZxNcvBd1aiGjUK0YYZ117LTEuuM9RXKrA0If9gN
pI2twdA6Ubb+uNIGh3aP8eMbq4KPdBkhYVMWxob+3ccpdRLlxDGUQDO276vpTRDP
`pragma protect end_protected
