`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oT+hbv1njRKCepzsKJhtQCh28P8fR7+ysE9h6IwoUgOkjbzbTjcutOCk/ffngUlP
naY/0k7LIyH+0p6Z5bi0nfaF/8rNXyrtTCSr097ckklo2hxAeyK9ybWIsVr7T91k
OWjVL3gAtWk6v6baSr0oflYzBhR1tjW6Rv62GxhQIMc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3184)
Cw2qU2fpVNy/mwB9hiVcckPlZMU8YaPqQ1NAks2Fdp7qTvSsSzZ2eybRS2WUzhvv
mXBK+AVAlOiStv+I2bZ2m48h/IxmsrvcBVh4KnqngguZdjRmmKmZqZb5VmJW8gKK
dozyjvHsDBMG3Ttbj2mj3no2FAtkAqGxT0NoMGaXgJ+C3yFn6vAN8h8kCDhRCszF
fEHQdo2TN7tExaTgljFANDMTWGLOa/sS5w/m++nVOynQaii1GY4TroIxgMWl7V8F
oFX8OTUcATgwG8i/62QO3laizY32P5FadXvBZF6dB+itlyJRDGCv2wMp/3cS6iFS
rI2FIgL+k4jC+NfvOT/gTyLuW9UWkBCpqRywy0fsNtR2AXgwfvy9vVfbiZig5cVc
kEXV8RXDdBm/txy2wA17HUCATdUAA1uKBDGfFSCfeBsWOIOjHaB8bul7aVDB0J7x
RsGZRVz3icrMh87HZF8KodfC0hF12fdtryxUFh2EBQYQUV4V6s2DJsiKdP5oAw27
mXtAGgzuF6MqxGp8Ie6Ibo06nlYItbYFJztN1vK7lYcIZrSVQT8JLF9y8ahYX1yY
9Mdsmq/S0X34XnO7+IfJ7MWCBqCsg+cI/qDXhonbBnrGxbLFa3UBZNVph/CJc3K/
gRTFdncBmGF+7kmb1Pc+Y+mbk/gNWzHacf4miX9mFynCBJeEVJWSd/RJa3iP1IVA
JaBtRMeaKR7UWHH1t1OJyTdD+PS1pdrtD2ZVB+V13/7Qj6Txqv0o/XPMMh4Qikkf
G4Q+t0YWJgr8tEOjzT8j2n5UhouIEGRXsNcE4Tftm5xoVoplO8OIteYF/S8OpBTr
yYCU7/M2/kkhqEBOKpdUIz15+e7zMv3vZciv1maSvqMleqjREImh7+u/YnbnW5Z1
/2UoZnqI3NwVYdXYkfFSf86bxalC3uIUAD/BuhVSxOYuMdcJEe6t4RYVWsg0wGQc
W1egIVgJqQD1LiMd15VvAb90sZ7eVXReRgdanlle8EqEInRIeYix+TQHpg7+2Tn4
VcTOCHGuq+hncKuUq6j6F/Uj6BzATRtphF8aQeE5oopfrS6MVHxwLqveh/PQF7Ih
mindUC6KVtSyJCv/9ny1q+AlURKcIQZRWk1KzkFNHE+vuSbRgX+GSp1gMCHGtKrk
PXAfmIstthaaFFIUtL+f3g8Fyt2KxMiiUz+MhBqoracCmrIRMCxOgRNSksPCDySL
LHqWIuZW3FOLL1d26bWVFh1m62bK5BY+K3aDKetT5Zt2Oqyt7kIA/V+TobeqMdxq
12NRBaC+tcVAjfAVoYmBrmuuq4mW4M0xzg5hOa+0Zrxeku+VuYA87cyiw+oOGgLJ
zNrDrzCGMpRTsMxZXEm+9PEZSH/vseAPstlNEPtvvYOhYnGAqq4YUBcZbMFmbsOZ
abEN8oEUZ08L9PWRSYFl9bAsPAxOM8nq3S9V5Nm9zi4B/uZkDr/vFZFxAGzjr2Vs
QnBwiMYqt3E3EnDcvM/CR9pGMe2Ov6SKYxlzeS/bW3wnlkOJrEwTk8cYAG4b8boI
V81WnSKznrUPlHSXigFJvdUM47NnzfjC/v4VXGkXrXeosdM18q7vkUoet48Om9gM
9V4aSE9PR7CiAqaOdaBBmmfqESgFAHcK+Pvdzei4zdwxMGnjA4ml1mWS4WO/fTzd
8InQslC6908vaWOQ+W0AC6dgpvq5JxM4+prtDSvtVxABAhBkLwE4Ec7oelhBT4N9
vr3qUXmeW0vDWZCJZpklWV0rHjVeGS8XFZCRtOmpgVlh9m9gIGZ1CSZHHlDF0QzZ
fHTbwyIBfhc3cMveneFxXABlbMa/w1/f4OnCpqVfyqPTp45pDCPW8vYJxj4ghDAa
qkiqiBeFUgHhv7imXsN0uN0T+FY7OrW2ECHZW6Ng1QtQqr4d7YXKyJyknDhsxEVV
H32kahT8L5tFM400jccMY9MomBNvekh9tnMoZPIk1pXagu7W03bvoBnnt8qU692c
VSDswLpA2NP+d8xVolhgX9anZbQun4+1qLa3DbWELQYvccwWwnYItVzI86ruWJUk
egu9NTnEi/C4F81jvwrpyzKLtc/yAiCEMOn6YqMIwxy28dt44Vr5jRpj9RlFN4as
piQ6HJrx4XgMLTGGnwkf1WiNsC00YSCADqb+YLOHsVxPPqQPxwdsg0JVYcwIXZfY
zSmM3d9LYyiedEjO3MGX9LRqCNAw/QVvTd1UN9NAuEGkv0s8RBH8T/H6wAmSThDN
ehVvONfXsyy+6tTgg6qEO4aA8W8qq1+Qn44qRsLp1W7Roh9YGAjkmtHOOZno6GPd
E8tnZypsursnvz/bPjql+HxkMCW/w+Fvj5C5RbGhvafNmcLTMArqvIdyN5NEQDbH
mD9EoY40JcS6FnYLrid9OPpp2KkpNnyrhcqOOQpGk08uH6jlqcv337T41gO0kQVM
PSiWZb+tovA+kgb5Hz9AwJawo+wuayxsb1w7WjdA12pMqLcx9OdXXjW7tTli9zub
jDGLpb9+5s41eelNLLqC6OZXSok74gpl1M0KXV/LmWscv4TKDhbfHwfpLkYnwozq
iVdT7avGWYpJWakMMapMrsSuQqmJae/NSuNJfHagoM2ON3D/kHNefw4KrOVfZWN+
oZ83YvyHG4zC+bkm1pUEFHIE+QFYWfLzxqEwFOCmdMkd3CvBYPRFaFQhQAqGukkp
ZUWlTgUwJaKEiV+QSgjJNN4MGahX0rvP03eDqEgMnmeaETjywusADADbYyXkRe5B
3R5U9pj5FSMuAIUkSSFw/ia7HSUJqwI95+X0XWwM4QMaYP7yIzDR9Xg42P8pF+vf
WW3md1APEY35XinyuDBvB5JOo8ufPlFdrcWSZxUDk5SD8qwCrdQL/DpeRhrEvIEK
+sAqr9uV6ayGn99nEKDw5s5n8JeX72Yx/oxLqtNyOj8OwtwYt3euLMVdj++TkAFu
03JNUaf0IAELLwC6+FIjansQbe0mjhuGMGMfKcWwY6CEp4/lREyqtHfln9J/b4HR
EJtRnat0H2L6ukyao+fktllWC/E4DbrAPHGm6qUiCPljBUu+6c6JZjhIaokubDSk
t8EdT+EHfn2uRWYTWPXoWc7NixOkcDKC8HJtNqxG40DsiyO+SAAJ/T6qOEt5DadV
ipsewnqyWD/wICjfK2ekoxUaCB5LhTmi8H9TTCCo0r5G8cbxUiPtZo+CoZoKBO1W
TFM4vDjoEfymX7EN5LZJnD3Mea6qJkn4+s3glmmT59QsRZKHNPrMBCK5pWOLCCHb
c7Z3kLWj6Fy7KbS6CwrjRQfqG+To+FlkCUyL534+4kqFBBzMK2rUWOBlZBBfb5ub
U21Im8gx1Mwp9osDQr7862adc5Omtrrnx5q5atKXgMZFTwXA/0jYQ2WZ3yMlMXdv
iz5e88PeqBGR9YcTs/oiSXvWF+pQNEcD1bH92kRovgVj73oZJ/8OzqO+jQXQGV4H
A0EKczAqutseqbBEe/VZkTSGzBi83zlROQS5OASMMSMRTHXuyEEQ0PnnWi27+KaI
PRONBDoX1QP9JB3t2YNPQa9t9JL8p53z2mJHbc37R45nm7qOFo0/1XpwPeQtQ24z
oSrDuCvuzMCcyWVxPfFsJtUmlFrckus1b4+cJPqgpXRZ2rQrfBq4l6zejyv8pD1D
2qPi6hO83x7uSdvHUKGbRhADoiHV5YCqD86zwLNkWa0ZqrwhYxFomES6XWzBMVU+
4/8BFu4IZTAuCP+7yJHZ9OXh7VqflEJlpf2S7JAwVTJDxF7vySpU3+QhO/WQ1fMk
SO32yEZXEMIElqCDBioXSx7gWXPrBFCA4ZlQV1YJZLknqwV0s/lRCD3KKp4z9g6C
HyXUByzI5o0CmXJBi2NvYl0/mDtJkv3llY2+iQXrcVd6gXOY6OrAAghivZK161yn
dL8hXfqxwYXRBsdLZ4v65pKOZisNf9jOveRSyenST0aGSVUzrdt1xDO3pXheXmqU
kQDFr4pFkMOFTZCfSH/wAlb/s8veNo9Zfqxryu7VBD89zpUtYuq0TwpIqxlt0NFu
L4CnwC+STHKLHvGKueoIXBAaTHLgabiJaNehTN4+mW9HOl7e2iaJETzAl2z/nBOm
VRKHo5Ca6EDbRoHk+ifEDtGwrJwbLNDe8jUlF9zWw69PT2tnfeYBI3o5SsB2gAxH
IZ7NTlz3tMSiqAHaCl08KJYxc9H01FMImeY3JbbYAjL/XV/60bgkCENKlD55Ty/6
Oo0ZbfwHUBqbQO2vOWU7AA==
`pragma protect end_protected
