`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Qiy8tEgjAi7/x96uYoQshsuILZio8kcvmagR+Eu2K/nvs/WFnoalN8y+niIgsUx+
CjCsbFlqAwHIX6K9F7MQwS3ev5p4QUwijl1Gs7M7vR9MmsyiNN4dZn2bgdzJ9Jgc
gcUevFQ5IaDLU/9bvb/n9bUYRdcIfVAAZEIBA1V22hs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27600)
dQTvvfyvcsEkKeS73Sc80oxCTNPSk8yXKTsSY18159grNJV+fySsoOqY8u6on71/
EWfiRsBsIBcBPg5SoyAPeGAeV2HsffN0f15RU+YAYzA/rk6Ok0nJe3GmljoebkZX
tY6mISUAOkCPeEQIQuuIk7x74XXSfJ67Zu6VgBBChScDMQdzQZHf36AFqAlK19DC
COX59Cc2cMqFgjn42Qxhh1xX1iO5Aa4A4ek4kWHCeRzKs+O+ph+2NbSXeU9c5xrY
TGynfSOFCDQqL+uTp4JvFLh2DnuMywDPmdZvsYzxr1EYWUf6WN6cgbVJfOj2dvMv
vGsGJiyuwFL8CFtqUjGMBHhJ30wdz6sXr0hAHiVOMuagiyhjOhdEK9v9qsEMouP0
o7rXXO0M0wVQR5wGnhFb/6xp6fuRhm0Z3VAxOiL4xvSFpjk6NqAHYx5UAHKv4gCF
wyBa/LuKNl4BVZf01fAoCB3VAA0XnEU4OTsQX9uHrVFZU3lmFmfQQlD5BOVbWydW
VJfPbnKToptXm7OKDE3Lug6VRoh4Y1GFULUKxkY2gfIgU4rh7BgUJAZgKHppOu78
aPFpoXBWdJuFRoq3qYud1bMo89VA3dT+su54N/MRT6Dz8vLiBduI62pAcNHyBc+f
qnNSzvZ81gZ+pytF1USf94vmlV8F4nhrMP1oX1+xBiS04s1+QKpSFMG/d3uugmRm
7ebJyBREFRvv+oInQeLoCWHrCJh3Vz1JLLqWD0ylpa1vFsiFiApkSqYS6KzC+bir
y4lcagwrgprJK5xb70RZTGBpwr1W5Qt+QhWB482+zPJesyWyhCheTxRpVrFU8DID
IBuF/nDROJNWFUnj91nhGHswqGvZt/SzTd1ZkKvRw6s6joUbHgpwnmPfyL8K7vby
DPUEyIcg+XeENrQEUB4TcYu3cr3zVPh5iWEnnLtl/qYd05Thh3iCuEf8vRPPkY2B
vMQgzuEMCBqtxsu/7GH0u7xfPAlsV6QROoXgI936/xcYFSD1VQ6LR7pJ/XCHx6/1
nTJ4/PhTrVQNVsDR2nvJLR5q7HMBCkAkf3M6FyUCbQpeKCcLbalppWKGtP/m5yzx
ZynSlbUMNArGO5MNlzeG6FRXXxdIVI96W66KRnEqsNEi7DLG20v+7wYLAHBPYmaR
iLY+uFzEdWSdBUnvbQuvc6U4qBPrM73s/96pfSe0ISl1gSdHAwrAzbNT+WcwCWkI
2WUrnopnaICS92NLPqdG8RVKO6WrCvj1447g5YmGRUVQDwXYdYx9DAa4qILA0laR
9LN2B4O9fhCOC2ooVlyCtQhyRLMIExPPxd7m4j5pFWOYaT3j+EMLm9jl2BQ0sf5H
V/RzCXzpW4JTytDTLXMPQw4MxCRSWU9/uvsFRtQdaOvcF3leK/VZnHnjD6PoZBN0
6+6wGRSA7Be9Jr5MJ/GikWLVaYNxi1/fc/jSxsOXVViavCFUut19zuyRuqm008TK
dKwhId88/ZuQ4u33vvZIk0YHypAuKb//D8ipiLSnOAXMquUNRkGJnyveQqmh1mLr
d6eAuZ4hfzhNQYNzovNqli8w6XHoPdu/tp1o89rnzq40BUyIC312QhK++Zy6fmue
lQ8HhZNCmjZkyYfXCXhpm7VgG2uNwP3tJsobU2PttIYTrfzpqveJmOjyGzf+SlAM
mYfZoJCQQnumLG+5TbpgLdJc81YTczXIwjWiHfb6M8UJ810hL3sG3FP7oz4ovtUd
KnHn3pTvjeorc6fUYoHVNMhpQEt69WGvLDDzLe82Kyi2BQuoBzwORBlWrH4d++DX
/EY0+6b1v6A/AwM2MspMsbF9rPfSInO57Sfb57qffcdbj0cmN+susyaUchl2WUcl
deqBtIEQEJq3hQ1S0TzMqTVTn/e1/EhW+u9vdZFlqhJ+Z/fuHnaJEZdw58IW+V/g
E0DtqBJp3ha6u+14LUCO9cxyHQteWoRweZbZszPwxPllY5YukbRBfjnxc96p7yk1
JCB19lIFcTcOhdkC/RH+oKe3Qsbx2zn5vBsIZwQ6doloV6WZqroD7532zv4OuS2Q
6IIwKkiGEdmKxK4f82bMgHZQ3WAVw+BcZHOK3z5duaKZgkKjn0TsyOw1SGK6muwI
ICpwPNmr6AOBqBkvDbz4Ez40HB3LtOk/xlcTTWW3PXegEkWR/KD39XsXwgD6y6hq
vdzpfC2kw1BSodRCO/JPyRuad2HuuHRg0SI7M7bN9OGCIBgjWCAK9uy0dQBcMdxE
yJtUaqmPs5qUF7h+vsgqp7tBun01zF9fA2UJYKzCGvinm1Qy+I9RPSuGL0Eeqa7A
U/6B/CVsg5WXZimlWaP8ZpoSeRbWWRQbWx5sQhLv+8BImG69MXMUHY1cdU6SjD3n
AWbJjwqG6EVgirthMnPzLZJTq38D85iWexmjqm7sYxiFXV3rARNN81fvupQKjOzG
Oo25OUdlOj4n3LnCoZipm33KMz2wXmVOQtILoFLlpnQcSedMdjlOHifp+1HBCD23
IDaM4C7A+SqI/wW1imSG+5oJ2Q25kJ5kl0I7RiLIQ9jI9jEhKdpGZrGiG2JCbtiY
s1/N548WUxu/hQZP1+ahLoW9mCC36cmjaZOIuSJuMmfZgW25G0q+P1dYelRTWYCT
lePJfWfujDLc9+L9uB6ouA6n5snFmptw61gPQ7mwOOf+6lkdIS49jCYfIaIq78w6
605INc8lknw1sezBNp27r+6aVOQQ1cXNPxqKBHX64PnKbqlE/W/HX3AYu3SUL450
h7sWEorLvDnLZSzXtYmDjHU27SIzzmvncfpJRkMQxmqdRaooo5cj5qKieLDRrZtK
eVKDNekF/sb1jk//tGx3dBE5dBzREQwMvI8jpaGH/Ib0i7NhHoa7fOK8vKIFA8/1
kq4kgPZxTPrnoWloDivHACYkZaBMIn5z9zfC56nWN2HoMtlvq6PFJmfT9dgglo1Q
UZbHFfZtggHyC425aW4hLIXzzOQm+8cuOiUymixzwS1m8J5I2vAh/gj/xEk+b0EU
zZxAdCuAf7bzAWEomQcKQbjtvhpDy+++DXc1y7WhkSDd0UsXbwnPy59RHk79oyum
GU0+/6sQEznLG5gDrU3IIpjN0G8N4W5JQqkO2KlhquBxWGkYb2Ul0KNCl2yiQrR5
1WVimCQdJ8pGIUCWXFN+o/0wT7xlfcG+X0YInUY/XBma0hE9ISYWyEkzqZDBTQIi
Ccr5iOBs4+MHEwyeDr9JjaqKyFVz/+thMUi2EPFqMXH+Ea88vY88SVOXzHGli2kk
nlSIikrDXpWyX33yXEGlKRekVLJ6J9Y4m1arEbtUiw8jSH/FZECd0AIavoGlUOLS
8D+sS/Ch9qIU8z8bxWSJykKou1wwF5nBfETNWVaukcS0j3XN83DmePOhfvb/VTsI
p/8pVElyMicspOanpca3nWqRnbVbsyc9D3c9cm+RcWF8nKcNjSf364Lchl2EEduM
4F7kl0xvjx/SZkjhE2IfnPr8vCZdH2YiQzK/XPrnqyN8SakHjb0HNaa0e695mmzA
erHAu7Xi6aUH+eGQRjeHiVommV+rZH5s6hyK+SJCV/VyBaOkGpKuyrLwMjC8KjXZ
0mf8gfgxzKE9sJcecbj9IDvbJkyE8o17uc5jyBJ9YHAPUaHvFEqz+QsbEoGGdtvK
TtptJJTAOoSawd9rMduguG8lZT6HMeFZZIH8a3Emoi30yX4j4865f1w4PQT74D81
L3hS0fcDe+1ldYsUyASrg5sSP6IlQoWdRp9FmB/wjTuzBriRHbkNoF7L3TK9rLNe
TSqYOroQ7zI8YamXAN7QZpOrlmnNdQDj40fXYTxP4ljvALaw4szUP72jsw5EaJO3
iSvRcMQpvxreB6satTEUkqa/2SrRK4KAQdDcz883DHtXXkQV+4kthHyft9lAzSfc
NRqZJx/XhovMflfAqEAAWCmWd6psTzyXPAJpFK10kZin7IEgLje1iP/a6H6zwcSb
5Pb8crQQI/D3p+QBC3DOpeeQWACJDqRP/wvnaYUTJzF7na1KgasXZq6i0Ia64MNf
5thzcdtdwZAZpQSwgCurNUkjYwXjb4AqFatDtZYyNISwDjF0AhYR4dLifm51Uizd
HBTIKi2x+AMmEqxsUJzQ6NM1gVNIOgooyTIm0M81R9fSo9maPqcFXdxupOGZ7ILJ
Cqe+baPzmpSPfC0BK/202hvtbn6YFvSsXwBzvEv2QORiiH/Jx/hn1ZBKQjcXGR1S
gKDO0spabvRXo8H6ArstmulfP7Tn3jueBXMrAEvIKV+JyQ04dUBCa6CHW/28RsMg
fJrLjTq9LngITkYBqF2arQ3U8boh3RHDRHMQ2wo1LSqUZwFHW0/zvXo964q82LZf
K3Zzpg+UJ8F09QBIpfvOJjqKMMu2xfoiAXM8FRmTFZouZEsMol220PyPkwokzoUl
90QTHHuJX7BUgsUan+78XVRJdaY7YrhB1pchsAy/8s4yt8enB8BBhgezYE7xHbPG
v2/ave0ovEeZIFvUu4k8taMV7IhKIJn6Flfk0KOvi2pRJJX96BIZzYOm+o6mJAUq
Hxkc8UyZofZnoPvN8Te7jZ6YKCTB+sW6j1Ax4B0BsysbJfS3WnWX/xtasumrPiwt
bGFO5q6iWSSifJ5Gc33arMz5ISueW92xBPMkvP6V19WjyI+AI0UvuS4Be/Y9i86g
8hzY6b32inW5EAOOZOdcOPYhMNP5pJ9j20oUs0yp4gwjUdfVuRkw5evGsRyUryEL
rpnx9oVaAeAEjqgLxYP4n2ImC3jBWpND27aTZTHjbqVKJ3Gnds17YyRtWLYztINH
egkA4bQe8JwVEGgODNSZY1c7rhTbFYcONC7+ZAXGWpIR3jG6X7ncAF8z4L0AscAO
lke/g/zcLdpvFaXl2Zv9kANz3yKIBQ/2Zozr/WeQQpUEQ+J1RQTEdwMg07C0nq8P
vetz4SO1pc5zUQOFs4L4v8bkrv2wF687cSkJ1fEpLEbwmKUB4vVlDHCAOmiJB6aI
Nj6FjfGl4gTicdwFbsk/BfTn58VoYgIy025S0pefnV/EvNEsnhrRR564X02YrFME
yDj+5neJxV5bdTf8GA/vPoWlcjlCqIIdJVUkOwwp1DOvY0oRNLLAtKqAmU/OEg0S
hTNRdT+cJqEGpZOPFJW2Y61fdkagUI/IbWUi1OSyzKhIJTUtJAdCj+Ib232bYcrj
1VaUFG+mzXm+4a3DSZWvtSQKPEzxBn27Sv4im03Sue2iI7yW6deRbyvPAqJnQVd7
Lmjl1fkSv3pV+F05Ylwa3MUkkN+EzElTXZKQVubwwthaY7nrCVhWvm4xZ+G4Eq6l
+BzIAZ4hNZx0Q70Gon6ZdGel+akKnNPsGp1BoLUPgKmEzG2WR6TbD8AeM4uz8R38
1Ap1w9hA7DI962JHu/JgbQKvrGQA11zUnk7ZGA1muS9XINCZnR1JnnFYstutEvhg
0F2FztH7SgYGASu/KXCTKBATwJeoj9n5J1JngTRtpHdFf5I1HzluRdmgiyzbA61/
0DcbOSK4fASOTodDb+agFHnrWpOnyT4F+oUxdZghVwMb1V9yNZa/2g2VIUCUyR3G
bh513lyy9C06qGh6KiQrnUsH9Ky9YCf2UjgFDSIgBhidEKIGsbBjloz4ftaSN56N
86jKZiwUN2Uobp0B6pRS5d3Sf3F+ahcfXq+O15LXDJ/zJ+lBpi8UhJw43oH7UDMV
xypUsbD5g5vojgbwV/Wo/Faz3sHYSrsqv8iUymEjfOEbKEtnjGFchAAn0UlKhDPw
IYVbrLrDjioGA0J43m13xinlB2svK8S0N9iZIrFWHUw2alABcESayInk+kC39JQU
NmPn2+o0yYPvInvvGU2X7LFqlMFXzrznsQmBEoBhyZ9Pb99NgLbEtRmaUm5XdyRb
+lbbj4ix1c2v+0J4oMJF39iPKPZMN9dDVxIE9jHcV9U75wvw6JGhHQiSNyI3jZV3
ELtXmsLzCC6QyGF1BJAKgZJGo5er94mGZudT0dphC10cZBSw5lUXLxOPoBjpsVH7
c8nPjR6glz4rQ8luMePPO/9iK84uNrNZJtxsamoBDcueZuxLTcuAJGwN024pplUv
375t/YTwlhS+ybXAJNN9ZYvX1kxFKcNMnEcPcHRbQ8Xs+BRkE76DyQxBoz/uuSf/
ReSKJ/Iisj/xm6419qxPcIa1GFfoyJNlTaEBPaQDwqZJCXcojGwAXDVNkLcFelI+
L/PFry0t01ENEME/CYKnUkn3cQpZAu97KIe2ZIvrJmIgAVN56BfrUHFvCgQfs47l
eiMaiIOgHdtKrnmmAw3YXgkaWUKtzgANhae1FTAzZhLsEVPiagpPDnkr4ZRKMihK
Sb3kUyfUkYi+XpwzyS1RTE25JDWPXXdcFU5snBiY1Fv3leHGuKQoj7aVDF7BH/QB
Rh784y+FpRv0C4aGCHg7CPBP4qATGiUnv0Bdh1ImsqVXCuZ22NSOMjHplsbhyZze
aGh9Ius0U4QOe4kHidgM5xFrSyV6EOYfsVk5z/T8rc1U4c0FF64W4GqY7dMF5P0v
5i/TcsQ7cKVQFvqq1ibec/Y/Qb3/fBTt9aMp2q0160L3z4S3J8q87Ki8tcdAgHXF
rV0AaGD2nYB9MLLmWtZnNN/Tl+Otiup8BE2iUu2WxTJbZ22dFNieiWQmu+P6Q9pu
8wEKsKuoqSNPmIq8wQjIuDivSHS/mu81rbcETa2Nl4cmF+ZDpewGRQPO7cKw9ToY
PlinQ+GIilZ/8qK24EfxCgEpHSVGjyxUk1Toxz6dEuHxyYTBuo5wkaxp85cE1VWF
0lTR+CEepi0y80Ld2BkPa+xwmnXWnaO+jTf8oT7syeF78NotJ9xTMeQs0ntIXpUQ
bJ5qOlvpZvi4efL+3+L5dJ5Y3VnLcLo5JBccg6nXAh4x/yVxWnHyytAMzLJ+H4Ay
CQCSC/vbx7/B4ijNs2PXNlF76uook5W1qwjqaTD3OFIwFI27FkJgYFtJywmN0AAL
+Xq/l0QTf7KoXAwbQzfft/nUS2dP2UWNFgRIZKa0d6/F2IDVSq372aU5gNyjfx6n
GACez4mMbM4kxQZKb6VJIG8Ips5OMSCKOhKNahsQN6fLYWUgAfBQUiYq6AsH7W16
EKR4MUVQQdgsJuKaHJ7GD4VUQ/uZXHxQE/Fw9EB3PI0Anm1VGgKSV/3bOPhBhl6h
gEX2olRrWTAVeYP8cyuP1ALXSg1IYC/FGiYohpYUuLJmFO2RCGRM2+m7ZYCzSNcF
T/39oYRKAqvsAU0L+rCAbzmHjlHzIoRBjl0xFP1eRMpGYJAe3ejYlDHij+c1W/jG
OUpnSQmkxJBven7lmy3mNhXC15ajspZykwqa1diTF3r2QwS99BHor42SHTLgNOG3
usYi7qY9o0+gycIFxf6CNPsfwwxPwbTFTslyAwvICYyFtwPFg7qP6TIjfCNkhxM3
4s/6Mx+A80SLhijshQH7y2ML2gWt1OtRTI8V1bcHgnOmoUJ14oE1bXDUGVHcpFfV
7vktsQ0iUg5E2KbDeHvGkdXsi1vV4Q43EnMqwkiSBxfjrCmZ07STmFdEpV32XVe9
MsET7by4layHoOe/K5fggqL0+V6NuAxmTk7+ZgUe46iZKVkHSuHSWllsNtiJbjmc
Qxq9hrlnawJ8uqf0KWvOMpPx1FQ5B+07FRsbxoUBKcXlp9+aOJ239YptDqeAbIkF
We6NYT60g/KhxbXMJau/gWXjBm7gJ++qiPvfMrv+11TwDqpJ+2yyyYC0M+TFT8JT
SgXn972NXeupZ00+uW5TnF2V4wJyU4XI2JNR/WYuEAH4Av93YvsdF1JP6zVAMYLe
0PiqeREgb43FKFkWU7DUd1iHYO+6r6HocIIEjZsgxY9lG6T9lFSlNKRVsSSznMRS
ipnJ6M2yGkLCBJW2DfXkc69JxmGrsEWW6GAB6RiOwABikq2bGr0PN8KXYSDGgn7w
xY4O2UKmHdJvl9L/lU7TW/RIswTimQi5AGYu2IhpRi+KmrFlUz+d1JVCzfb5MJae
L+bv2mYpnxyCPb0DZANiEkY/VdDoUepsSWIOR1MLzdYoka7SI5sbsCeMH3jriRPU
yhNf9I174V9haVTQn9EK7Aeuz7s7JPegWsmPP03yBpS/DiGq87EaIfdhr3OBWcIA
2za8yoJ19AgNL3upHUMyVP/ONCBmuPKIBmeqxAjy5wg/53DyYWMflc0rO3TqIvml
TBiASC48mQgn6OTJ5k8n8tXKOkOt2iVWTeKMFmhlXRMbHfe4BaazAdVr+pnB5fOV
UW9b15AtBe3zmRbXuiKja20emSaQl+O/HaUahsPOE+Xc3r+ZR1li5fnldcUMc03P
5zQVkLgWEXaqTKiUC4j2czq3wY4gxjuR23Kt33oHiVoKs3fOtkCQ9MFUt6wGsJzM
mMUYuFBTdCbAlyTg9l0nZg43BNbyfh6xNrtlzPngWml9bfUcZozJxT2C++Pstc95
AOetkfFcnvJT7f296NMaXpREH1yoFxrSx99WoR98WRlUdvjwy6AKKzatTk6wdtlY
a5nPll5j5HdSzXy+t2mgYt3hC/IUef4pqvTV62Obvyex/xcL3mEhAjXhmS8M4pJa
A9PjS4LzPBdHuwinYfzotPJnfVolgLZDRkoosKyFoYPNzk/5U+D/rSntuoGZjOEi
AyY8tDmN8ebg18uKcvAV4IWwz/AJHmax187+IZ0Spw6ZOTWa/GIc3OBZCrNgPmx9
NrKhHsr0g5o0WvOVdjpMRSwOfKdOKTsrzNYE3PfcFelU95Lm8GluWS549yG7twMr
aG/0c5cgqfbSnFEiYNY7YQ4L/szfCVpNCKOOz+jPP2TSWHvHdAJytz5vuaHBt5l8
SH2d4tfV57ReBPLq7mowfslaj+IL6C48XFAo2/LFXWSL9UY1OJ8FfL/V7qZTOql7
hjUwKqAjL94rAYn5Sd58P/C4vvH20sdfyo5rywvE0NWWdm+pu6EaUeUkHLMHbBT0
H/afETW7mikvQGSTW7VjK4VPTpIN8w1QcCZs99JRBeM59XHSrW250Xy1YeYRxRXt
+Z1+YOTlleKjdl51kv+2uYV97skK8ZQMhmQECZlmi/+ebYd4+v+M9cK5IHBzgx/E
MtxVkVETyZ2NCdg+RGxH1joBPI8zfEXfz7Kk7QjDx347UHxGcc4yruFhTXo3JELP
EgVbmssFFaz676k8b0QXSqlfSpNvlxW1ZQnYE663hxVPm96+eZFpZvZOAeq4UkYb
/RB//yfIS7YxP3rl3eF0QjApRjGCOTBoQithsaXC8lY2rQHOeJojqERvAWWWzOvQ
ctTIahuMQpOwrNX5hU/YmDKi+eA4KlpJLj9BIIxLKW2KGpgDk4pihpM/cmY7dmz3
cP+p8hRc3H7mxWrIJWjWqagploz+hUUs6g03l7RQeOhm5lQF8yHQwLln6cxNj6gL
l7NV9ehLY5edmRRpYkHjknRspncBcXDzVAcp75DYy5S5mQ1dARZiOIR0LpgV+ghP
hQdB6SgYa2ZJs8NZhqeBYzmckojlXAgh1utm8YJEOVYN4MQuBNmDvO50ejEW6GJ4
YNf+qZbaIXrOgEJRe42BvTgk/0oRI6RHAqVJZLJ9oBHdRX4ePDNs6AT/P2z4Frts
dB3dAShp1fZkXq6u638RZVOoIssJOOd04sKQpeokL0IvzSlAn755Dj8ua+Va2fT+
RWwjVLuE+MV8d33H8F0Ug75on+B6V6kiLgxywUsjr9HNeH0CXWUxWCqF/ODDEEaJ
mID8yf+dw+Uer9IGNXBkUskUii+rDnJ3hwvrr8V7T1jfqs5PnKEzf19DoBiqzDPv
i3LM64OEJl7507r6Ewyo0kVdPqqDHvDD8Vn/JNUa20LyTqlmgkS42uQ5eiHmCUbt
mb4KhCd+njg3Svf8l1g1CNcXGSodRwmF87+CYI3w4hYyFO96L3ju0qmGPLXowVFb
/tRt9+1T5rQbl3tvzcLL1TRfY0B1FBRmsqAJbVBM+4YM9cwUDfXkY/u16P0EV67p
L6n4Uhch4SYxtZMxec8m33Y2bY4Ywgm6hC8fQ06u0rX4tAl9HTwRF4z0ePGWrDlQ
i5hAo5Sq3H8s/1SlYmmykkHBUx5J5L0sruHwpiIuKglHCJBHFgqidWhrwM5/0yq0
4Q8Af0ei+XyaL37RNBYsTApWgt8AfIoFW5k2Glt03c/FdcBdngOCO4iv1RZCYfR6
IgeSzTmeTpMdbSAK+Y0IExw9qskfVHFzlzB3OllGkmgXwfbkrcdEKZX0BRRla31B
ACi91lbE1/6ystr9cFu466gIwxbzLqAxaXwDJCiq3CZcf2vRkwggnp0uITk16B1v
GP0vqFWJV7kEW4ffwAoJ8aiO36KzDQyYyvxSG+mLFT4kqkLpc7aiSmFlpil5GyRL
M8n6/F9VVaL58UGRLiFj6aukKafLXP3/WEd2C8bMjYijtLpSfTJYDZlT5vhelYaf
S6Ali8X1Ga/D+jlX5JXP0LY9Kx51g+nO1dvxVXYBClcFV7LzQV+qTCmhCWaZaNkc
lkJM5MYVvFzOufTqj5C7Z26dSlTegMMt99zKzKirgxdk37p/nA42ECiAsRNrGJdo
P+UigwX1xqOyOspJCMWUExcWjg6OKRE2JtRYOAboqbICN3EwoJ34HNDVX6v+ivqA
g6fY2r27R6ubau9oH7JbLBwe7jkKKDQmGsW2nFjYPfCkfkrMDcUIynpf2+tBddUB
5PBrKEofUsegpmPTnvpzhoIU+Bf5UYn+/aTo9n4lBjSvk34eS8GU1ctn2Q32AQfU
1fRU76P9Xxu9mzzpSRlIubI/PHcnHey+p0pt1FpxTuFM3Y/Oj9ugstzjcpen6/Mn
FDdKb/ieUrx9aSVlOKpZ6Hw+1q0Rv3vLamDg7gOQU7uurxxt4xdyRg4MyrF2gfVL
KyM3mDRBfrIfeE6JnTtnC5IXqFkEkbTzYcY4ZqH2v2rXFzvEIH1A9usaKnPQUGN2
oPy2pRMiMYsgo5SkE+DS14RKpHjQb7XOmKmr0BhnaO9hyNYkxjuDHH5rWd12O6Vv
VU3NPt4MhPiXpUR5qFmZbzYBkPdwILT+OyUf5Dgg2VCpLrvD1H1/DNis/g/h+3Iu
bRiWP/XTYFfgdSde5vo72yAczzJWX6IR1C8Ajn3+B9O5sEF6bo9a9Wlsl9rx/cK3
P8ap6FJgTzX/QoZc2kfKPOam1NT5Lof5Gk1/ultoJ4Ejn3BWYStwDrWMROarm3iG
UoeghroYDlhZ9pZpVpNItmX4usZHM6vMZ7XS74nWLqqJpP977EDT+EeWICrHc6FP
uygbIzhx4QMAtCYgX2xWcW+r+NuolsVAkH+kRcoqIq3HHkMeTDI/lUCyXwek+8Ja
wbIcSQ7+m4IPerMXdZ6CGKjGEL5GPdBhmN1dwZub74wTVj4RQGu20x/LJW5/Snh8
oJZh8Sj6qIIjRpg8H19fcpGTAXzLU0bnoMD5cAF3qYF/sYvIaoebrDJvc+GyFaDQ
Y7Wb2tFAhDhcLNtFmbxcBj9H/tYKAIytB1iea+2AM+tcn+waR5UukQmfOTlPociX
lufm0LWnrSs/T81hWf4ekeKEJ5t7Gp90aIbpn41N+FbJsQT+Jbx8t42j88DOCXyS
6JfvD98F38K8weOPN0eL+VmklVTsUn/7Dy1UWrFiTtsyDxFinVII8sCqXz6ES8vG
W7v0wZFBfqhRSmwu/8stV0yqgQ1j+vRpPsuXgYBCBEuSIk50Q212WghYRdTPtTBL
YMpKCRUbEmgM3pCrrbxEYhgyp3p+34UCsO/zqU6zHAdS9q2+Fe4fnP0Dgh1M/GSO
Y4260AduAbhj4U1EUZIaucY4l4J0IUr4s49g93vqyLKbiHZ6CRyQACBkH7OXX9TQ
PofDVdASnklwcZPlmwQ9SGY1sg//uV+69yA3ICAQ0igXODsv9+K/FZRk4A+jML2S
GyXWcDPfg7OGCIbZPLZH20MAiKyHxiuhJveKuU4oxtgQPRLG+9VLSENjMfhx2cuY
4BBEEUjYpz2TNdlOrO3/rUJpv+Kq6OulzPMpS5wcOxFcpTjfRLQIIC/aSOJkmVv+
naP6X0Tb3xU6GOIMvwkrx0SrsKdbOGk/EHmQt0XuNCaJCin3ENVjWy52nf3I5eEf
KWUxNlUN/GsSc1zU52tL/Zt1jYq77trMojKsXIiKCYO4HBlNHk/2/hQyfEkXQaVM
GPoNvA23SSMA6WCHiugUH952V8HglIF9+EYJwOOWO2LqSlgB3UEi7C31es37ffiL
te52QWEXgfyvoRjFW1xUGdyvVQizUMQNcDfYaDq5IS8yLQ4X8rJzQ8okNGtncmF3
T5Qh2RMd0QBSIEGp/KzcYUzPFGywllWHgMvHK6j2BTAUL+2V5DAwLElNcOT3tk+s
e4QBJ35MItaZNvLSqp5kYrdz3381vCB2ObJPEqNYw4qan0dnIEmoYkcC6x+EyTkF
uUlJrdPDlTyXnlvqbcJI/fu9MP6M5Rmm29yKTMxqWD9d+dzIATLM4HCQRaPjmpPw
xaXC1Rg/FKewlJMcJk1u8u7rupGeZw5ROqZDso0C2ja59K0tDQDm3dVnvQGVAGAs
yQ5UT/2Os/V2H+AoLpXp9zvFFJcTu2ETfLYB1rO0fvvJ7zN+AYke/ebDdLIZl81a
d7nnjCMhHAqGZHEEBQYdGeNDNvI7XsI4yZklnMXt7U9i4oJwQT2w5zj6wj8TS+tX
7gDIhr5P+4YriD9VG28haOHpNL73sC8kzFUPWWYCQQcsz6vHXPBoy704ftBhfMzR
lshiux+wlFlcGf2RKiMIhipXtblFU0TKICuLI7mAhrmGTrG9YDOKU4cngIJzCCUg
UNqjWyPFg0TKtA32Or62em8Ya6iX3zcK37uE5C7AlGTACZEJ/6/AmIqMKRAoNcWF
U0wsr+9TyWOmL4bFtfG290EZwn/ORFiY9SNYWXgP57mbJovRq2KiuCsqoBqH1M+7
pTeKquJ0pLBkjkuiXVtuqMo226OZ4q3XV8nQtBaiAi3ah+F5nOsK+D8SkMlSKiQl
tekKTVLe8sQK9PZC1lKiA8mjvZAEYEIXPAOzKHbBVDrmyWnruiFPUlCvasfX8gnU
VXLrBY+m48BFdy1Zg7kEqSiaJIOCgZbQ7t1sYLQQ9Tp5mYiBK3mBAS8affpSCG/x
929DMDeJnHlpavjlN3NlflK9kHa0aNxciSoa3egZdDA0aKdr7e61qOA+zRcYoufI
d16Iak7IIBZJVtEZoJBhYDcWBlYE4GC6WRwdW3Dh1a8K8WkX3M0JRjnLPz6Ga9NT
yvxzTCSvBaW931c5RO+ZU9tIZnaeGieVc8FckbwzEcpSDn31NegPWWNixiG2F/+D
BrvqsAGE4BODDDKM+n52HNn2EHUf0qBQsU+QPvbLnjNfAPTNhNmaTUyAaB6kQgET
GMfkyMMxMh1BtQaiYnggZMm/irdY8F9gbBCNw5WNAVt7MLHYYkxwhrFbjvfZYA8Q
qLKTSsPbK3n4v89i0qloGNIcg5LTTyabWKRNX2GyoWRp2ZqPlEwdthiMt49dvU8Y
Q7hCpeLBt/6UTqcxlJFeSTMiuwPCkEOcD4LxnLt8wVIJc7v4I304TVQ3Nwc/OJQh
qu4dfTRF/hh/co4oyCW632qv25KqSaLgbPzFDqSSuQO+y8FXWrCXKe2j9jxtpaAT
U+h+UqTeNzZc3n1EJ94dUbAtKLey29kRzhihMsrtA3lKHiN96GhVjuDXmAppS3ab
weCtT3FMpPjcMGcpuQmAshEqb//otLYlA12steTld01eYMcFomZ8XwOQyR7C+oKE
p/d1ja7wMuXmqA7t60VHI7OLDgAbNeKCXcP6XGJT/yWXiR5fIZQ55fRxlKVUGri4
xrTRyGk5POWU4ovJrcw4x6I6HzHRqRIcOsavktK68376UQBoSasUcqg+I99grO2S
KwojWpIb7436FVAEXX/uPqpjosc6hiyoYgVMBlVR/M8mGUU1iXMljHHVW4BXy4gf
nXT+wQLvJ0VCan+tM9YoCf9LwjZYOrVw/DjVpXy4k5qq845yjNNDXFczLfhBK8hJ
eMZOyGKeprwR8DrFXOl69q1Eisd0qcDZyKDF+FDSqvQIlH+ybKffaBmASH+alsrc
1zyp/QWgu8AQXL9yXJWv52UgejOwKMoDdghjArzAyeX4VGLo9PhPQCKWdiraqF1G
HC1EOrGmiXNuqq7m5+e5fdsM3DDPAkvhNY4HBiSvLMuHI4+ImHkouQ3RLKOH+YLi
v5WdLD9LnOJYXuCb0hJOP6mMoBHeMD60xslne3bzICVibENhiowb/AS4x03gHuE/
SQkGXHMJdFKf5O7tpKaJ4RnAfEYnVmOZR8dPrTGeGYqHx1Vit8GG9ekt3mmS3Un8
ugL7ROWjKlrVdifbVnK8fzmiXm7n3vhAxp9Avjrf6Rh6aLQcz/6iGzj+L3ES6I/p
sBjCQxgmYm0TG/3+U6OjIXmYJjwH51qPhgmsB8OqePM7km/TsiTPl7VerfAmSYEo
doLi+16mBX5YKEHVvv1g2mh77EJ9eAq+moPLP76bLBE6f7ZD3h7KIQ53MHB3T1CN
s/phLtJ9OlC72YWbhqI6MNuOKcTf0oT5M4QADI5KZwbuFZRUmCD2FhFm8C0pBf3Y
eqDwS6j4ls8G39x/aB7TXe6t7NoJAx8Umukcdx9Z8n3SJXhxx/7ensxhh2hwsCKk
01tEZJI9RmAHDKezf6qoej3SGC6o34Nkv8tviy5/usCSTx7ToG5G8cUdeQGDoFWy
e39C87nLtz2GiO1MSuTspqveZuaKzes6QeTHqWK/U+ocF4lVTz/fW5GCbHK9foAt
iOAxTNLXaOqQrAFFpY6fzGawOUbn8t3g09CTw9lAzlJO5yDI9PXN7nDZCaDy5Llt
qS08pdFGKvvX0Yes8S2rhdP9OQHhjzsMlSxZICLvE5Py3k/ghRAzF9JNS4Hgu9RZ
h/pjIYzSxti6kU2ZI/eHaVLPO6I1XZhPKqLYeflOK2CWdDMUjRzUlkXMwcvL6uU3
GBn3G9CK/zGDerQyVm8DmHM7Drj7muFpgta9r8jInA98QDUw3p6SyWBQKKgldNu9
OmIEYgH57ODJdRymt32wy1VyGxqiAmeTB5ySAGyVPoN8NpTnQapudCfY1Ah8sXHY
yD2n00nW2s8u5qB5oBlwGlBeBM3EOZ/MCraww8GYnaaAxOf1obWzIrFP5aUPwWDp
Uc+dHu7AmzDqDH4IEHx+AZ/eA4J8BmI7f70WBHoMph9GyOlGGIytvnX73wYjepMM
Ua9NSz86jNf2Uu6ZoKpLtIHFfmkhzivniGuaOSzYDwxKuOEcNVaqEH6NljhhP2/7
Mp/zdQ2Ew7qcQaywsBUmSHxj/hJPQG2GjgWaRRaWzWHftSTX2TX9DJE8/4FYqr0W
g6eByVeQpaK3+35dITKv7IImVdvAhtTgagFBiczVTog7iPHgMcPcs7GMejDPlfz1
3DLWmRsGhgrboUKH5kcaZ5YHbuxqkB3BIM3rdPN8Y9/Y4aT6/xfpzKWENHZfy+qN
Q1+MJzxLOfcVtoayApxho2vb31duO/soeAUAo3AfQY70MtD1LCClRfsuJ81+jZrQ
WsDXhLBDkoDgEO5Um8JF9s5kR3ZQmp7/DjPF7S+xpMTgSRcDKMAIo4zNko8t1imn
Z7iq8+0aIV07MHS5bLloJXBezHeVf8ZnuRIwEQx6BzUQTzQz59XxTRrzbp+x0KEs
M7uSIlCKXHPyd6pSOTTg8KjXse+kPyNSDhNNbtvvqB4ZcfTFensKczgtt/l0+M91
mvZ+wuQ5lghZ86g9g9qxE1i3wMblIXz7Fy/W2wyUIbjRV+mvRgje2u/xNWvnrqVs
75OYG9QAaVahyzZrAiXl4BfWgbBii8yIn4++gknunoWPn2BPWZpYnZMzjVQK5YsN
Y8CFJCdfxGTDzlsk0OQyNO1s5tmk7+pFGdLsV6GRlZRjekt1x6W1VMUPgleFGYOQ
BfQbEmXyIMdWxceWH6oK8zPED8/kL1j38ygNaeREV/7xtCaWKSjoKnSOvZ3tw/yy
JeXSqRQOevCRTMKWDfW5TB98bHcKchVjFlpz71gvtMVST/IiL1679TxURoR4s07q
A7HfFCHPhJAMUQHvF1WWiZwm0buEIAL5bXIkmtuKKVfAuF/7yyx8w6EsS/zTqGiq
en8t5+MtyzCpctuMjA6dJmcnFXZtO/ayTTIbr5aXfBn37cRleflCPDTheNsJ6AYE
UtvqRG0MgY+f0J7w5wEHGS4zmBYk+rfnmaDbu6dLnMQrmm86EKx8yIjYry8VRIiO
MXuPR1TNGMcX+Hk6o5TlxRcekJtHG76TLJ1lSsOEH19rkv7OnymMM6wq0L/qI9rn
vPfJsIPwnYt0FO36lqQCMq5HIGKp3aBiLD5jo6LjOasyCOo7DVOnPvJozLetz5rh
Qaw6uLzrAq/6gcvNkYin6O+M6gp80N6h52Wm3GyLaGU0eJ4BJzspDqFKnUjRib0t
nHyVEbHiUo2py45RDHYW6wb8NX5+wEf2TYugiOI32m35DwDXsj2N7wOGAZaNW+NB
A5w4vP3Jx2nzBqOgH+z/laiT0WcCNd3y4ahGn1nE2kGxHkK3YA43tZRpsGRB1tSS
80iAOnBqIt16+SSEwgDL/Cc14oDBWlJLdM7Q1c/LqScMTR9hoGcJaTCerghd0OHD
htn6DSeb/+TCAWP5plCqUkOasFVIxU4kSkB9Xnu9NYxDBE66L0YbEWXuwTftpr9Q
xcKUfL3MX0b0z5g2YVXmxtE4fHjqXiE7jl29g8f7VznjTmU9TlDCDRVHHgJXNghw
c0NhmGqvOKKNcNJdKh8tVuXidhFkzarnHa+a8w9y//cZomD8BOLd0ZJ4zBmG3vPG
EXkDEWavSROdmXol6cHWfwXbBlajBNb3PDU4iupPneZRDkl6+mR2QQfTSG/ZhxiS
pf7Gt3lW3LrHSh4trsC1/ji7gMkdwwczlcZvnZS4CAS5Di4KwShiU1aLH1o4KLyp
H3AEpfRPJaEAXA4n5qjEuFkxg9DE5PIJnDUxCB0oCNFGg8KTz16Q/q8mmE4JbWtL
HLJ6u9An0r4M9H9W1wErldp1a5KBx3bibTz0ceEVD0/O2UpPTI8j1xgT1700qFnW
+bPHb535SwTWGyjhF5MDrZsZsXCXopP/XZa7Qux6Lkh3dUdOG6Oj9Y/xEAc9D9kY
Tu46ZoV2C5XUG+p3oh457zYU+nhaHd7aAqR5U8f/JdeReDKOAUY+MjsaBkvQfiEt
90eOsE3/sCdBEOlBiHSe6CvRf2BNqV5SMkpS+00z2lkVLSOXHy69/RUJI9DPeZ/z
hxFctpr3MpXtvsQk+F8ujnAw7fteHa1k3UkRxD/51eVp3yPtTTiC+uwyIhlow3RA
cfGERyXZEVKdASMaS9J6NTAgtHlF/meWxspY7L7P9tBAtT1CCAHEZbO5tuqocoSY
/L3c79PDsfNOl+SKffc0tgKWVC20OydCcRg0XGWcdEibDdHvU7SovQhptnjS84RW
vc3cSdoGTus/Zs09vs74RcmDm2SirFjswPtdq0dpBqDadK3TPSRFmN2T08K2/cOg
xeAFNL6//bEfQKghQan07RUUkPqZygdxfDTx43Q7jzdkQWLrzPO8ZHQoknX16lcA
ShlQGeF015OKOKfjO1is5bQjFhD8YbWWTOmD6H4qCoeU5tTocbK9uHDVRSNkiL6Q
cBYWpZ90tsSwQGeiO+FZW8OBYyXo1ZjQlnWDat/nZicGofmTRQRLWFdAZBRrD3ss
21bNjVvI6U4HCDBEgQGDFOu8LNJ7gZkxqhX+p8opcputJ59I4SKaNV4aTD6PuOT3
ZNKerGCgK0TGPu1NbJMrptDKl0U0Evmmy5fDGgzA0vvN8Sm7Ull3aI+PO812s2Bq
s8nWgYU3U/hdxgIZwVWkSYApOcSUYWkwzwTi4QOvzFq2lqsadGBxsCnPyPcLrQrV
3Lx6gSPzKKtf8NuN3iq8nIbja2OXudGHTuh/Kbl7VJ4MXEqIOzAa+l8ASFDLMddy
t8xyleNA5aM5cw9VV11KeFPJZ2ys8QXwB4ygY+xMycp9pSt8MNA8b7W4uPk94tWh
4MibCwMBJNQggdVXVfD1mkjWFH3ew9eOXvyvZ5FYCC49KercojZDdDNIKzhrK9P0
bMm1MlTbgI6+zCSk94+RSF1Vw8xYO4YxH98DbOJI0u+o8ClB5wfYzz/NaZcTWtC4
/dy6k6o56xrg9kFxKFARTvyR2JcYD99Kncoz/sEOsCjxL+txaaFDzt6HMsbc6TaK
uxrx2/5zn/l4PNUXAvN4U+WwoKj5UuaScNmTwDvoEVITCc0yV5Gw0gVqds05oalp
jnwSG6R988nWGo5zImhX31vxIk3VVgtBCnHhsV7DmLVNAQjpzmzu5DZW4vqrmVzA
qMZTQkuRGHT0h+MphIRT/We3X2ri6zFXVTqjbh1efw0ICZdNof0tWb1UUaah0lKh
ZW4q6/VAT9LOdo8RuUao2NgQzQS9UOX62b7PfpopJMOUMKIJVVzjEDE8qxS3c+6G
JWABU6XJLIQkj7awsssUjrb9ySYBCj0QzcLj49Wz1iL/4ICtM/W2C/7s20M75fdV
DSgjG3lBGc6sziXSRjigOSYcgDOO2djwf1aejYUJRCpPMJgmLd4s8Gq8n1D39lQ4
MXX5RVsVopJXA45alKhKkbhZWy4O4uLUT37M3UaAL/NQ/pgQpzpgKULfDxo0xPCj
Zwk+m+fChvCIZukzYban2Ag4QrVWkLk0O2KIrBQdb3nZ/HcicpJlrHQc6YTML3+B
AufuWBj1YhR/yAPyitVEz3NyCoEZmkoBSYQIDYa7uQb7fMBY8pTLNjfpXzorvi9U
jB8uf4wMpYqRJV3F3q1BkGUKHpcWklnrt88CDD4GNxCDEy6vCN8v39NT2zgiWk9U
4LBXcxQ/ZlSZma1HDZDe2f9UY/J0uaGUp4pB2WHR8UgWasFbWk7Ncqu4JCSACorY
n0qFt/RKVcvB+u1jjEA37WxKW6Mpxx/JOvs0aOiRD20ZM3RzpOoca+GYm4qPCjsi
A3oUamHdxEbnaAdZDNI+UtsbbbjctJ+RH1J6MeClgFYV5X82hURo+kp3nSfqnJQQ
hrbV65AKk4r/L9wvQYlUJsTDAVwQtw/Dx/a/r+f21aOLqoW4MSffJ+XAholKd/le
0mABse1v7OXw3cJjIMiC66h4UEP8nARupLgG9GAFw5yLMVc27QPG0MK/nMTmCNPA
ysa6kAMI1DYB14yg5+4Megbim8i0Enl6dG6a4WYSjvFJkaGdTCO3RuY+OCdvypXw
rkh5tjSJeX5C8gzn+SL7VJ0XbpQQUUx7zJ85jo/x8HpAS1yJvtO0qGS1BVALQ/S3
Y7lxW2ClhF5oQNYCBWaVieLZCGWilabuviTGkFlej14ChIsmRod8lbY6tg3LZKJL
4QQDkF72GeUPWtY0+f3nXd0lCJCXULMWvM8ubgkWydjKv0DsQuf0y8J6YdUnJKGB
CqH/WfUolP80nVCzZ82jUq49fxqZ4sQx1IMWrZSSZv+eJs2QXYGkOZ14cg93JI8n
QtCAJy0AANgC6HaFxTJxKpNTzxKqiqCWUjfnNRCPk0B7b2inN0ljCVYDp+we9sdd
0mwMJCspbjFKB8BX3Kc1nIJ6QruHyQbeXiPAN2KdLxEzEuhAJbYrW6dCvY2H9ymn
9gu2TQcDmfZ4OkB6yrX2+JBI2mVH4jpLN4HeUj+3L4NUTKN9wtMwnfyL8sy+2u+r
uYPiGfXkNyCFHvYz5pU8/EBznYU1bsW96ozEF5uhiSlghak4cmHWHOJNAvCnlHoY
7FO0ohDoPessbq4QLxR0ynBSVbIyheeVJ13cvV4b+MYX8wZ1C5yT3pw8WWv/Wo3C
uf190TQYLEKBc0E+VKW59CB2S1CZc53CsVAS8RfIilX+D4V1tDrDJSeLVaX+yAqG
JuTXXisLj3Q7GwxxXytaxCHShGwQ6yI0Em0p8T5qsRfXcJNlsbfYaiHZVv8cb6Pk
MOlOXAp6GW6lFUz+UMTPqe097vn5ZQ4jjMzkyZ0ycYDnvIUON32L631u6Wh+g7Mm
Lhd5TO27MG38/CEG7NCR06td1mlnsX/0XFRGUwpCDIhQE5KINkreyZzWJmGPYhYB
yvOX9E4ws47p3C6ourX3B3O1HiCOpat79vxKbFTeMD3uTr07YU2Qb5PVbm01osEW
7Jz+xzQ6hTu23awIRoevQKZ6lbfYm8lrGp795jOqO6dTMsiwWY9dmhTU72VhLJY0
ZGml2nmMYnt5cWibOFCOsa52CFUSMqbVIPU3Dwd8wgbmZKgu60cKlQ47pQU+bF6e
lgpp5Jn6UYlp2MG56kOeaBbSNsTMXDrxz6JDrrysIZFJFWTHo4aGH+TM6qDOfkgI
JiSDslf4+S2AiVEtkwzJGqHbFm6TYdTqCwWonZxklkRqL6eoudn5ovLi1/yqflAt
kRD6KO3tFa3/QGKMndMZdowvoCX4syIcCp232vrOlGVl7UzaPbZ48gP9g8Kgg8Bm
Zho7T3YgEbyKW8RsVbob9FHRaAJY6hAjq9hVRuVj3CgE1L6oVx93dolJj9BcGMjQ
wBdsvR6jMVPfAFA+9mPMWpj1xEUUtiPjuvae2ps2t+yOCvxhhXaBqlUZoPSfxwQN
6o/SiGtG8Kl6ILa+Ju4JbzEPWRTTwGioHJ0I3YlP9oQ1udgbumUBFedURpCsOV9d
H5eUrsvu5Mb3u1iBUDKPAEu/28TbYK58hEI1HBXJESySPMnPTodMEFb1vaQkpz5M
7/n3vxvxa6qJjBuPyCMm01fo2RbzoEiHVK6b55RnKiGqhu5Cu5Qf/bNDkreZ9EIX
k6e2SPVTEmYeosxMHe2/knjBvfrRI3FZdIwl4rXC4InC2eJUFW6ti/XxF9E4CWMF
KTyjmoqQl0qM5Lv8H/xAIqK5oX/764KtiU7SdQI+GX2y7/UAfgPm9mR4Mh9EGkyP
SOXqfCotiF0xquPhK+VQ1w499q8LRiE22NQ0QZtmGUh3T+Y1IjdgDzQn5++j3Xbf
GqLeKxGdcUufCBTGrl1/rcjl48fDqxOfynG/NQoRkGXBQxsj7d/slnDQ24TfuVjv
6B5gk7XlGAyMjn9BomgNm6h63CbVq8SFkXvcJbtWuCSZ0y+ULNgJVMVdP0asly/J
Gsei2ovABOA3SlWspg146lg8YuRPUB4O9R9aQAioAgjh1pw8E5HQUmjmCM+kTbnZ
LJSR5RniWTuQmkZHH7zVuvaGlTA0Uyk/0EFwjUdpfgvcDNT58qYojQnnn5mnOsrC
kG/B2ZOF9hU77BMOOPewe90DKR6Gk/nNC4fT3LL8ohD1hJy4WvcUiz1O/wtDVmWN
j5MxXSGnjigteUaHsPMa9DLMGqiLwJQJpjf/wrDUV1is4rxpaXkly803kZT/5DYb
lmq0lUeKs54WlM3SYFTCAXq5nuX3rWr/+9WOyrviCEAI0fedYek5ONdtCuN/hJ6I
d+A0MnzcQLC/1wKaVZkEcCqu5kCW3D4dq1j1ko8inXjKzuGgUiy9Uopx9Ek9s59e
MqRN+SjNKeF7e+PFEeqJOt/pi9CS7Bnc5IsaxD3ooja0oefG7kq6xOYAifNvd7JO
cMqd+g8tt0wVxAhWJZs6Pec3q8Dk/TQBtjhlTTHVFO9Mr+hIr4Mtc0iSkKRNh3KB
sb6zjrEapMLPvGyZ8YYMyyXoanc0LVeNHN0Th87hMPDitOuIGR2vbnHvd16RdbuJ
53B8qh/76bGsEFs8GJMhNBI0Dw+6p9lCGzOX1DTYrw+tXcpiBL48jQ/uo0Emkj6u
mATbWZEeDBfQGQ4+LvUdZM8DDou+KAV3AXUeSi2Y7TNgFtYggPFkbm990fhpsd6/
gCKhI9YdgYx/gDtPQRNwINeqBQT03P/WsoxrDKppz6p+A5lzI70d+YzRDnH/pPOl
dE79YTENZbdL44ixpP+JU34V8oNYHySYXmoTuJyi/8xL8aayXfsdnKo/W9Q7zmag
xzdxpQ0Q9yyg2I67oDNa8fg6eHteYYpm5IhC8aPnrjoSqfpfwo5cr5tGqeFxkEs9
DcQRCABrtaXDHDpqpvZhcVyLvGc9YAZ3tC6EPZinDuoAJKNfFKf22eofpYuj0Gc3
eO9ynCdpVf3nkSq0pNLR2wLE0ziWqUB1LBZ02CxLIejqZld3Y6D/u7UQCVod2Yz4
dDClPfXfIpu170Znx1yHuDVrAVHfh41mv1h7dW0FGjk3bmrYxekHLC21cT9fe31Y
YHA/la2edlYVKaVhovN9LW0F9m7+x8zH5upbVdxpNHbwQz1YTBJZk6GmJAfmj6sK
LI8iuL/U8f8+OYPmS+v6I3bKD7eFswNTqzfWg5Gr233ns+2i9ryO9HucjkVzCyOr
TdQAU21V4zWYZ/hGU9eVvje64FuwusyzG7aJruVDhP30PLennGxKsKnIFhOzFa+w
gOJJEsnfL/EnpDmZUIO0l/ijkxnWdvO1CSw/87VOzFEGwSg12HvXt/wH3QuLPI4D
4GLqpgSPd+FSqcsHfG4QiMaE26lUZ65I2UEMjov3BEEx19cCamv56ZKagzFOQ9Ri
/Z2ekm/95S1hL1ryo/E2zzPtgkRB8BAO+4Z+9Z/01i2nghKj8/wTVfILQL1K2Shz
Q6FdxHNzRQTkrnzAXlzJLjz6KJJFoeDUiUbGFGwLiGSozYlKsQdvh20Gr7rBjX9q
dWbrj8NWnWqO39FbOQQj5l+wXIzrPsVRqIJfi8mOvsjd2B/a8x1lPoc/tEvB8hsK
A8/zyL76K5dMz3VFJGA9c+AzEQ7vr+LLJDPl2pHzMucRtC6kpkIjOcu9ZLHixj3l
ATg9yMDMlyT4hN85uRwQ+yRl5EOHH3g5RBfaeg7zERX3alEn50L06vpOyndQcBoa
M4KDsHt1sdj3txmSx8y/cA0gFZMnc7CbSeT646JQxDi1UQrqIMx0XdWud1oHPIZ7
eahHTf+i7SvuWFrQa3SFm/jlKBxsGP4wMqnVdFtUtm2qKNvOdhBTmbmY2KIYOvYc
SGvun/KM/keIjaJ16mHAK8KA3iQrvFW8Ircu+9rHGGAUAlz5VMsD/WTO8iu1ll8n
rkidFbaglCiUl2L0DFauf3CWVWA+yeY/Q3LVnpIlkOefOf874dca3DgGiHAJWjDY
BWDxUGce1Oem06MDyEXJMxwp7S/qWRXLCcsmlOcWGoO1z6f9LMSdTex3/2Fx5I6g
OLzXtR4zPQ08t6ilTpoo9YBCfGCUmF4PGiH7KSGrLxApOlZZ5e7u3hX62zxp6xVY
n8nY3FUnEyPwIbuuGv0USZxorkXl7yX7ZaV/+OBAP/5w8G0YhNdRO1b83PRTtTC+
D0/RpynmR/mNFwp40IW8G46ZgD4ulNezyikXUazy4rvCR0tHPSX8YVQHqTpG4jYN
HOtv23rvD7UCjVvtj60SP6f5DAWwcR/sxAIQvIgMmL2vEJV709R5Nl0wvAqL2CMZ
gOCVKhT3umjTLld9tNMAxBGz4QpDzHLs99c0Kfl9pm3oV+E64jge80F7kA/QZv8Y
VG5OtVmyQFtbn5Z0wZyzfS+B6hX11+z6YILCdbQxxFzcVy9Ztu33K6f1urDzDb89
6jKiI24vMOKnK/PewF1Ltal8OvheULfYgOYn/jM6UiZEIaQE0E0JTceBDrxX3jdt
kZkNa8gf2Y6vS7MVgBP0uUHuX+B43IsEJ79RXnJrtvJHiPobsuvdYWhl6eo14Yxl
gfuPeP46YjH6PYrvSXZnJBWLUMvYLUnhFpApdDVlNZfCsq8mE6hHU9hGpRzpJb1D
w0p6/9OmH9iPG6eIyr9wedKWVIoiJFl3l4MEkbSeiKA5VgP+KJrJU+d+LB60orcR
7vQzVTi+2fxpzITO+XgtK8Iwm5FHJPUPN+4A8wivPEwBzkqHv1/0IE786uzWfsGP
d2qdow/taykmsbubd8rbPFjOhkMjhyStUpiPrdSfWj4SzG7k1A6uiUdSTyv6Ce07
6mrmB6aGr/IyMnVJ6mTCDEakCEdjkkZAiLTBhJShHaAMEDuLnHALvGJIVLLs3P0d
ay2EwMtChb9UaaZBVXXeNJKAiPhGprhG4KTu0OLUYehDkTGJXkWT3mQzKg2mwaS1
RCs4AnHU1C5rMWfVyihT0XuzqMmhFu39SDhjvvr0l2wlXwxX1nfEeC69EEI5yl7x
Y+CHGTk8dnCdMMjxZaEP1LPISljS1ehoa27D/77XI+D6ere/k2vB00GbuHNqK+8P
xxsF85SxPVSrn2OJ8PxqG+SFoysMrqGxtYQNDC3uWbl0hP1VdckDsIlDDe6fCXJp
eyYPbggZHMxsqTYxuxa/NPyPcGWADClbvbU8TU9lXa4fHggGUkj7P2AdmCUYMbBb
rI0VAq5XszKzCQZbUB8yqps7MLYS6mdAF5KoDqPYDEzTa4Wg2L1n3RoIFywTgoXF
I9bttc/y0eTObvEwOwnZVZWgTY/B/l2hrOidpW+coBwCLZzMM0Ld2TXbdF+gofPi
+RDu9KcziqUSLmERJx5nBZGucnAscAMDYXNoJaz+1f+4PCBzxj0YnYmPbG5piBYr
eb2JBoi3KRbc2kAu/GmEb5pMcJSX3Tnm4/tYbKX2unOxzijnFt0PHR/5GS6JoHjy
GcPydUXwY+jDnLnAk3iuIGgMpLT+O5hwHZsRG9X2a3/pUg0K0eGcvc57DJnWX/Sc
7zylR0GZS0cfgx2fx5W9RKvnlJBfrqlGdbrI9bBMc2Jh2m7lPSTwN08o5JR9b6LK
Aypn9EbeGnagvRyAeAMaZiNZx1RCXHFR1tRRBOCnBkCRASN/DckueSBn7sU87fE7
DX+TpAXTVM/Od6tpnonKHHUaO6jXJWUSrVSL23vz73jp7z8YowexiP6iFaSN404J
G+wpNki8fsbTfmX+0YmhCEpGubMeHFXLmjCH/LG5lzkh4Bcjv7UuaSLHhuH2kRUS
CYaTKzpi3sqnoMiVofR625ZWau+T1IbodQna0GhjwHWV/A4BQg6gHjQ68JU1xpUA
QIR3H0xkT6tFbgcmxWYXxqXz0wPjp19gCal7S2L2yzAbsfJBMXxVCmk0LBEn7UQw
5hr0Onnk7f0DCchuevji83yXJaZIuk+YxuIfuf0ph6KNMkOO7LjBqDcJVHIURtxW
XyylNqxJCcDuQkZyraOAJvb+8UG3/WeHcYBw5+URQss5+pv3tyFqfBeKE+jWjmek
Q/6sgy5MV21i1R2bxN3HN/SYpgHtRDiosFeVuiuY6PrNqLZqVXwzRSAB/GL22Y45
78Kpha2lP+o6eMqDn+Q63k1/64IZCdpQogHgnxoO++VVpZ9wqVhjqZJjNLQU7j4T
nEsTBRqV5s9ZA4aWfODWVp6Y0eITxeximnBkgTT5YN6F1Dqxb5KIQDKxEVemMADC
F9MHC8ydt/z15txjn3ZYEZJHUA0gcykpZ5tIJMXpyJaNHl2Rk6grLAIDc94srSbu
0uAjKHmuwNsx9YGnPATPmnvdpmIOC48Px+f4PpN63HG3f80jn624hixX7u0UyNSa
aLEj52c3XN6i+ZoPKDmdWknIe16Fmf7PjdiMifBXF0XboZySQLWZR3BKnYHitE1m
GkloPuDhr2TvWGCeM8ISZDNymjx6O3tgTtcWIQ0nk64NQXToWRCgD1Ezasmz7mZy
ow4UZsOs3+XRbdGroFXoa4E2gAGbrUEQYitdm5mp0Gr4Fj6xyXcBsOSiYOgI6Qow
pWJj7dbwZPj001rbrH8bTQBu7lwdoXAH4sVdS8+NjKbgcsrxYudaczSm+8uW98v4
mx4TcMjK+6EL3Mft4zaYlcIvo5JnKGTFHZa594mGpn9rIg00cE2yLR0dEOzSG3xE
DJEFps3n8MxR+rgBOy5eLoBgUNt36Cgp+Pin812nEadT45DU2/YRNXOzZR6/SoN4
Dc6IhampXf8HlmrMX2xXilYLmCVX4NWNhioi6t0UmSXmaG8pEkKAxt3R2YgVidwJ
lcx3As9MsPVfNnrSub2vEOlyl/YDR2ThAAX6j5gqomvFpQ8pZwNFQZRa+T5FxD/d
eBQvu3H7qjurF9XyQw4R7pwMbeI7vn99sQz84zpslARhvpVdur+WY/3+63mZxsGH
0C2YZtYknjBlgSsFlkalDXFu7KwDG8xZVE4WM8fTRpHt0jtiAZUJKei1+ncfI+gN
GkB1JbT0jTz1w1gSHK6YQgLw8oDU8OoGcZZ+YiqsReAzvolyjfwD5VYpSbaHyVZL
cXGU3MbIG7bCt0enZCeUL/DkLui6nu07NCUhnnb0rKHuV1gBHSOPNrUMDoWz4uyj
CWUHBLeVKkuUsoNLxrVWrMh86UpCQBy+5fw6GMwHMiseMzqj7OJ7YG8TmOuwWKmB
46j3BdQqU9fl4cTkmIfMGkMs3LtslSU4gyabj9QDWsfXuPRg5tJaQNFLC4GULc/0
G0r4sgjx+kRz3ayymICQmUNcNRU7QoofQvDqaeMLufuUz0YS+ZACU1hMXas6j09h
Y1FckiyusFsBUPXd/Vc7VQHkLc698uwU+jiMOIPyD+ce6NKfyuKyHMnY1BktgeiA
e+3EY/EGxFjguv5vko8TwaNpYn7jmDFSIXMuHX6nx8kNADe1mY5PpwSFV4Smq99d
xgoFQLgTNpZGtovP7WDyi76CfsfnGc5VODSgmNC7Rvf2XabRYG3noLQUK1EEqpRE
qkMgxg/Dxk4WuFETkY13u2khRGK+SnnENRxeFEsEODVv62DxW8m+WzspAoT7p1SZ
7Vi9tSVEBVg/odqt/v59bDrP62P7BRcF/R5ao8b65BqBahRg0Ux21KmkjqINSgNy
/0QkInJkloekIvO7DFOqjwmvqoZboZp072qRyT1a+Y0SpLINzBpju9+4dqqKEkzB
w79AjTPnmfxlyeLNgQzkZ1tcwI8aULrcFOVrFxUtcZChTc6xtDmtwH2FlBeOWvsB
GYg5W+SEuXAV2+UN1X03aUAcHjlXr4vahVEnaw3/qo8pg2NOrS40d7slSvAccw5V
mTdMOgGyclz+OD1nlaa1EFjnAmnLPFhaadR5hBosJiWVMCpB/CB2kgCx4uIwJImT
5Zw5Bpc/EB8ZTpIDgISSOkWRiTeVgrjrwZtqp+c0GsUTAFHLMMvRLT5yzZpPUzrx
NZ0pWnTGTCKjmZe702RKt4ih9Emm+HxqkzhxqswAKfJzUPmhiKdBPF1uNwEGB1rM
LdxHG/P1mvRq9xfq9lLONbk5BTgMmg7c4ajXUw781/xRPuoRpItevwvWsaQghIor
EVVbNJz98CrWSqAgESemFPtx6DetzLDV7NiPFyl8ZiS3FH9IXcyiVQIIrE4v+ecf
HCqNGv/D1FTtaC6BfY2iofKIS/VgnsTqtF1RVeJQU5GFoBZ5vmZEslcXbAgReTbx
bk/2hbfgLP3g7oxccQlBhh7iNDDugQTyR+mPzCTmihEWA3jezkAULCAuGIlUUXjy
NgAKjNC7BR479KB1Q4IMwKXH+KF/Aq+JOn0+v01nQwZRkkXCF6StqvlUOG55Yi/0
4qbFovaGWx491hEm3S6t5Wbtavb2mnGkwU98R07oEkOcBgpdm9GHwNjJ6uxIXGAH
ljRvb+eMMgTkFETwKuaHadjmC62MidGYtuc1cybj8evOH819NsKTk7Ktz7eBXpRi
M5L/IlS68a4Oe2cj6sMORiTbEqfRMWIoEO25ckQMOphZLGTVd7tJFKiq65cnMRcJ
e4DGBFan6S+pviR81pxZudS0Gu5xA042DmVsipgE/ZwA7TeaJV6PtdpCSw+MVrQc
zJ7eOkIAovoD1QDMDldmC5QprtXv8XuwJFMIHmXJrAdNbwcd46La2AsYtt0xG0BD
5m0rb7t012HEMk0OM+I6mB2LPEOUwYa5VpZIwkfBXA3odAUfJ5FWCzKLKpbm+1wC
5NfKb7179BVc7RgMPePznILzKMozbgs0a42dk1sPuOSCpfAHtG3YWlJFKyqGp+5V
GOFZVWHvoVC1fR6KeKnh/OFIqI/FVzAwjwwyBq73Ipl9iecdVpNx/i/mAod9YG8m
8jcCf5eT6dZVXz8uc4028IfWdvw4rZxo0eT+jmen5+761OHGcD5MRWOqdS0a6oEE
tNMMdN+5GuqmSTpwjWvA1wtXJrL64UUstUXCR5znwMjrw4SC172VUmDLMpeeQn2W
2tVMiXSUutA3qfleNU2kxQOxlJlXKWLMeGA8vXHH2ZJClZWOWBOv7CKYeg1TQws3
vsZfUQZjuXuPWsJeP43ThMbAaUuSMpKEGlFpzXBM8VWuMVi2/B8d71agpw9h9lC9
fXdLVjpA09om0RoI8R0fqwKxmsi6rbJm//g3xcSn+JifHiAvvmgB6PzHaskvZfyW
dnEmNp47sEZYx8+NOb8bOhl4kpdd44EGEvc9cfNHI7R6SMSMFPQ4WrLw8cIqvQTg
8J9vF0dAA/44rOKPO7KVgWmDcHyqjFCmMmEdmrGMScuBCwOHcB5rzZ25y+2zIP3A
LoG9jSEFg+Z+h/p1IDIvBkGyTheHx7wBMEFcsBhAotZhuOQiqmEg5Y82uQXozGo3
6M3dzH+diYv3W2C6UpsrOxVkodcTPqUqIzNdb4J6Y68syOFPqt7JX4QBTvrfqs7q
xtlOaO6O/+YIdqJJqhzBHRUkv7TaJojwFPyrbiEWK5wEFCf/zwX3qh44/D/Ab2SG
yajGu8TaaMZPt0edmF75prUES8v8ISFy2ZDMB/tNSxoZ6yKE3ojwiOrkPBaHeXN8
Cy65rWdkDZWpNK9uAjUQleuJiJbLEPfKfO2BGKtK5hMNv4DqN58Y++/lUvbKO3aa
dHuXftf2Mm3EGcKWi8d66n9muUoHThth7JYtMeVmk4wO0hE/DzEOMD3fwBLvKlO0
KKyTGqfDsgMd3nTZvloS+JGs5cBVUdC0VOV/so2o/kQR7RNVDLR1wZtRRoKXBPDF
eZ1ttFct5RQtkJzG7XBTXTNxiffQr4uGikd2/irfG+tdE+9JWbkZFezelg0E9u92
xwBhDt914oxBIKhNuZKpKSYOqwNCrSLPDMegiaogt7e7+XVy6HreUx9mza7PPUdW
Nz6fl5qZC4cO0cR1k9MrDac5TNShKbCO8s7t9jcdEqYPs6XAyRvF7mKYjvPGooaQ
kItF13BNODGEgHGR9Lc6tfSmwt9tYksMmaPiZtRWbaPFofOhYddePFj4w6EaAv30
8ckqArE6OW8Z5IhxhwdjyrqFpJqfJfX+EAFgNBlACUQ2sdhmpGDD4/FxWq9+WeDO
WSBLpNy/EvlAdw7rKngIzZHIX02EUN8aUiBPNAXwiLC2zlbZjCIBrh6N3HJk1bZ5
AB21Fv1calHvzdf+Egtp2Al3zf/6K0FtPUGkx82l4206kvoVLYyaWFdSgl+ouSzV
apG97kdl45kZE/wdhW+Q/yzP7NBSS/ad1dAH/zFOE3+EPhKokUuGD2bYZg173tD7
oLh4U2MCsCOe9M00293upNsYHLETmJXfdkKDipCV0jUsr4j6sIn+ieqVhp0s1yAD
00blwrTUFeDNX5rs7OqdHE4bwgsnm0NKqox86aYtqAjB8XuPBo8vvS4cP7yACHig
omKf8qlqtB238r6dCyPVUMy7QiKrmJjI/VuE4cTKr6mZZQ3gKLu4vB9iAo3EKRy8
wv5BxB8K63klm+Ywl/k3t4AHAcZHMg3JYdDwPnyKmMASFBzUo1QzO476hLEAxn9f
FdSIkkzRr6jNUHLWlYK0Il9UVxJiRTzGFqKe43KOk5/jrbuUMZOECYilgSfAEt9h
howPIUpnD7Rq3dBX+xVlYTnZRR4yFGz68WwKvtI477q3bmqbPjPiGf67J8RQzi1V
EVAGWOM7hs9kZAeH9O6TMefZUjOKAygv1N0sFLbCgBec9WI7LwFTBmQFSX0T9/h6
oxlLBxTEPapREeMhYUl7MbWVUigdFfupEburcwHLc1asZvvm7yYP9BIXNLSwikmF
OwQG3zjjgWqF5+LrJ/Rth0VFqL1rhLufDjZuTfSKvY0Rg/twkuKUhFikc8I5lyCP
1B4oxmeKeeOuTyYYfKLVETJSMPY2uBlc/49BScLI7V5nNpFMqIjAVG2I6uamJOgS
ySEzr2uxUtEJU8Aw/l3xiMG7xs7RzZhgGH068IGIJWudNaCTZOE5iUxzR7I/b33H
KfF8NNZV09/ShtKum2fp0EhGRUKvYqxlBea4uMt+Q8BinrlcO6vzmV/55DanPoa8
F2BZU7QCOSs1551S39E4sa3Ok3fMdNQAnm9RAAkB9kcyF8aDExDgcnMw0ydbsiKJ
xggIxx+0vcqzA8XxEH6tjiIyV/XSJijR+/XNK/X9edKiUsyPhv3UUxC5V+ZrGekR
5fCwgN7WPFlHZVgHOvGEbvG+MSSwcpBw88XD1/uQ25k5shzSAD4KdBp8erodgZ2o
Zsgg7fb6T6BBKZrsdIAJ9TtDnoSNV8BAjEyDlDChOe3ZpJmOLTVdQKv3nBvW/4vw
xD5q8UIPYDjuduixd6Qp56415spDvoqRTNX32W1qNjW/sfO5lWsewR3TKGMNREeT
sDKfsRt1JCxpMUvxQWY4vTLFJLkNnxJ6uDmSl/PHKjdDgKnkFizGL3nTSdxMW6rR
id/Bn9Ty1G9gmS1kXHJ6EybViunSthKUSolK3yBCpkRaOxwo/XWZ3SzldqmWjtcP
tWbK4C1+cB904ymRd/q8ASErxwsTTYgrG+Fr3UfbPlHdWQ5rHhY6yUTc9Efn5jqn
6V3Pc2Nvj0u6cnQoYy4gFP5i+JJdogGQNHfHwxaEG3dM4T7yO8kalPrHIj1g4+6R
HWzvNEdWHDSszAqdZtRQ71Rq7OaD4N+8bxS5skD0075zbjKXzBdlxU7Nn2pScgoG
qaPOrbHNn+3JL4A32vIHwT4kj4aO3B9KxNi5Zj2BEkjRdzqwZPgjraY3/T7ny4tb
LwRYNWwftpqUaXp0lN5X2Oqb7qPRzGPOLX/JjjIG85np7h3et/R8u8I6QGmTaSct
N3bt9f0Ete9Yv1V65oF7ACqMxqJ/CYkv4Rslc+YUGYl40zWXSVf3kEpHueTqcKrA
Q3cgzO0dT2lO03gsf9sjjLT5e/yQitwcszDlucifCigxxZxcAzVhcpainlf0+mHL
DuQAJK4emistxKSCEVKjjHeh3ApLAQRYEpagZ7diWyZNjlDzSHwpsu37PMgySsdQ
SHl2xiPL2mmZRvczemONG/S00zAKz0FBaZKJvyhDViOJaZ+W5pI64be67XrZiQIW
5rXMomvfDSgo6DMmA/sm3DkI3CVivMVsYSE4IJOBrxDSzEcc3lM/HsBppZVe/1Sd
8H2RhTpM4/GWn7par849QTPRxoekqIilWxYpBvcziQTXPY3OzSifUshUeI3pmyGR
Xn5dhdEne5ABfARSeeNHSC+Es2Wyni1hzMeNMX77j6SgunUgtdRBUAu+quF5nIo1
Y/EsVUKkcsfufnWk9kqDBUuD5zTtzfeUdDBWusrzmpxEw6XdJ2ALZTSXnJYym+dO
tLOG3OwoSLmg3GZRoDyEsoc5R2EnJLXIXSM5NkaQMgYoyACVb8esKXd+8mRA9jDW
yo+6azf+E3WS3m+faCitESnhxjZc56bnLgJDVc3IIwQzNUrgzjMyyJVoXgO4lZI0
3KHfeQGSxb934c+FtZVM+r5cGWGQ9w1AMoztDxSoGEKu3J91bY5oMbHTpch1a30J
I46LjcYaQQ6ChfRLajJhwaCI77bgNMeCvkWMmQiOhvg3yY47NCQEhFmpkAE+htpk
UBpeCbPVM3hWva7EildcwHqC9LTLpNX6pCNmmiFQn9cwdgbju9kpXJRS4dfCI29s
vowKkHf5nmrLlR2U2hfKt4w/wjy26Bv/6iRDddlb/ri0hNX4kERjrS7zzN5ji3TW
1fv1yTkNxA8V8Ap3uclx3gAYTazoXpTfHIdCRQXZwDjc3iHC1wdohLCh5s8h5TOs
Gazgw+bPilTZSEsyDnKye852YmtvyEGlFCemF90qQy5womFHpmx7xOzIn81Dw70a
3e7hR5Axr28DviWMYhLMRcdqWi/+J9IH/KgNjjvgbfxMzPyhsaEns8d6oWGlqZUc
tF5pbvqxi9Oza3cn+6tHa4BF+3Za5+G6kvzL1+rjeez6A/5vQFqJu6rICMLqOob7
efpQdLIrC9NO65uEViznfBt+8tr4yNdn1To7wQnIIJtnMqYFGE3HIvIo+Rget9Qn
vhldPqCM4j4BuV3c9bEzdsq5FjI5zLSxgVLbcSlnN2CHTFP7GaWZ3EYYottLKKnY
HZ2pACnuOLlQ4C9pMQfwcACreeR9OUoxd/15HaXxEoc/IZ30y5KMEBOXVw0QvsEn
sQcX+3izQs4EQm/aMdy2uzEiDJKHC4SdBcdvVMAYzthpDUB3AddLwHJ5sn5FYdnE
8zzZVGNyC/HEhgnR9Kpgn/HXab9sBt7Xr4RXXvSCAMeoX9eXavkk3s+ht19rr25v
uuS0poZEpjESWkXJya7wDmeb8C1mG9r6/gSolZTKiGjHolo8/r1bXYQus4ve5hoF
pR/pfuzfX51//O2Asr2OkIfsZcb8Vlpy8GAy9M9Su8TRzWvjMq/R5OKe3n1FeDBe
8UTFsP2ikgB955jmFm9PwjxyRuCIgV5gmC5OKb1/QKN5Um/m7C6+JVetRGjwpWUD
mnSC4hsZmUkElARy+E1XYBaKn9LV3RLCgE2wr/Gli8jt+GxMXjaHPfJc7FQ0uAv8
vPzOaHH/SuwEgtN8iaSJt6qxv3ZyTy2k48RoiFz2R/wHZAagpPyDzxj0De+QBr2h
MFidHknMP1pylhz+s+K5+P4f19mB1fzWdbFj/+GCpjLYpGBU2epS6CdqzewA5LN1
XqIK82dinUAimf/6Fh72X1SH555Jv8bTq1fo+LOxTmPUIFIgfvsbfH3PAslUHTzo
1v30hCf92wfByXGjLhiUFd8bUtXjbz8EleR6YnhHZYRiGBtr3Cv2yhOSTL6F6sYK
ghqXnuJ4azEnp5Pbtu46TL+edjG6BEMxgII7UKaccC9jBwN/Q5qTPpdCwMQtAovf
ELbMptBw00JgQGeQCmKfzOLAK8s4z//pSIFc28khl+nT2M5fKMhQ3eFsPyvkdEwb
FCEVc1EdfgzwkdBHxLQLTsfgycoaEElRmn2BcoQoJ19WfKSsJFmpeIu5X9iUp7Yl
YtRvko6+Bp1qatJl5wlxUIU3dm1S4bDNO+cplgp9gqbyOeTYmEFxhXbtmkvAJ64z
Owu5yTMiaBqOtzSAkF1Pahrtz393Ltke8ca0vAjmStD4UXA9SHUvKnmtEUTvqLIN
DK1oppRt/AkaMKWDQ6gK/hVwCsd2cAgQDq3AShFgOBiAbrtmh1Y5iHGtETOvfeSx
+mU4alOEhh3vzGDhTrJ+olUos4Lo0WJGsIjNJ7He5Vzi2yaXmWMpKb7moSYRezGY
jI75GqRtoRzqh//UjVRLhQDMHEoPm3c1/6QRR1VtG8Lc0PHCPyKRImliYyjjB4yZ
0JxxSYjT1GI+OBBde+lUJJizuObGFjjLv//t47cr/RhitNVg7xiCZ12qYjlxzlbG
hlCSgr0PRFxr5P5tRhB8kOUtqvtZGa8gtyMBZ0ZgidW42h9PI6OlNJuohqKm1A4F
Nzq2EAUTAOAdCLyinboJ7DLtEmqghnL5+rsRNESRoa2gYuA+qLHB/4zgHL1FSegl
yGBBC3itnwcocezkGhTfytfx9rMvwcWz4woRpkJMXjn/p0bCsTPxGDDGsWbX6ODu
TYNZjClxzczbNHBIitmGDHiH/kMjr7mwVZQYYdz7wsH0XHe3ISpk9NplR0FnQm5W
cbAqpE2xqaFsFttS6saCNbVxMMWchxYD9yai66uJlf2rmcD5MZLfMiYU8wkKG9LW
dTXw13ESGHr2PFIrKeZIyWSitWtIm6Gwpu7HeRdIifDdDRF5Q3jQ4WsP4Lt6duS2
JOo4s87rNYEIaLyZUP5qxZ6FxzcJ0Gh3PKC1HGAjbhbRsWV1fp++rfbORF1Jy/KL
3RQhSjmNFsK8j4Sv/PDltru9LPuqqh3Dfg7gdLQ86uGaXqTYukc7Zs7OApPbvzY8
hrw8SSxj8blGbtLWXZ6UKB4N4kMdVyZMqRt5Q4iMzHAXVWkpxWtyjqhbgRAtbx+I
2jKncTeOHOzQyrHhKmiB8kuph6q12XI+ggaYCdzGLA4IRM1BbItXquv4PH1H7VBJ
yoYJHS5UnZ8RCcaWqoxt9dpDv3q/WME9vN4C38rPy/oi+dSPzXC4+9/BWw3tFfgT
Y01qSHx0uPRB0ywDbrTb2VGXRQdsifvp2M3k4x6v9yaj/sVIgtSNCkbhojJQJP7d
2lKto4pJzw08Tqe1D7moWZ1GHF5/hl5RMq4/kZTKlLtrW78w/FC2jEpT2O9vKTwg
8vETL3F2jKrQ0g5AjpJe3OQzpr3zkHgLwon8ad0JmNeG1voPw08teGRt8w8WO43B
u0bSvX94DfHAM8fGgXTJbMmkPvL4rywO3fKuS8mDJ401svZiWRt8GS7wdxKvmFKq
80I6ihP2SZE4Am4hXrJJkJU2yy8i78jhCpj89n/+Pi4hptE1SVZxFSaoPTKaT0T7
NV8qVBJZRUUSZd7/+YR0MOnkJNOcCYX9PEx3VvTvVbbN70s+FlPwDM3oEEBUMT8E
JWCGuzIbNe9AbjI8pkaUS+q2vF5slbipD0rfjj42zy0N0LI9zkkxxz+MRyqwoVhx
lYS0whJyibF4duRjwFYbx4ALtPcKnF0HnDYcvEioPW38uXKxF1uPGrBKO9UMQ598
VCKndlPjl2oYjTOTKC3BChcQaoD3x53kOiPdibWe6yczW3SmF8iR/iix9N7ws74q
Jcj8b6//nvO4H5qFMqDnsGWf5VsBRqFDpuc88ijwztwP2BidWraKNsDRnnIKmBeX
DxQxS+puZX4Apzyeg7eke16fc3WIK94j+YYfejGE41Z5z16FnP2dYRf5s2DyLTk/
97fKNhjnmnSCeYK1eLHdBPdcmeO7vDLvONXMNx9LwiS4eBaRRAAsYDk7hFcxz8p9
0lNTDjnQc6Qa8jBC3WIqSdtNUN8MARxHkCGG3xgqamqgioaKArPa/kfJxgMnxlOt
lKsGNAjafm6oXOccvkHNoEbpAukRRXVDEOLPaCEOBjrwqk3w1ogpJ9SnZ+LRPuV3
hKtTOoiHgo8YfAeqipVD6L17IJRf1YsS99x5FsB2Ik5KH274vWIJAyRpGncwLXWc
BzLYXFQ3M5BSEvgNXSUf9oVy1md+xmnUdV+rBNy3vqTYYd2rZFiMpMOgutzueZAl
oTZlTpdAnHt4Lx22/2Niq9Ct72v/U/mUxA11CEp8uUWUJJ8VXXUzozlO/ly7aEnT
egxTkZgU6B+7liszoiwI5HrCLDiWR1/qohaWM71J2y+vRvsHWWPhc1HsNyx7JXqo
76u5ZkCvFbLU9sGAoGGL3R9yZv/tuF8LW95ncEwWpedadyFb8fgF6kjlRIRsprDR
VzPschfv2fqr5HDpQ6psCAN605dIZAMFlPUWs896sLYziWpKfwekeyfRz7hoOtmK
jY7zA7lcAW05HGolF6rKOdhxXFi6PZKVVzeTXFd30d8QAqkTleUVRCff+xLVqtTN
A0ql331g4m6YYg0G+ftqKzR4YVufYHSq20vl1mH7ObfqBIHz7dj1WdxsXvkUvikD
RgWt/2BIN3S7Pt9iQ0rX4EAPu84/q9UM6eA+T6AFJvsc2HLfbIPsb+0k4fSJuSw+
tUKKyjd3fVzxBX6lp5NpLghovkBfD2mR/to+nIk5AaTPtHnzJA/NWlGx0h/HNTWZ
MRoxXu3MT8prUj3uNRbxPXVLUtW9FRe7QjQlq/LGK28ARRGJX+Eg/PCklw+xudpI
OnP4PSoA8VFWJfRGrn2E+XjfNQH1PPEhfq2RHZmoS804VObvz92+ppwdaj/Ed0Ee
XNjXHrLDkDmEwU5KkBF0c1w8oX0MuG8DJ6zpaXg8KSBiacf1gFfsYIaMWQ+5QFqT
m1RDoNmfA2SjZCAk+OILqzXh1Uwblr4O5ihTM6GoiKKrvO+0Vta9sha1BvbN89Fh
nuF2MMjMUrF4y9aibd9yMuCqdRprNXa96ghqIj/VQ/hpGJJNUshx9fXLJMN0i48a
R7B7/GXZz1TFwOYUjuEARozGjgzs9iuE6wVMejSLl7aRYgesWNxpf8uJN7f8jkWU
jXDMjUAr5WbuD5NoEeDhCa0xNW41YYCKue3LNppGKJIHqENu0+NYb8jAH0R9IsPf
YrQZXUmT9UOW/t+0ZLsf/c0+dXZXCISfCNHwJr1E98iwsYz4BLwJKbab+V6+G2jL
HP14svOxx65YD9oAJMMX6A5XXmvrOGaZbkcVNqbZFYRNAeaZ/sZeRunF7RyQzjjh
8n6Tzh1KLcUurDsk2h5mDzbIdRtV7ntZZSzIg3kPHCTPARz/9wvW/zTd92oYD+xY
JuOiyGEPz/mZoOQFe4XL1pB1L9Ybi/73CLiXirkiMwIuQLbyV3TYYmFw6yHm0+9Q
tC0VKR8eV5mIC2BBN4fqC/0c7kBDEBEiqQ2NjgfJP1T2Wl27WPcmFzGDKZmVUJBj
RAufcYrdfOM2Q9eRcngrEXfo6mmRbvgEZNS+ydsY+ZEAXPMVTbcl9fyJCYUvxlIx
LXrsIpL5zJkD1GgiRciq8u7EpgFg6ggDPOH02w3gF86jnmvQZ6j1lCXTDU9oBOIy
IdywoNZSzVE8/L2poK6emrAQFW6OTjGgsGIbCN4oZuup0UHlDl+rWmeTlzxZugxj
kyxGB5vcbyr//ngewjEZWGzmldhu/6UUm5p7BCALEUWqNIHwvZw7n5xANQCEpiAb
54x/nvGPtq62oKs8WttGr37NbqPKbosTr5ik4LVufEBcMEjYfePhzqV0/P+oCi8t
`pragma protect end_protected
