`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kjys85yABO/KwdL0XdWjmdGd9hGzuJkyo7Xoyd+E0JcVIOMR/yc6La6GSZ/YmIy3
ehqKuS8uQfrxZBRRKPzeuNYpvCDfiyE73D/CM3rxIzqnjVPLJCVJipnt0HZDGIY7
MzhEcNT0BQSoTvdvgBRV6N1NtW/VYFcDFavhyaX7g2s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8144)
uCHvkBE+S52CJB4su7JMgHR44wi5d3lSqwwhiHs3B/ySfue+8tV3T0382g6Dyu5K
/mM/k8BDyiRKl6nh0XPnjhOhgZAe05ZVD+1ASt48ezlUB8269TsIAEMGy0UZAX1y
a1BfyHWharw84TOIVnSMa0Lqvw5G5IaMeeB7r93TZIV3VIGkAjcnImrWWTVVlpNG
fOmT80HBzgBR9iqdR5Kl6PveQblsoIcc2vgmZ6ZPJDXgZyx/BPcdVQfYvtuP4ZiN
pxc/86AjJxumFKrzi5WIAW9AcZ2sv7TjkU+sqhmhQdJSjziklh591HlZtf6KaKEZ
fmbDjG0poLLqdo+Z0lsua/Ugf/FKvZUfYZ+t8kG28pKoqEbhDxA4kyMmrwnY+QOx
n3NLEQbeyfjMeUYOFYkFpxpFjjaM/fWoXqJgw32GNLYIyTKDFdvuTwsah4EcykzU
l+odrrfwNF5b+OI9uZoPJxpsJxWxz1+G044wqUMmUNXKpUe3StyfY1KRhycIAM+a
w1DtaZGLlX+E1/lhVJRrljPDkMpuKRtXsZMS9574IfORkqubO30Y8FUOG5t0cDxQ
VDAAehr+wwbJniW86B9i788DN6D329O1uqoZujNwEQSzY7JXTVKsSeE0//5AdciU
jleEqaVK66NI1PfRIwZeFvrjllt84yrM/Gx610QGovdkKr2x1zdVURV40todkJGH
eXkXM4jJa/pSjuKFc1ybtuEo6fQ/vwwkqdh0Nqf23hUiibzmyEbNN8wh9PwqOkBQ
dha+uCbeOiTp89hTSEFF2/z6JZoY0o8eoBw4i3y4Yt0OJ20neZyXtvSyp6U25V7K
XzbQR/yEz02gva4Fmlx/u1RQaeATDYBxI+B/TTicFsurFOJktQMiv2wzEZIpeBSF
0ABo8gpuW1fpJ0h3TIryRB042fi3H+Lp5PdCzW00z8+AUuXBf20a5pjqI3OervTF
zjYHEe04aZN3HbURkuTD8DbXVx5xXVa/7712cQIbZZsRJwKN2kBGRn/uugzTN1ix
mL8O1YfGcc39WkQ60LKnB9LM16uYrmQk502zRhSzkN1D6v4EJqIkRvYzHyiwDRf+
7HK6leEjmvlqXPaUEePC/iHOncwNqdytEvMneqxK9eR5G3mxqgZQAnaS3ZiqvIao
thy1KI6dBRaoDu4T09gxuMGQC6sSTRkaMEGJgwffceIu9lbT6wr2qn+CJjIoagSK
27ciY8j/5R+PaF73tCq3hLRVj6Js4f9a3+GX+gW8U7ehkMmS1gIQWcNCkCisSh+A
FsZUmgcMv+s2oCkEtuIXUTv6d4yDPj37Yq+7u8bYQjolf0Zq0W5mpPDQhhzYiJb0
NF99MdU23URqJGhW7/Ozvkko7IfjaJHHuVoG9NYX1zv/qPlacvA3NdBjkcVFDW5e
ltQK2BasO4Y+Qh02FNcFQXYevafC69i5TvGZccjlIj63HnSd+K9i36bFN+zYR9UR
renM3xobIpxexLbTKqqZ6N6N6fERywC3tWDsaVH0iVl40a2Ctv2BINcMhuQKGI6A
W0OmGlqpiRxTs17RL+W3q0RlE1xcO37ySgzNfFh8usai0MkSfml0fn9MSCqokRdv
YEgbjJhyusGcMINpXQIk1KTQxKKmMphku48HSk4cn1/845SIgd5JdgaFpF+4oq6k
moeMwp2mhHflAbU2GK6JjySasSHuhazJbF2seBuLGRxdL1GZrP3TMP/0Q1i/7PlJ
s+adXcAaJ+gXzEQctfsuxOL+GWiG36jKUJk0E/dfDGE2Oy+Jv3ypD9w7u95CO0I7
TRdl24pwWjluHBaB8RWFr6dDv/nZheGcwqfI1ZzUvK24TCdkS3OyhhbAJCjnkx5M
GyXNMK8ljLDFeDx8uwX8pDBFEbxZXXsAxSstezypZgcK2w0Ycuu91ErNfCFKlcfS
eLxCSzaqwCkBWw3KOWWpQmO7MOjhWmm/ljGy4NJyOb7Vcwsj9y9uhgpZLPbiKmbI
18f3pwMRAnboh1SCqPQdMLFLvb99Ml446qOt+QVHD+3oryWfW0+IJxohfH6ZT3E0
RPEPUQBFpTSvGfgllrmuKnuCd1wz7em/V6auPfFeaSlJatqRJAunLxNw/rar+zCU
/UjGO5E3K5Z5Uq0eZBeGM+Re03G9EGpwqHi9mqdKFJLLIhMAdOBgGGivvd5v4jGH
tHF5I7vHpHhJmy5ed3BUgbdbdkvqtRC09am35ZAb5PP/NmsHa3DtZGv/oyi5+2qA
qXcrSOP3chlX2u1BXXrxOsDRgeQOAiUh5tvSOekUyXshFgMTRmKLuktqQmIoexZN
LcxAZESEgvc2g8/ZWvg5rjO8+K4fFPfNC6LBBGJWM2gMD4SeCab5MiNwEMalx0SY
JufhQUnT99mRc7Ezf/7gvLi0iGkDzIX47smurnz2OLKoBTTrh+zg81uYEoEARZIL
3zw19B0qbqzpuvO7aTtcIDpni/cP5eyj0y/Gt47sSlnqQ2frZLiYqnQdp73er86o
v3xJo9LsJ2e3/TBwsH8KMiZlrlk8KSa8ifJNOuGJTYHYHkt2B8/gQR/rpQReY7jB
uhqMwnWP3aP8jAnF5Zs6psT/xN/p9olI79j74ZdqE6iJofEer6qCK1vmPCcy8RRW
tVTYaQyhOaA23TVc/nhJhcwpSibk6xGc2n66a9AJ0sC2FwL/k31LANsSUsbJcyfO
Nymn4cXaoshgCorHecC7bL4wr7KiOj7fingsAbIBsnYDWaX4ZZPjl5FE1uigrx5S
kC8SimPEv5SJ4rgZFXkVQUVIt1xfp8dv1OyXC9tVy/IfAd/mY7cilUiqjfgXpE52
UFOfgvo2E5r79+4vmrRFBI+sPfSq8NoaXQxslm/sXAxKCe8cEVYz/PakpIkYU/ba
r6kmhg6es5xbttpDWDmk06wmfxAYGBx7aDXTwSDbl0IrMUt2+Zd6C+3/D1ZaE23o
KgX5G5F465KSlBpz33qJpZATf9S0KagMHhOnjUyd/Jo8l/bU+duX/wGvp+xn8V8w
7iTZHrrn4AeW68FmbWItQ3ykJCEIpvX+DRKWQX5P8JI8ztV2lCREeZs9LXgfK/mx
keuWqHnJqVOivu4AjMUrRbGG63QPjwHr7ogLBzlZiaY/DeCAF5JD8EXp2hZjwbFf
0H/cTZFAQUiE8zLbx1ARV7sDSgJh6duLBuiGts3M2vvi2GyQfvLMutqQxLOMSKEZ
nZc6R+IsDM6vFb+VntxmOqvNOKE/psWiupWZ/1ZJN+drFugua6LSMD6iPYkmU95d
fNuNfs5GdwiiLVHeMf7UE1A5rqK4VSwKuMnSW61BBC++EHYOWKiJIktid/TEPyA6
dVHM3k4TKQQEORKxkA/qwayaBuZmzXKEJ0mWbF85Vm58M2aKHWXO7H8EBRdllvfp
BG28VeyfsOLhsIEVhivPWnk6LPNRyaBwitN9lP3tT+DIZObGxblaDaCQuvwNAEAc
diy/DMnf7jnLbnMzIY5+/JTmML5OggfNNmwdRCHO79XD7GGddhMZFl5T3OKPHa4Y
sav3hqaCqXyUaywpRyZS34CKx/7tBGTaoY/vGfOCuLZAEAWb/wc4uUE+1lOlP5AM
sSCsjy0wuekCSXqXtl7dnR1j5E9hQZSMQm6CrdfAxJgyAFqIi5l8yi/Tkf7lchfN
vyMSvLvXUTLj02hfzMxgSvgHXXVUCAW4wDvULMyX4JtjTXcO30B14npDS6DVTIn+
E/BLdCMQ8ENyCUuqCfzP365kCHNcuvIBCCMs/zUP/d1/0exn86gGtXUCv/C5y3B5
jVn2ecb6gZNzBc+7+PElX6mz1JygOmkN+ewGah/ek+PvGpBsvUGrvIDCKdM2stGE
P5e4DvRnL/A4rPj1RrpcEqikCa2dUcA8pCnoR3q6F90g6icUSWPw2VxUqxFeuVfW
tt3O1r92ZogDGqviGRSRgRgPvgEWAZi9LKRh0wh3fQAUy2ocUVM8nDnJSsuRmax+
tM4SSBhvKhddl2fVdvNI591iGliDgHZRWyOQwIPuvc0SwVK8NmBKEif92eyfz17N
qGzNghzjs/+2cXkum8MPxyxErRAsRtyugtJyxiFRRC98/WeszGaOfVGzm9ZnwvYc
xGppT5ZDod9k7Fy9GHYaNuUYJZsK/bLMzM7eOTxLyvEpnvHavMic4QiKYT03OTwX
zi75t13Tvl7sKwFqAUe//MzOdNECoCcY7y7IVNAA/QpwP7xJMb0flYTDDFL7qmUW
x036Abxtwp7njJZi+6PBE13d59OCWSuBTFCQrAQeJnj8jImELUa8evV8hDO35WNj
Iaasv6l8UWJzrYoZnOXtEE4z+cLYhX2fb8kRjrGgI8S47lX7I7/olWbphQAC0IaU
vepywvGGT4jTFbU1F0l9YwMl6xevrLhnzX/jEVeLhY7CPaZdTCYs4rHMveZGvo/N
52ycsAtnPHN5fx9s9df1/HooGhkcuRd8N1AvsWRg1Cx9bJraPrzN0PWCKgX8TAHw
b8VWSayr5YYGliK2lWDl1PRkwDSCCeKv5DMfWuwui4rh1dFhsCoK/TQYIFuKdzI+
PiTJopT78KIrumLsahuJq3tXyff55/nN0DMkjxhh/uESxRKhDFvJRTtpSrXVg0zb
acsDksow8A3L5UI6qfekbVYvbUE/yb+kYFD00j1b7OLCLqVEOLTcJz9/ZifrggEN
9F/kPHmUdJZrpSsma4HOBniiLQpvu5XkNXMBIMjDWThpP36g4J8FaskGiljaRtay
vem2H2dN/K4u8EffePB1QrLsPcZZDNeacF0VxdYSUkr3lAofmN8CSS5ZHZEWTiPN
KJc3EsSE5UcJ05jpTL/444VTgrlUq22hQ+vUXtKs/Kpl5L5lDIYxjIjSzYAgIzsU
RKs+8oeAl4P+YDCZJzoNcJklSJ+rqxE0+yWIhSMOiX6DPXZhe7j251AnawCsVbDI
sLSS+hg36s5CtE95v+YuQjbGwq/eXluUlgzCCk8i7eGEHyrfe59AbQBVwDvHwFrw
BjyhzbNWTfp56HUx4kGtufemZ0L1UXO0AAnJY6f78MWANqM3n0vNScc5DB2aVl96
BzMqzhB2trsJ6hHD4cF0y/fMNx0oJE4Q2QIrmwdy0yhYoyHUDwcMSMsSZ6ix/KOh
NU7JnzpbBXYur2alqrdpv7Pdp/8ITTYvLkZFZJ8bhymQsmHZPp3LDbvlWd6KYJOw
4dqCTcEZvEeggd1n7fyF855Sd63yMtMBGMEAZPJ81cjyj0IRC3jJYkRAiHq3kREW
QnNJaKFyywVcccSfLBSj6d8F3RqhnqvrnWkvNWe/jKR34aoCaf1IkXo5Qpi0Xboh
i+luADm1NR065hZ8uPC52Az5nU84bcQ/mHR9akkfnkx6PmqKouseIZ1Ptv4tKoZH
knMP/iTy0KwOPMUZxiDnyvRMhSOtt1JKT0LvhRF0UaTqIAfPiC99/7qIEDCvqwWl
IDKjlMA2i2oKkH6Wd6fOwNofaT0ItGGFUaDT8av2cXcgFWU5qSVGH+XPp3XbM4L8
PnkL9YTXff7sot/m97AeP6Aaj/vmiCnvdVwEyEiq95Ff1pkwdHw8H90D9eEGkAEC
ZvsArBgh5xoOg9F2qvpH2OuGGraTxfMh2Ly5ForpYvUqaDfJrxW5Z1EPN4b8boWd
MqtVbu4G5cNuwM9n9x5/EQGk2TWw/zUSwfqH5fet6EMC+zWMsMv8+REohCuV5rjH
BswZD3VVSzieOVau4dkRrga/jRb4u6+Gl2HflFNbNa56706mpBhozq7cEqFYHCkR
YOWi31b3GFajeekgn1hN5gAyO+IfJOsFu83it1XXx7tybTXLsUqRw/oaiye2KGCD
Z1fmYC5U46GOxCPkVGM7BeEI/w6sYX1RoUoQqAS4hnCcOVNRPpe1X/6iYDoOT5HX
qB1Jo4+HwhiWxMs0b7y5CYRPEEsLD7DlH0ttkuiLTogCe68tyHIydw+Rrcf9m2i+
ljzr9zo6FaPBLVZyDVklgDeHVrWyhclqVbbMB/Pge7U+veJu6jWtjr/JghvvcLZk
dhWn1jvDSVkbAVh9YDtUtT4kz6mlCrBYI2tNdb++HJCKZyElK/x3SCY9VkFPUBs2
gJm8zkw2j4ercpxHfzdiDSSqUmyTFmERD/M5QY7JCT5q13n/BLc33kJe3SyXUai6
oC2d9IBIH/ubVE+gLCB+cQ8HCaLFx8ZJTVILcA88Lhe/NdiX/V6du9Vn+mXnzrQS
UkSFZ9V6NFu+vaQh3ydkFUSy2D05Wu6J3Oz5HdQpBpzB1oPHTnX1UcBN+tRm1tml
ZofqU9DOX/lrOAKVZEpMm/gGPbVfLsXjt4uYFvPlgVUX1LXDQGmYtdklHPdCMIjN
MaCwVlrLV0Se3Mws+7E//It8b6mFDFfLNsrBQzQ5zkIjchn+uJ0B2etHBTFYyg15
rqXGcu8MQcdDI7EC3hdAP86+BGIuJHN4a5NzqUdCzBs7DHf4OCmzmYxrLb3muzvh
XVgBCEFKjAb9QxwzudNGs1FpFh2p3stmdddaEY3nuFIL5EK0IFhJuVgkg3LG7bBu
J+0e258garCr3DW4BDWaVudYlgBYe1cK9PhgXvGZk3HV1YfXo2/z83KGPgg2mDAW
i98y77Wt5oZ6PkdSynSB+k9LsE7i/OSr129+TOuZxkYPgAYqjQq/of37lXdSpbPw
YpHWxSTpcnZe3rN3lUDZm688y8LyaXu6gy1HMKS33p5rrkVsv0+q2ixuKkVkQUWZ
TvJt4JOdg/IafXsSOfpQJv19i9bEnMG2mfkJUC9NXeWpmR+CX1ZRHolGv22QmhCU
lH7X7h3eNwAWQ1BgMbCj9Tt1TLF+FCjzH9zl0/PK1kP4Ol5/T1rDYYSJhipTWYCj
rddBRSR3lE0+Yp4NP0iZWv5sjz2ikkFhPWm573Z2AG6oOpyBFtt/0r89xMjrk5SC
9cn/5FMGzVsLc7+KWU9dPYCwj/XDlEdnpLnrnJCq2j3/FMen85xfwOoAw96QhTbF
Oo1/NHCknyvcVOzpgPeM2dLj8Kcho1k+8IEwSsxuYRFiIEgqftyauzj4570kqHJ4
9h7rkMXmssVCedqnMbmqO5JAakUC8oRnl41mTLsJrwYjF9xvq8d3LH5+AzUmhKRZ
klO4FV8Ona9YX8oRTVukM4yegVwcJlqUAN8PGde0iaBp6I4hDxMm+MKKnOKk7Bj2
M/vooyxqoZUpWjMzrzSRYUVydoS0rJ6ymm/Um6orULYIjDw4CDtfxl6b05Otk7nn
OpIpZEMdGnzZfa18IgXhSEeW3AQQv0WFU5gfMEs/LyH870xA6IdH0j2Af9Bv6dyH
bYwic3gx9gyqGrXkuAKL28vJG3XP+X0oc2rExpf/9Ac8hS4uauSmITJKRHMHP5XU
k2WbkHshjWLXI5533XXRS70Qu2oqUs4vFV3Fpe7UCSRebJyvj8rmPHNbRqHbSH+F
b83i6z4nL+D2+eKx8GESL+zo45LoxnbD45w4ai3ff8vpJovYGeq52qn+55BfpAUr
xx7t7ZXtpqDy3uHxDpXyXIOknFxgGc7lhHqC6xPY0Cp/iXpY3tpNikWQPQv+1tDS
CVh4HRaPoGGs3Xaclz+mEaRsiQhLZyl+25aT/IHfiQgWPoOBM0c4oZFV5uWcGoEj
Ze/j2kJUFsQL/YqUkTCjPBY3UYq6e+Qwn9C9gq0JXAua7FLJFJL4qDRq/7h31HSN
C+fISdydCloATrVpIdUMhi+LV3/fJMTfIwTXAE0t2JZEQjEKRC/MEnudUQaVQB4x
GiWB98qMHVaetGi40b2tBeDnyQDJ0otDuHZjGAVbTgFoeKBTwRlSq3F8NaxIkxS6
l9VfRjwHE+CRh7qRzX7u/D5dOsjf1pH9T48gW3SZw+DxR4zCvFrKTGmyYvKRQEXQ
vkVFf6IHHqEi/RqvrrlP2aBt0ZnVPjRKXRG66P7VeVpVRMp9re8hdBYrP9sVdMIW
E2CQgR+u8rgzFEh+eIjXTTWSNCpLZLumOej78x4NJ9PvwCTq9MUk5wrklOPEjf6V
vrtVGHafcAzJh+tfRzCbynFS5f362K3uICW1JZuZEEfq9221M/RvZ6vyWgCv+0f+
DLvCb6ERcHytkV5p73mkUdL9D/DrNfURroaaNuMdeWr0gB16FhgNlaJpLES/olwo
ACYEgo1cp3h1DZXE+tMYAHLG4Ns/6eFgr3gi+/mZHwgGFMX1jm/fq5bay26GbchX
nlGvm7y/Mw2U8gdxFGMAXl+oQPKWDzOQ5sGqjI/HwZqBqUpBlStu5uB8YtjhTGUX
qzcXlKkQSwOf789TXsg7L31v4BAkM+WOho7Ds5xbFaBeF5huurKMFPEu3/yNP8MY
L+YKCSxpnJ/Ly54q3N1HoKViOjN/rHrgbIk+H6OiIMtp6uP4BfKZMIi8gHBryTs8
CQL3Icpij3TDPnvw5B2Z/dC6qX40WHQ7wqnSE8HcNKM/4YK6PuLCDzNuqMF5EqxK
nGlzdWsUVuhEKzX2sGgnzsLiQevG0PIJJhImNkjoWxdfMJLLmkzJbNvvNUZT1d2o
wyP4mDfcaBOoY7HZQA44UYTeoEycvXSP5N8XcGbrjaA9WPpq+HPOuSw/yF1Pw0Va
VkvSPVKxxYkpA4zJ10toIfHrDdCLQBjojq4oNz8mdzISlst6ADgna0m8EicQTB2y
KcFDw4x3+CK7OED7u7zIqSxpe2M4Hn/XgccpFJQ/wqYa33VTh/tNeFMQkbegUv6m
kF7+SyC44yPg6Phum98OGhdCbv09eGezbSNQf1GNUc4DIC06Ft4xRgGUwcujcuw1
dh+lC24lHVqynogfambO3VKV0LWJx5+N4NRg8TgFna3lX2hI5Z2t2/z5ju8EenfW
oKuRYLBK3VDyo73Bir8nCOnOfXLH/IpzX3UFNvC3iEvQyuewzJSIRI5+WEIZveBC
R4cGMQlLZSmbZhnXqklKtTScEGZSiEf+fkP07XYgWOGWCqEXc/Uzn5vZwFFScKYN
EU81wzTm7oNoXUVMv2xT08hFf+9rthc78aN5UvoDXKwMKCSUcP1iqod/kZT4PfHu
Xysq0LYJNIsoM/k9sKCJCdWNZrhjbvb/Q3lm9MN+Nvruxz39atdeo4kj/tBOEHtE
py85/krtb604bgIZT6vHWMk7k46dyXyNRmzwxRA5m2VnPp47lBBYCnlgUQoLRAt6
UuEm/chIUTGVNwYgsVATK9cjwMVTh0gDfrG07OrMyYLjBFK/4KF/zU/3bkQspmti
1T9BVdJDXS5yQUc0Fald7Wc+NF7YvxlOA95z3EM+cihObc+N31jke7s+64ptF7zc
fADSC6DfD4zW3Ma8iXdqifyBSgcHKwf4MdShQe5dWb7VgLUNjxdreUYdl4M5Olc8
yOw4innSzHafSRRj3nCGmjx5JL4FLmaCAfJ91qiGdBPdThcbcxknINKpIUClqjve
sQOdPbqetBXRsvkYb22H9yzkjhOG6KAPztNpsfyKIp+qoOmIdwjWYO/nZUKpTWE+
GhSfIchPB9WfqG0Z0AfnWrX50GqcuQvpFX8Pad1Bcr7gnE6wKuRoXiKeitkZ23iv
lJEqj5lHyX8r8WPX10adyH+nwuvAavQVwYevVnGnbVy2HRaw3ZTO/I04IBAa97Bn
viMwV8r4PWix1XlG/b13/nkDh1XugOZGDm3TRBou61LEWzyeOkf48U90n5Ww8oNy
ruCRWBafH/MU5zxz9mnbWFsWw4aJkYSUdFaNvCeFCakTpCsICzsxzlMDloWDEqz1
ubjJnURaxH48IYp9kriFwA1sQlXZPJ2bedmMhPaywm2o/JGSY6Ks5EljeF/mZxB6
Dn67GNb6xr5wDpDv2p/FsIRLrE8wB8mh6ZT38Bb7eI8e+s2bPWJTy2fcXXZZw4tg
SfE/ikckQ1lCPP7+Vns68TrNb/taGHMz3iy9CCdn6rgOkUd5fA9ACTUAFtneoz2I
KfRQV3CXOWozzx6vmGTWEW0yyz4PwQC16DYM5dHk/zFBsEc4h9uJBNq5m+m+biwQ
w8V78Ub10OmlEdDI/VbwfmE11YrnHfDx1/xRYDwV7FY5xZ5VvQFG3yCHTxA9qbU+
Mo6opJJ1/bUdkb+URyJ8ZFoZa4cVZrt5LoWzr2Mp5j0qrZZYp6zgHlHkz+lqaC2E
+N8KfOB2AR1YilAYmCg4nfgc/+8d/G9h3LoWIMsZ6OCf9BJScOF2IxPoUOsQTqMy
LvTSNgvWjykoSGi28AC6YheuJzfXISHzre4Vk2xqom/VmM4gv2k61Pm8O6s4gmp5
PFrO8iStbnM8EtfWGk+u6RMXicOE1Q2FaXtYwgNXAz0iMhLLdHYKWAc5h3OamJlu
HutnTey5H65kBCxcyXsTiMZnMGkASYMSozuZFpXzItyyvnLEVP1AobgNRfx79+f8
TNrD7zCVMd1KF58FRQLpnC59e1GFKxsLT8vgtqaJ5b8fxQI8aKC8U5vWONKuVYxc
9DgtUdIE1Wpyv+kMaJQ1N8KCD13jZs452SnawNWx9WMokfncPVgf6Z/urCI1wgzu
b1RSsV1WNfajijghgw1A0W+/Bn0yDO3/v4ZGViwr2/OoGCcm1WLNvtOF3Y5Jriqk
t71BaNpP6MS/HPa5gnaRmqGQyDEFN502YGUVKPnQ+oq64wfMtwHIrJqWsn1tM7x5
kC8eI8wt+CTneJqboTnHE/qb91Ac8RuPPqYgnbKy8Q7n+K0hBm+fYXOnQbMp8UNQ
d+AMlcql5FF372UX4kaZxuve5fDJME6I8uMQ+tHUxyGWvImlq0zXKysjRm98BNbf
9a0Kurd34EmU4/Bfh5n/08t086J8hLxRFvB9HHXv2JRv5+XDeR4sgcf8+C/PONHN
Ay3FbJddKgVCVB+oc9rwOCSnPjfaSiiZAbjJ3yYhrjM=
`pragma protect end_protected
