`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jOv1suOqyAf+DBHw+CaZ3MntHXMSds6MzPYUeFWzVp4i1DHb10MJItqFubK1JMYB
st3Yi2ueMCyvyqInDUJINbYeqgDTROKtKqppq5Yu8QK8dKnerOq65FSi/2LURqkn
TD2HfBmwoJz0ViP+7KmkEM6NlE5zBmfh0FtNx2SX08A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 45200)
MQVNwCqqHlAoxlZh8IoyDbBlJSGkRgPLb5RdulNZLJmRHZofR5aUddXgVuz83/lv
RZrWXDlJFcvPRZRRjW6z7n1rg++eOgkJpCpKyUL5Pe+jJ/oqHPLXHnHV+Rl8Z5+b
BlH8EqkTWFUYb5xHyg+yn51RF2+PBSaPLi8KXKKVxTM5ENOYKAGQGeOn0bQtYe4X
iChq16VeAVQXJCd9lpc++eipPNZuZc7PkEzQ0NqYL9tT4Ho8AAmfXUWo4qdmTxbE
RycoZMHlA8pn7nuvAwESumkl1jIVgp2nJYOiELVzsZ9dY2lnRRxs3CKqO9MqPx8O
dxtIYIyonCJII6FyYHh4AMUBjjUFZZAtK2bwtyzv6CeJHQfwIO/V5FjGjb64kK7t
qSRjpCh52qZO+J0+TIz9icF7WlfGl2xM1uhlitT5hNYogt/etHY7T7rS0YjMwUZH
G+iqhSoI1uIPZGFcIdcDePysm7TeZgyrplp4hL+ybIZFZ9LFN0QQuVdZ9nBGpgoX
UV64GHGe/9WNjA3tjrGyX6/mcQbkWbCBay5MDpl9K1Xbyk7mZVVSAlwOBBiEVtnP
KkFPuaQcJNFOXKthHtR0ZbNZaHVJzL8dibnwr2svx9e4zRzsxVE5WWaQ1Hk2zr6s
8lipzlP+znmt3IQ93yTb+Q6p1S4l0N9unN3WdtrBuo0GLodrF2xgTYP/uveIWvfS
P9L24NhtGUu95d4ZkOIweGZ4EihVp0ZzcVrnHH81qDPUzwvpHwLNr9bOYCogJ9p5
5UHKREo+GViGaoWxqI8iC6KcyDQnOTsZ+V360jTqhwhq2/fR5devrSWj8oJ5G/uN
uDCpCZYM7DCqsvQcxzjC0c+g+HQqutNfcSW1CEAEsi/JhdgVs4qSPrMF8YejaMXa
TLpePnSA5LD8CXczSxeHT0RTxscFvNQh/WlEIHUy9LIWf2qMC0M0S+5dU5M4eZce
yTd4SqixpRyFQsCUrOE5NcA9r/zDmA2a2OlmiMFiC8xDAFb6beS/N7ZUW1DmoEXm
qD0Cx2aSB6j8ugFyIDK43A3cje+SOChEor5NDJp63mlQNtqpdt8ThiD37I2f+WnR
ZRxiAUYxm9BVTfNQdtdpaDsXEX64a42ntqK1OO1l2BMl6LX674xEw5/gWt07rWoc
0sDIpRChaI+lBah4xTmf7QBhJUMEDuNUStILjAcuT+CJ2krWyL5kihzXmxrm0hVT
VrotoNxLoKNaHLQRw2iWPwrqF7+O6HYH8lxn2lfj/ORqf/Aw7I85DsgS+PLWyj+e
DLweQQqLjPUdOmaj5GU6jqM6Gi+Pb+jN0SFC/oWJRYAKbAD4Zk7iCoPPjZAXMo4C
uJ3ZhWS8e3F++13xwGQFgtQyQkXDWBXUh0oDghgIREMMGRFXlU2F7fV/7FKWkUz9
1guHzKHpLCgk4tBAnORqZo4BYsykH3noFx3r+IM5qqSu/BuJY1IGWHOKPiGdGakL
W9mUjK9ZWqc2BpdYFm17oKIGY6kxt16TSDwqVWy9fzEmKw7YR7DdNc0wGFai98/q
f1gknyr+YnNQ3CzzIKMedX3WnfqiLbkXiimiyK6MSJ8DR5BhbOAnT3Z3mlLpz3jS
v1eKQWylsLfl4iB3wRgP1av8oxcLnEZFk53aGb0v/LUT+BHvz0F5rQt2YYjSJVez
NM6ctIFgMVALJ6ASTgZoDK95pBjvn7mbaosOZFQvmqLFWALbpQSnQobwegOMnedr
AjzDM239LE7aZM6f/OqXbwDfPfZJ27oRnpZTtW7tY01K2AekgF4SNEZJHiK082rB
carBja3dz714Z/Ritr67h52nb+ee3yuSnRbeFwsXDUHcz4Bh0IFglG5HTvahgtTC
/fcy29c4MIAI+KFAZwZhB0Uveh/N9jymbdOb3f95CdgWa4mXvmxkG8Nm3fcE+Qjn
dIBjd8U9NUbMbtB/BMwDSXxNP03yddX13+B/Oc5i48ha12w4K9musV9nrOzTFWPu
guxIwtU4pq3Y59c3qrNztL3tckV8vpCiDOJ4oGq2g+jjXZ8yW0/RHsqJh4H2Crjr
YzNLxmpDsYt7ESmE06U1dzEwjE7tcQsXNMzl9Rjm4PzJSduH4V2iy1/hvVk2nL+B
7R+rgihndZa/0eja9sJC+3FGWcRjhkjKjL2A3Gv3BYiECmur8HqbxrNCbZlneVnr
WTgsoVKjOJ5wXTv2mciVg9w2bvVYcaTZC+1xluEKzqMLv1NiwsJtsYIJOke0b62w
XMYv9N5puKf6qe/ug8JgrXg6TkV1lBl15aQvmwCX7edq3wBm0rzI85ohnV1mF6cC
wFMXiua7jAdHaeGhRZkLTv8vpeBmxV01v0DWWN7Qi1lcahneQR4ip//t9RwzI/v3
gR0z6bre6Rx7jqMEie1csaDagR7p89t3x8UWafllFOtf6j/dCVET45zW0dGRP4rQ
IIQOz8AUMh0nRgFWu+KvURyhYXV7H4QUCjDMiRF+Ub4WlBq1g6KvR4UuAo4G5FYm
iH2wFufrYFutkNkj9JDP5vcbZv4Q2F78axHH/KjFpMiK+eClNA/kQFhUsk04hgm8
4utcZ21HdXDWQ69pUGokMBo2/oxEVWcuZcv++nLS1BmrdrmHKtp5KSOBY1WPXRwr
dHHsHrU7MQ8C8Np0KlQFZwTSqUL39evT0KoANwOpLlqPaTmGWGqNhOhJN0PSTIPJ
gkpFxE87abAyIqTOYsNeW7uxytdijP0YnGJyyvlXRM6WtQmXcogy/ZhtcQIJpyTO
oFkGG33TA+cMwIpegIrXrP2yZ2KQIcPi9FZy0hPa/mbdNUM+SsBeAIvpAztn36Lx
l8A1tzjAaRjKOHQ7hfTcEpTmbtClraTfxsdFVUG+ocKSkw1TY1RIfstUg2Vhsgt5
vutrUTP6E21UMEgHG4F2mk8wqXnkQrbWoreTi9bATzbpSAC7/8iGYG+SIcc9DBP4
ifwkIaS+eRZkdG2uaDwsnDechqy100Pskv5Dg/8WR9utHo/6Mp/JIK7IXNTLUfLI
T6SjkutV7RxeG2HaUXBkNN9jw2LqSEQ3hLE7ZC0/auRNjzky1UVqwHx9hsSNfaHx
tgp5IUaHDQoG6T9MIPkNazdcUXklblzxOfojzUGkEzZrv2pjohb5CbdJoc9HVdHj
GaTy1BluLXE44OYVYyMxMtsxyEYf11hIl+wFDwm94+rbsc+WZJgfYtMnDEUzZQ4l
o1tgoMZWqCT874sOXdkR112z/Xdg+0IQZi2CyUzKDgryoBGev6mO4pn+rr8f/+Xv
qwzr3V1eFvBLMGFrG8aV0u4mJQiTEObzrzZJXUB33QlGwE0uH6iRokFkO/F+FTrO
eASgykOw2WT4QcGhwCAk2AIzSb2LEJ0kHCSn9qVpX4MYvHVqTONAu8l5iM7koo+p
J+0ED4/9ML7ILNAmggbstE05AUvazMfLgAhmpzw6NdTuk89CLoVk2s+AdMUvCJUA
DaHm008s3nv8Bl+06P6nFQJTx1cf70mRwKAhiMsEIrfXnuJNwd7B1jDJmlsPr1ZB
2sg37MYMWn8E2R+O/hm6g1wSrUySlD31LbmCfw2H4C/PD2nT5DdCjjuxf8veeuHa
brexhzi2tzSL8qzcG/tRSqKXVWn5kPCI+joDAck5DLbJLznmWRGJ3TgSV8BaL+oX
zHKlJSx0c6ZPRMW4/BQFu5wDmg6HQfGjSlbUGtRKf0b79W0aLc7LE6DVc+Tdjsz9
Ugb1IPVkWIRE/zmCUzkIKuQUKagOfeI1gvaGYAKv3LGMqLrWac63jZD3Gf7yArQk
mwepeQLX2MvprgABagIbLhhYu2i1/voIVD/BLpI8anRNrPmY7yz9AZKOwFya3Y2x
ywjNx9KF2b/kNBpf/Goz1a3P1/Dip553sIISfh1pR9BgupdUTOCHIn75NP6fpRyp
9KQvdljuMHmENIKgZPrZRXkNVlnTlD5h8YzApqTi9CZy193qSgM4IMZuTSVP4ebB
JDkc3B6wmkHHNdaGvUh2EPQ+U7n2m8G0lBKiCvwMwcQmRvbFpwjid48aP9/C9VZe
iSfHIDyzFQgbYb56lmb+ycP3T+5PION2svl8hX+MGJwJPRyT0tdRoGqgYOhZRM5O
e/Gum6nIFPlV9tAj1XN9WgpOfYNeQF/q44QhZI1PNgKQzb5y5iROvTWHg5KAOg2P
4imFOZVoXfTdDXMR0xMZdCDrLPHvtg4glmhTlvH/24UjJ8TtTkQq/+7dQ7sGGSJs
xkL2vEGbtDPGHrQfn3W4yQ3RtZ7VAFSWTRHgoMhtNT9T5X28EwfOSEq8fiaRXUqN
CNMUBBgel25MJjapBjQScvqTmJnsmUy8Qc5qDBjcXjypCbO4e44yC7wBVlThhM4h
yxRFzdzaN0Z+rcRXk9iazGXTHqCVbC0lKHwXGN3mEyY8bFMhC6OBpQLmg8L6oiGC
slyP6VlGJr/NyUR8SwUrzGERjFxrvuFsIMdtS1C3cErZee+Z6rIQWUI0q2gsWBSd
0PVlNzAswxT+uzV1Lj/cbvWJgofL2ohllOUqjoPjnnGcLz4uHGbFORw4OTCFHE43
TthnMU0YhxU7Fx3PWCygUk3BxmDZ8Y7hHVDzm5VOI0FshqWVEHkEYmqF8x24rQxn
4jwifRkZyoNPyjr6Uw+wOUPtqJMWAkN1RWOSNykz3lqwsvZijZOfIPvQPktUMjLc
h6WmH+z6y5TeRjInST++zHCUSfa2dwwj2eYlD5px7M3jx91jmZkB7qA6l2+1Ifcs
p+lrkJBNVsDCbOTojJ/XYbWzZ4C6BLFRW7ADyc+JgvVMG5qxNnM+aGC4rDHExxwY
7wxgiU/8kwsgl2WObyfX56gSkqJ7HwvExpqaxDBTDzd3bSXVggkFR0BS9HS6Gw4j
saRcKhOO2ON6YUL59LW8f5o+2XYU50iyMbHyus3m4fu9neOhIDHQxof20DqlZtJu
AtcZSPp53qgOfDHFjaVTenhcxY+KXmm/6ongiRkjWtxnXuGiEXk88HCTvF4Ij4y6
aSMFaJS+oTroSAmUPyz5o/dRxYc/TfcR+eYZ1y/yzXkRP1vUVYy7DDDa5xvrq6Y9
3NjauHujjmdbLUY4a1SC8BwGtjpq1xM03r9+pQ8+uhFp44EYdajCHxebBtvM5XWG
ntGRFbgR01b1HLVbOM5Fit02QOV8ylHlaWcqG4St+CNuxSEtDDu8LnubU6rGK+4i
C9zG0+7mj/RLIUoVgnI6oE79uCOgdtwH6iwx0+nnqLkn6W+NT42nLpURkKU8sT9t
9E4dWKc9Y7cYgvfJXCta92C7Zcpn90OTubvgZ5hDaEpjESGj5t2vBpS72T+ejxzR
uvA2HPM+jWSnqB1VdFbcQRrQhHHdNre16+K4jYipa1IfOf+PixlGMD6CV1m8Dosq
cCTK/AibgulsAQmXOhKAXK5nC2Arx/16X+R7ZgOcxgnXT5rAJ+uhP1cyl+5pwlHq
W0yNj8yEiNDFqjf8bupTtBZwaGUUtcxBswfrAg3hhrWqroScMeGuBDR3LBQd7I0L
IoFAR5x9zYVv9V4BMB8KXIl6lYYvqGmm1IrlRB3LC1E4sLTtV1rTbJJn2hmRDMdd
xU0BABtBaRCSl9N5rlSURkzQPzE698UpYsQWTy/Q0h1tASNOcbCY7Ilv513OCMjn
EuPNRhC01EJePoysIrP89CWEy8t6Kg22GkWkj0LSWi1C0vDK26CZ+zoJKko2DckJ
9eqrkK6/mts32kT0fHuVj/Ak3BSwwnOFLkEKt0R2VLVBa5ucnKEDGZG0+WFSyREJ
0dhYc3xkY+Up7Tb6Q8GZ25yjALk+NqcB6iGHgWaTdJjqlgkBEPwXCMBvN6yiPNwY
bsD6chNPz0hVBJJZWFriYrmXHHOqVO1VSToFRBXZLNnT1XQmwb5wSfAnnRJ4XHVO
cxqpBu+ko47F5KaDTl1AXUOeRA5CkSwltb4wDaXqmTthDzHZc9oDzj8bN/HuPkhq
dXipEFr2HvUG8cJRYdc3vQXrUtObuuk+4OHiYmQqcH/L1n6n8HOwdCGBIWZsr1jG
IImhJUr/4Is8z2/8NFb1kCEaE/TxDK7zuXUXafPjHvzRJ3wAcMPjI5iqwqV+OoHk
6NDwH1PfwbK9p4hm5d1Wvy3Zo9gcu+O+qMzp7S0eV35vRNh1gyBEUcaBMgC7YG7P
3ZyP/CVf+usdwczJM4QHZjePCgy2hSXbxHfRnM5ipPonLhLS/mp6KdMgDHAxqPZU
bqqZ7mj2WzgvG1taUMduGfVw0Qq6C1OcGrxm33ybMoeaCgvUCy7RbkQAh4t3xrqd
QcpOQE3QXJGOGQkAQ5+1zdY8QPdA80oLhLycnFPoOJubmKT98OcNm/byUrxkEmvB
VszupmOywep2VvdEeRZkj0nxF4jRCVxESZpTFBUvoKjPijFzKFs2ONdFWdlTuBUm
ZluiLCO0KudGWcO1HRE3k22lgnTp7kdSarm9ve2AqgBY1E5PcPC4bLzALqy7hIu/
k34B104ocji3C3xEqWrbhV+pQ1MEgRClQryvSDcVL6eBa2/B/G2brB9mYuV9TcKP
lYK48DUNHuMsHapZNfmbGJcj2ib5lw7gG21CEEmkWW6tsHv63sMLWf2je95KEHSw
4E3dAUElNzF6vAe1M9veraVykNbpwFC0AZSsGwod5Um1EL+SLWtzVJaRtH5YNFbc
yWJcC4oM2gKg0cZvG3qeAvEiBVS0fPPkYkKe3YDog0XoQaG4mqbvN1ZFNJDPz+k+
cfgvZE9xu8aQpQ84oa84pdIQLpqASwwOtWW89WpSvKxVBpKii1l+RV2Ongc8tDi8
Tgk1PjbfGFo4iqflhR0djf8/4/qoK82OgLeTekGQ0BOyMuMqbEhgpAigB2dlIlgv
aRZa+qlQ3qh7oWQUD46rPC92IfpgIgI+/sZstFY3rHMo/8bB29xdcudBEPq5EQiu
cyhmAfEqsL7HH0PzDIWBCHW0fYBvwhRljozEjds/n+v86MeCHdcpA3uige68JUEQ
a7+eoXwp2nkwTjPCFJWelgDKsDqr8HvRhiiigveOeaWolje4HvUEJIowcRnzyyWd
AA94JyvClPk6MGKjfbfEKSLjfcunJdHwpxe8mUlYe+TwQUZY6ZR4S+mw+azQB8ys
9Tqpr6DL7yiW0btZ+JfYC9Y/zEFHaLWbvQDAIMmbwS6oWUSzPl/IuDVMMRPw5gJS
pmw/T36imJAw1gFdt4X8+6/3Jlghyd7veUSPvGltCfvsqA0RAl3H505Xh3ZuSvHe
C5vhodL6c87e5IP4JN1EjREFBkk9+9syUPqVCZOSmBJrmluwQZg879Imu7pP5l4b
+GnOR0s2JLqK/eRCjCsRD1iENL79WY22aHa7AQJFVZfni9EyQQpBVOboVeWjuZ3O
Rd9VSmj4c0oSjWkcHcE72kRfgyfelFOOR81VT4pD7bvNAO4r/5R1oXJL1S55P47T
oK0QFtvzBAFatYwk2/P5WW/fKfBIAQVQuxNdfKoQgtFLqah+z4OHMDx4s9eeqKNT
nN/GKogDMrq7UI85pXHr4s2jhgu7ZZBDmPKJg3cwyLYf8VLLvx7/5X8SyARkrDI6
1hl5T1ylsumZu48lRlPwJNKApbw3kC7Tj9sCzu2+tSiijwLg9UfmLywFmnjJkc+t
aUEI6CpmgIK0BGF7kBkrYqp5aavtGX3yYEmYCqlRW5UxSwyASANlUmEcXXiete6e
mUebdpKEXDn7o/yNFgysz69hWOwseGU/Be3Kt/nmwiKjHo74CFEd4N/gIrTOUH/D
RM2WQmaFND04oMZG6fPpAwXmGz41rcQSy27E7nc68uQsCLpj9W8SOFVjCj8QrgQH
lE+2rCWtpqKdl6F9yA2K6AdFKmFYccSqSqIZ8n8VdJPlpTl2n0WB+DL/VT6baRGz
vN9k56FWzNhUc9ovAs5+8arFl+mpXiOTHyH+vsNgM13gmRVrmBxXoLG26/6iNnHD
B3SrOzcZ8IcFj2DMaISrqilZDdwCZiJqBVLxHmj6NNfN0sT9XbdFRIzY4SPREbb8
ZsLURdgk3RNULfeDZDXFKS/419Dg+h6MbhuoOzXtqczDByCUBO4NFw1KP5zGizUj
JEA2naoqiftRqh6vLuoybHrLprZW1R3elJExKsGFqDT2YkhOS75+GyPpdffUeEwe
KwU9JrPmWs68PIasUY4sOBzL4nqNc/PaZBGd3APbcJ5+Tv0Y5O0NMwR1oUUECnb4
1XS+9ISh31rJqTjO63A5PxAhI0m5dFE6h6LW6SpdrXrxin5P4xx45Z1u68BUUl5w
sqYIB+2Ucqjysg0jONM54Hfcy7EQvAzaqlyyCFeSOSGACcMyvlyFWob0BJ9qIG8a
UEdKfZQP5JM3TWdKqor5heGRvvLUoQ71sXIcTi+GruVsR5OSQ1oN9kwZLeb2snXC
M4KsiD1e0V8KshCdXfK/eklG2KS42W/UuO40yFnTs1GIbme4gTGYTP2qQa/ryIkp
QG/a4iMZ8SkO2LrzelHUb0hqOzzBgsbvmHzQ+HDKwt6flwqOZ83CcPt9loNDwU/m
GjXU+Nzy+Ahbb9a6Wk34hGdNa7xAgBW8eQ0pVBXRn7TGDoG8KR0rLUvs5yW+LPqU
INJb5W+Lxpt3px2P+SjDY3ctI4XDp9vfFZ8ajc5WMGBYAogJMDMqcJ0/5WwlNQuM
ysjtMegJkwiihtf1fak4ehRzFDlPPH51SHgCjLMOQ7BXwyvtVmMCAiAxTxEe1LXc
x9RermkkSRP40d6YRJe1IjillqLJdgELyHdugrQTkvjp5ABqBjsxj3El/JOlrLV/
oGDa3tLU1wLs1QnxN1Qkl4l5GB9gF0NjtJzyXGt4VTMErx87Tr7Y2W+CRdpRNucO
1/dVUJwck5shPGvLFEf50THnKbsOikNW9lSiU2d72wAba20BGC58UehQnFbU6DiJ
OazZrAwv6ixU2EQiDvafzFIz3dRuCKY/S5C7bwtYHmiTwsy58rkqxKqRvnU7zljv
M4NccmNnzlZ6BmacsEIEpOiqKOjFB3eGcV036+FUIWSSoMFmjVqaoYyXyem//rGh
sEsmo0ktDNpNRZNpeqBDS64LpEnQAGlgZz69YStOeaoq6i51IDVrNItLE2ODopZ/
Nbj4a19SYk1ckEBXiqTxUsFV0B9FoJy4LA+cAMIAhF5UonUYHSs6pxdRdVRlQNx+
NtWpTK96mGZ3cTmWeBCnepVepil6RF35FjHHlbuRLQy1IICWNHenh1CfDyn0SfX8
0hNwN49rbYY4XSfTPs9VwWyvEH/VVC/sNkXgOoyHeu8m1JiVKR1DQEA0gED27FQF
2vKpkK9GxosiMBg8LJdYTNZ/BwlvFMfiy525ZGqNQItP6vsJWnzG+bZQrOcYRIvS
WbrKdtAUNTmENNmsE1y++Oz07F/8oeKdSqXhu9fhcha/uTWsDpQTuSi8gy7fbZOB
Rw4xALBp1CdPNMmnh3KVEqVUcnbqdjsRyxezvr5lruCrubfdYqlJZRBS/INbBuvg
tz4DsdW99RSwO9EJVUGE7ozO6IOX5MiD90bYQv1E5FE9MdCgXyLSVkAhNsMinWLK
gCuUrltMnQF1AdBTT/7sOfFqwVfcR6DRC3MxGelnYmdS4AgZeZOZwIZT75PSYnrM
8KhcR9ESBnY7JAtCzsejWE4O8IoqyAUzE1JBlqR+YEZh+kdP//8YV4akIyVTSSZy
muQtczWTzPnydwGtKd1yxKlMwksCHywf4kEiUOIhsTI6bFvQryOezQ5wzrAxZ+lM
QPR/VK7qNeTrjVGISCEJQyG6P1XROXM0AZ7/QwhiEV+oRCgrtQBMTq1fNGa9kPq3
CW9u51aR1zw4dM3Uxmt0RslqLxr18nMOrvVOwUP/T0/Ugut92q5jZ/YmezyJNS8v
Xv1tFi3QA/U3HqFQsNpoLBzNTc85nqV+yKbbacIqzPchGUrnWzJsyTtQmFo8QOEe
IELEt0pID5A/8b64jFDrBA5S/en/t2iJse9GO/qz8/yc5c3X5gkdJcdlh8NLYWsv
xLTNjwTeAU0KyFdO0SpUW53FQlptKhjaUeH3mpEQPLWiVcR8D/Cd3mqTLKWz/etf
7NFmXlX9skJ8mkZOMezGyVRidz0VYp+NR1uNcpstLqg7h+CjGl77/21rfOt2Tmbg
JqVI+2UyAc96L226j6m9+/m4985+0P8eXT6XC3eZ87F7JwKRiDm6sB4ObFjZ8T3w
TbO29TY8EnBIo4d6mHqyJoBBn/j95q7K7OhP3y1JjiBQQJIYs3Q7xbnEpXy1yM7X
SDl5cF2khnGO3D1v5sBMnZPWyFeNJs1QNJt86r5usiD2JUrFzEldeGcLhXQT6ZvV
4FV5Sx0vU10KFiN+JRtEWBUzYJCNAPuTIlMBewEaGHLnHAp6b4GZY8HuXKU6qEST
1q70SZ036sNMMunO5FBQK08cMLxM6SqRL5lTpPLpooMR0YMb6l6Y4Pr5M6BFG34r
4nD89jhl4BnzKs2Q3ZJJ1s8Agw/VqdrPReXrDtOJxkcLoIF8C5tZfASFE8DvS/al
24eiN3mNyT9o6dTubzddovvu3MdcaOAM+EG+WmaXioG4udk8r9xOjWFpw2XJSet5
bDvNhV3sKLLM52n4QE2dCyvWIrcODPwZF53GOt5XXWZy+0x4XGj6FnrO+YQA24sR
RwGEAMavvKjuXuP4fn5Br37Yh825ro+VvRuOoJ40SqqEVg35rs8XzUgwwJzRhEb1
CCl2r1KNx9rzOsa4lFBZ8lXuXvwX+VNs0M135gBDHaV4txP+ojjQyMyicqOcJXW/
Jhcqw6hC6ClezBweHsApMIMwItGS4sxVdThJrRmb0isCnJjJ54aSVbjOUc2Z7Hn9
2JCFoDChYdWwzduUrH4530z+c6mHk+hcfFNvI74aq0YyD8lx9dW87Ati+BnS8mrJ
eTED6mvO8h2uThqBIj/ZF9l8hDWuKPKHn/EbhepCaSOjJIe5KboOUALoTW9ihrMG
Hdy/Yw/+vy02+TCNWr1CIZEsnAEkfzWqedIBuKn0HFk+lHfeeAQOWUOtoe3flOPk
c30gCuFC3WqoIlGJnwK30Euc4gcc7eHGl39GyH/zwBcCGkuh3RfZiYl6Yv9bg9a3
n7aUBrR0lRu6zQso1jU92aTXCSJmD7KkmFMTvu06RHoB34aygECbGFfaUTovAPa2
T9+srf5ZqvnG4jgfy/CHK+y8M9EZEnj5vufaxPP4ck8LtGRZcdbeaPnMvmLRgiIv
vy0V/X9r54aww+sPnb5uokCzx2vxbvE98Tf61/pGWPWvrpHxmqeUF6AxaMDvmlGl
XlveTvrBbO3J94H+pDsfTf63arv8JDxva28TcmWKib3qJOQKYQxOw6WbItM2P8wb
cQ9Nb6DBoi/AOQ0tvlTUrhjyUONb4TwvEeFGtCuLWOEkBmKGa4M62JDLiKAyrM6E
EPtipWhHc6wynTJDo1BHXhKwu96ICDzV9UlhPZo3YfJiKitZGlShvITSlkjxFwu3
gMJyf88MfUJy5mlzS6Qm/dPvp3QhUdV6Af66OCUVY4TTQCLu8hsoPlN8/baUGbly
+GJnAqe7/aHrHMJdEIsJefsGsj50rtlgHZ/jVwwa2PPf5L3g1Uaqs+tG+pyx7c8o
2Ecj8ih/He3lYwcZC0vnqrrUfVwkI3nthoHt53unMOt+lT7Jw2aJFN99Bf/k6R3b
n6w8xn4cMwQ7d1ro69YMu1Z6Oj+te2+omqhABRpKHvJrT+bIsFJTt4UTwORawX+w
jmvFheTaSbU+kAjusUbjvAuh1p6HnEA/X9fLKMzfBneoNxyxB+iK1EBFTSCWEfcY
vQqNI1lZE/50M7OKP1W7RCmInAj8rQBLivgHCFCxGAkI06oy+DY+z4E1NqgSB5cU
0lFLb3qBDgjaT6IGnSSJiLm+/NQN36de2bidgx/ZiVtZugukYapHEiTAriQ2QYIa
1tgq9NIaSgvq6POL8/8Gps7rvi/12CsMgIkFWx5v916hVpjOHRtUy3i0A3Hff+Vb
vZN/NiNIAkB//V1ilZnPMzkTDw4NTaS24Q4aTxh404gBhivfNPEExzaw3L6/5OMc
VhDTOYZoica99PfubNBWrFGhEOiG67Qkp6TfIPfpmddqt2XOs6NZS1L1J7rlX2TC
tsr+xF2Dr1PlwY4syUARmis0uGqWgtDsf/Rb2p6XIx3aYOshzidAr0NlIaDoFnvm
AWa3RBoaw55KWqvmy9qnTageD+gekyV9Wqo5X53SpVYGg+8CO4U/rXF4t/Jai2XA
/0aoW2nT24ljqAb0UvrdO99+beeuTaNO7Oxsh3V8wi+rHLZI7tF/SAc+jdL3nQ6A
ekdxopfiMqdktbN3FXIp7Oat1lK187VcP88KRwz46Fd8MI27Yk6r+hs6TOF2phSN
ERpLSJ5MgnZzXKARHZhVyCFB2dyHqqYqLJsV3r4zUtONbMdFBgFwHbUeIWhhF8mq
uD462nUc4CgnE1SX73cv64kos2yMV5dPEmC4osHViSQsx37Uaz+ysslqpQ/aOhbU
68yEOHuqhIKoa26qXumtJtnScOxnNDaZ9M+tt3GyLJrIHFGM/zFeCHirc6LRJHyE
gYSGlcZ7d4AIBOP7OavS9Xo42ANi2jZ2f0NddWQZFK7GeGgiIF58sQPTOeCFtCMz
MSnEMlrkoDMfar5CLt9wsuJU7Ib3sbMoNoOqR2cOTS3NhPIbm94eipDu9P7yIifJ
nb7we0klqhde15Wn++wNucfsu1DXGaxoZgyqKN9YKN7FGbUks+GFm3vWKB07NCE4
e1YRmWvjct1uftjapgCBbYoPEta8Y0Emnv8SqWG4f0JtOWYhmhZRBBrdHs/1vHvm
AfymhsD2LsdcMWxaunsa5NBxJYQoJlYV12doKZvXFAvH93tPH0oZ8AReeFSpuOnx
cfWCwLp9mH30Ao5U97GmaOtH0NH2i7KLMdzWUEkXVm+XfuYGkyqYewJtyBPfX3KO
pr2XCsKZK4RgFY74B06c3GkPBnyqliVgyKoYaMfbtOa04ndmQl7LfVHZ1R1lTJZt
8sHjdOdx5Iyk4wXcIGEAkuVs4jYfqbVu34KLNlG7mwFzHqxWhrtC6et44pPcIwEZ
IRvkbVEegHFypgFHIY4R4Nvzt2wfkFPLSl0VKmWZxKYjcmaOy0n5gQ3jHngbE9x3
7SzUI9OtTD24q0y5bpBUZSLsywNXjQ1LDVZ4x6S1FMJ4vMHtb8sZ6kPXdCHJ8EIy
SxWPa4AKLBd0pP6cUbVZ2vDu2ZhHszMvGv+t/nd/82kBqBdxjlrxSupZ2p/KCBiB
OjloE8JtPINN/+eLBWCy/o4LtGBgB2kSbhxXbnPDGMQmcNJ+DPLma12Jy5FGrOCv
si5o6LkCAUYlli2QVpMNvW5Wbvm6/qEZNukoYoV2zSQ1mENFYcohNOkMIpsA8YRv
J1NIfT+Js9mGGuG2z+2TJrrYhSF8F/FM1BZzkyyaCELgsCY2QbUHGIhSlsUW5s2v
dE6S5al+20u9z51ZUqls1UA+A2vn7wzfK7ocvXJ7a4HYhN/0Kqmb7fPhUkeD1Dkp
yWVPFvSO7CWfQt+mnJdpNYWlMPy7rdW3fH+ljwMG20maCyveH+g2bUhv7cuwZT8M
8yV+CX+e7T97BnCQ9igxtGb2C0wbPjn+MUS2lf7ALaJwImtNPct2qOFXFfbHii8M
ZpulNypd08D2cGOiJrz2UuTnwspavzU5yculnFP9ZTpMYZ7vcLqGU4cTVwhKlhnC
zlw7734+g5Z9kd/S/p7vvniyUq81S6R/4cwQYJadeAgYxKq2L7S2ltWm7LwMK+pg
8LOqKTUVjhfWXuVXypriOVvhJh/XciLF+RHaZYl6+vE71vXh3cvE1LkganGCfN0q
WFB1iMlbVynCtrhP4WyQK5n3j1+YqJXvcQiN9dylDXvcEPax0TYjCUA7b5/VlbFq
i67OGJEjkYCUR9IrRLsME0hokGHGMGTb3S1LEu8bWZsKzBBfb5oE9ywm0EbyFwHL
eT1PFQJHox4fO8BNQ8bmMZB2yJEJ26beBR4NebztyG0hlfYCZM61iAeQXS1n1wND
kwQHO0uLE2HnIp4T+rguqGnn4ISYLBjRe1jejgS1bjx7Ac7SF4rtWYEPESAYZbxY
MTftVUi0ZUZ5aK8GKB3gvf8gccX9G+Z/U+CdgTzEWcmg/nQv4ErdarBUuC1m11nU
LaOUNd7WB/Qgkdq7Mr0LX5vXG2lNPySeO3aDm+ufOyjewNUeZLVlu5G89KNxnPrY
g/EdT2fShoGZJqk6slhD3x9u71+Dz0datoipZAIisKzU2Tj5Zw+rvY2fz6Ht5jNB
bxPg8s+bRoOIbXWTfH/q44AZCzOjWTqf4ztR/B7LIvUUnbhTWUhd2zCz3SZrm+3G
RM0Mxbj3NaMvKI/3ChV6xCRMm0+1bNMiWkYaKfoQG6yl1vfeCVnwgY5d8KaPSPzB
Pmmdjj35+x6VQGeDerS+HISUok1YK/outuk1Aa65jKl7IGC1nG/k7kpli8y17Uzh
K7xoxcx7zuJKZV2Bzs1WYbR71nVpmgqvKaWdD5P8sypfhcKx7B0I1q2i+4LbdhA/
nd/EACYBi2EOWxdUXVfk/koH0C1e6Yhd/Lq4byxg7hrVICtn2aMse6LO/D4Gpf9P
7OmjVS+pO06inVVOXJxxMnpzZNtXKq7X5k9FDGLSKYhHMY36m2Q1VQyIP2F9SNZm
4Kr9HVKxLPO4jUzXvmOqzxcNZsLH/XTfLim0LN6swzaFodlXSkcpVL9M7lGbQl+f
OWqju7oh8U/4Ys23AyrZXEHrwLny7jiNicz3gqLdycxCHGqhwi4/hIdkpfe2e/CI
STdS2AIOkG+5+T+B3SaF2tut2UB/EPNqgF+cUQ0MWDGIGqM0YWaec5ivYlrab79y
6VoeKm81I1YsSbpaJhKBui8r+KKF7ZCt1GF/wCqYv4zRFczCq5gnyTyeAIPVafmc
aiWxkdnJ1GwXlqiw0ltwMc2PPUxLSGWi6NKV0f2fKXLU2PX5EXBi9JON7X+uitsn
XJaKMKymYGrORJTPNpEQ6I6CcJ8gQ/CNHMwhgjzy03n14yG57+UTJeznbks8RzF1
WvcUC/lrg+SDuOauTKizpFRpoIBc/ezvx+ORaSjuQRTg61nwa38u+BFzZ5+ghnF1
xqc+wAEzBkAXHbWVGBmbvxX5lfxhvxZMcXARjEkG/RzY/2pTSs1IM+7RSZl8gd/r
l+TX2jKI1hWrYrL6PfjlRRIfz5zIx2UERre5J7xJUg6Ah9Qt8sap/moq8PfzPU9u
BXY56RokR2CO1jDRcR6eoACEykGz0xKhGzCMydMJWby3Yb+r4YimgPLxVpu917iU
MHX0geCfS3s75WdpYeP/zhUD/Td7w9TXof6/zUI10MjUkJq82IlkQylZOFwQkQ9W
hyA8w1WPzAS6BWgI7N+nFcbxw9j5yKxW48e2dZpJCV9JJ4EfvkczP3X3stQRHLmo
spzz5UXESldOgZFVWVP5Kw9FMcBLFsLHjl0CapbAy0/VFkaMuvERh3xc+RTqNjHw
6CwuKUkK4l6izOdnUPbaBP5AOULd8aa+mjZ5Y6bJtPbkKNuxpiAOaSXCGKY6hcQ3
uYLAwoKV8HkQpp9H7dtzxVCC1Zf+It/wCJxkDldayFpi3OkRIxkJUgO5sEV55RjX
hxt4iraxHhxxhz+Q/YOY2jwjF/zgnjehBc8qAgIkR7qeXCRHtUHpFwC+IcuedYON
jVL8Tqdyxa/+Qx8MGDmf8R+t7wTLQIID5+rxZScC4Zh8OSLe3/f72Z1uXeT/dKts
iNYESECxj1cQNvzAMpfc5w7LuMQyYObAMaUvlndMHe5G/6oShEbMoUywYxjxJh/+
uNv0c/d40Hx0BgQ3JZaMDxVzGr5HNgxaMRoesHikz0tmsNiy/p27bVcBs5y9QoPL
mlZzFI/oVPkGDCY2jyZsL8BcSCta5vNKQERrKeHG431wYvfQdFmbsdWU8bMbWu85
4pdQw/ji2euBezRCGOeszJndTg0TSlZvfoMrnTGBQnwncyiykuf9use6gEag4DvL
QVL/Z4b2AMPPrgiqA/frRRrr06VaBh+HnutIn9RZA3Howe+V7EFoLChWZQoeUJVS
nX+k74AG58uMNDtHrioiBFjqINNLyJjkqoBOpeO52xf6eoGeClFiCYY5bV/Nv7Gv
237c0bj2EHPFojS6VlJrGSDNdJdF2/SZ6h8Mq3MVxnydjDeGDsZ4jlHEpBd3rItZ
LHp+PsuEDRHz75Hg4SPDbNE367aHHvPNXyFRSyO05BqL4MHRmGsE6EBMc8ieKUoS
K5mxW6T1t87qWFjPVS1nG5DkcH8qcLqmguC8Ct9M7eViU1nzULUxCgq9BEM+7vAI
M+QIFUon2O19WGSgdnXux2vJVszjV9XpnM+hajioE7aVH+GjhPImCT8/E6NqqJx2
bhZ+i+bVczWvJI/TB1mUosx2LkjDOcTviEkzppUCqwwaoKORtSzhss9DAaWrNIEH
Kt8nIWXXe0fCG8WySc/Pxh/dy8CRSYQA+utpn/LjQXZGVNLgUw0U6JrUX6IBWlpJ
rRLyZsoJEwylaqFepU4h3ESyPDm7MpyQLQJBan3fYJkIes4TQ8vZacR2cLprbjK/
HIWirzZz2q56E+mBBF1wP5hgQ88wLhQBSyROiG7JQ0wIqwtm3GajFHkQUdVq2saj
0sUNPCaWYQQlxpBHuDneKVtyJj/I486s+xDmaN8Nk2J2TQyUB9JdZoW0VTkXfc5y
573qpMKmXZ7viT9d7l37MGQON0APU8lp0XCaH7dLbjiBiGqU8P9/IDkz1x43qqnR
5gLOcivuTaABH42Sj8/abE0ZSxHR+GU4xAcAZC7t6jH5pPFAUdUEZBMud1vWBZGi
eAYJzXY0tZ28hb2JOv/KY9DKfYmsTXAWV+e7lhv9cK+NtCGPPaxlCH44kE9jjbnH
mL0nUO02jmyZ3Qwz1PWJKPOQU03+Dq0rCtJpb8QVYmsfzGttnoDxBwoZatnL2ELR
6ORC5/JXyBbbh2gycvG+zeia4Y7fzlI/mIKUKPMaD2Yv72+GJkJKz08iPWndgbBO
MacA/CV66PI7HU9W2cW5JCsVwkzOmAjPwnwg6QvPyZrlISj1drjZfb/+S7188DIN
S6BwAfVfJ8V6WDTsCecyWUpQzW9jfgGuVjY7WJc8jDNugXqSJN04lff1S1Oho/0h
RlV0Zytgmx9kDcowG+REd1vCzjW4IGhgy/1zdaS831oYw+Fp9fWdmA185lrhO7kd
VnfwNu1lG7CIAMaux6dALkDQ0+Bz+pOlreLVExgQNiZ/ZKkOayhdwwjQM27MH5fP
/fH3954riXowDlHvVZSxu1zoiz4V3Xa6ofpb04OILEe5iPQNdu2T12qMGSdIlSQ6
o596HWqvswO+ancV23mI+W88l1Mm6RbZbWa157A4+20c20Le3DysPadmu0dcqn62
jFZ/OXlPtX6QGXWY1Ap97sLyM2LSecheve7v9C8MydKtfQwVW9YW9ZPsM8x0Ha7g
+eT94YizuzWrEUjzJE6hjy4gHbJGZo6ovJr/hcp3T6x3zzjwTCSgVcTkVhpu4Ikx
5vI4WUCizCHC8bxIox2P/qBFiEYhvtMz9+aHSCz9qrahxHavFU8McZuSOkOwXmvF
Im2vnwrOsdQQzA/mqXpgNSAq16uw31jsqwWhpUwoCzJSdyXfrsxijMF7Ijxm1gch
qnzN+h4INkL0oapZ6UTM+KpyK6anQ6BqrQALiqq1tjkAdNqVgo7l+9TD5GzeBAne
RGOjmZ78j5e5HB3hb3bqcWvkO3TPCdo+Gzj1GVu8UC3C1TaBeOXrb80UaLYQxM0B
WhEjMxnmaxl6KRtNGCgxIoN48vwwVAIcKrxCN65DTDxO6rWVHlR2yhQo15JfhrE8
6eezMzXC2zQqdTKXkb8Den54sEf87W7UnwN2lVkAa/mspLStzP8A0WA1q2U3tZl2
TrwCIOdQ9WdFotMhjotuwTUGxsjLd47VKMRV3mP7r2/mAuQGQ1jmFLZsZlF3o6U+
Z2oLY6MOZeWsVW5+TDPl+of91nu7cg2sDalTJk5/5UutxtMa9u4lc3GyKKaQZeaz
saz5vEmTJrXgBL0b+KH2Kgg8LFlMH5rbXt3t7OCRmVsz/4z1JdNFSjl8Hp8MBhfx
jeTv3NiDC4NfybAiJwL7oyzD4YpnqMqcrDDWmdcyJIif40NkEy/55+RPzQ8JyJxL
odORE9bLX01rE2Z4nJTQAfGhwTtNJYDbF5jV/jSKGZBGccbNuSad7Am54QkYNmtp
lgyR5f82v2D71jeUamwj+yOlDZDlW4jS7BLOmpD8CI2V9GoLA/NbWCUoYAN3UyTr
6MXH3bdRTkuS6sXXuAtBkySBH5l9z/UspoPKekaQhetQMk/VhWzTI2GqmerNR7Ec
FDob+fJk9ZGaiJHcs1A8yLvCYctVyjd5EIOoUoe0st7n5MI9Mj/tR8ledkysfsAn
pCyZd60aHW+zUSZDP7e305R90q0O7ITO+tKkipoYgpCA7honGj8fMoYcsNfxYGCA
2UhEJR0ZMXqrmgZznNQBMZkqnUTiqak55Sct3ScP4Oo6zonhSA5mEZi1ZNotPdUX
Z9S1nTfBBOMbKOyAbmvDrTutNGfp+NAOBSnSdhrF8G33d4ZCUJnlDWvwKUoYuRkv
VxT12iiLTuoGJsivFsIYBWfJgR8bwuxgIJTUWBHjV9Yq/uDkYPiO7h6h3EkxSI8i
2ySufXKA9b3QEDzTY5PwSxI+CmlisvVMyhedzYWYwVf4oXNnNhh5FiO428KjbeGY
n2yPcWx3Cvd2ReMVA06xP+8FNXeNs9mjjSDJzUCQgmnUqOLFaPtzF23OymOtRf3P
6PaC5rt+xuLW2ZigR7E898/9EHjiQ/wtk+70QRaRrF+GqRNi9SwtTzzMujh4NI3W
GSpiHxJqgzRJENJJ8XaidA3zd710/Ubam5nr//I6wR7DnbEFuJVMWRopndCnszgD
K5rqpGnm5axMP0j5WLiGk5f4x8dL2iWmGvKaCWsBSMZ0bpgJ+ube4P7s0l6tuLb/
5rRnzXAPVv7GfVaFzawlm95YXb+CROuVvmmsagl5MpXJq6JnQqXcBcvED9kuKJfd
4GoSSu+iOIIKqKW8hVwqsFFgmwYbIk2aKBUtXiUtLoD4JBq+OsbrUzgyw7dWdcLB
avJi1ZUWi0XETrQ//vYquqrc85poSPPfMoej7Bt7TY/hrYkrTf5PDAoipxnYCB81
szNS78wt8M7kD+bVuMLM+Vmo55dQkkIF0vg6YSFwYr5PuhLVwmgX9hvcuClzMoNP
KGxkvXGdBFMbHyH80zN9q1/PADYgmp+ZOmPhP+CeQGl3UFH0GQlSD9PJVwTrKZBf
INB6XsWEuamGDBW4RVpLqt0bxNMRJvCul4fu0+wnemNCoCFRXxwW+ClaGmHjywpf
4FeKWZX+LgbUQK7kTFCr+NOpVKfgez0YJKzF3PVgRvyKIzYgS8l1xZK2zUxMpXpT
g1TEaZmweUxojj/RNYnSuxQb9TxgXHXheE07WrDaMAiNCLLomnuGucoTYM+QKofy
Q4WgrBOOKddCA6X4mvHI4sUZFCJhzDW74Cuoe9ZtUBEcZU55TP5uJ+EvyXdA88fU
0ZGPLBrB7+okmpq0ULtY0pu2BKvGaNWHq/1gF9uxpO8fKZnZV+9JlQ9kuRD+yIC0
h0juP+XCk4WTejnyO6cQiJXl0FporCMHzL++17R8A3kwRLU6BwBTBpvttNJR3orp
RKIz4aQrFnHplsNqB9Fx9Iey1L1wZhr4NZktGVQzwCbktymfXGoLhtiwztVib8R2
6GvIv73jFHBBroMsZXslg2xPBgPYgPDLcSOPNwUwwBf8IjAWLY+GV9zL9nuWgTOT
QpNcP319LW9iHNA5pApo8h636PYz0LrGAfvWRSZjdoXvcHS0g0j2qXNFPFMkM791
ul5cA2SMkSfeOVN7TGlsqBfAg4W2lRoUy+pexIOosuk8mcpFeYSoDpvygE/dTPtN
Mzhc6aNWAM9/+dxdrCzEJMLPBMrJaSNYC7/2ddCKNYVmJRK3zdAL7l5Toyqd16f3
KiJYTv+kylT5ljWQlzpdeuBuZSgknczhzuCiZ3TMDpHHkPAMwsrJ2+KNQVoQ5e0I
fOg2vTSMgw61lBx8WhK1QYxdp13avQAuW8jJKz17csI/4T4nRmgpNGWTOsQH/x0D
7fvHfuvveSthAEWU2ErjFDfgJ2PIpFoP3Bi7eD2JFQD8h1cmRRm1O38bREfACZWX
fMv3kz3DrN41a8EiIOOf6HIv/pa+LFkXDH3bfeung6eOUZKoCxlAjFNg86wxvSer
7zgrtVzscC37JjUQdDXEb5SL9/8R1s6Q6FvW7LYS7xNkAdNwgx5c7cIWrB9BqAVV
BS24NO/ikWVe7pwTx67Ay9sUp+IS+5tRTuGanQ7o7KDxpce9Xu5AGd6JvdGDt1Lx
SzJdPJE6T30fBUQkJ0rGzCDFRt5MkStGx2p3+aPd/xsTbEkSNqECtHHQnrS1MKhH
J6cBSP5fkudL1AVqRVwozQ5xTldXaeLAjA1GifZUioxXDCfupDglXMhMR0AhXhda
Mx1AOUfrTC/jd6+BnfPU6SNt6WHEtG7HQ/DxCcGav9E6GN7iqNLwom3aH4HYEb8w
bJ3HGoo/mi1ySlDcdP3MHveesGHebOCxtiCidDJ/OAhtnurQJBnK8HcINuV22T/B
xDieCP52RRWcIkYWmvMcSuyyYMCqu39CWPWI4lJLi6f49XHdP7RBai9mMO+RD4Ol
Cd8aiwyPor7erjPLWmMOs8fFEIDZJFt9LniHx2+jwy0Xf9rryicnC6sLFktYtQtG
dopH1reFec/qYzMFo3razoERUlZfgUbwNyCYC7ucZ7ZK/qM8ZYfhZqh5wym6E3Lv
dwhXboapmm4ULK9CVKdQflfB/Q9HakFy0mga/j1OFC3LXn9wEQNz5aqygelYegg9
zrYjNyv5H0n4fRp92QOszdSeXg8I5+rhDYp0Wft9I5NOQpHvsSfYtcBDWOvfDbA0
deM16gWnQSFKbbkjb2Fd0VC9MUldEjYjCt3vQ7aicLGJ/bexEjr0gC0NwCR7tf+M
BJlBgayZxgLakxB6c41CxEZn3psI0ajDRfo/zRQ52PxHlr9TIqnRQz6dMUBp/l8W
UxgE3BPA6y8vL5aqhuu64UIL6pJuvIfTwcBs8wxUyJP+vYEJsVExsnUb67u2iXfo
bLcXBuLYAhFq3Z8ZSmcphICbJc7tqkfjLN55pkoYItm875qzJ5HQi8hTp3xqd30e
BWLAheGCN/o5rIoor/fQdiFxSxMVnouyP1MNP9d2GYO1BOT8/hudUNW6D62Rh3ia
ttV/Du/Ujuz23JZGegHVsalrxHOi8zXH2lYJDvWUd9LYWbb6Vm+ZHktbVdboPfa9
/L0ubBQgFORU3NG8tF6zY87iCWNh8OSmRg6TdICD/VS3o5csg/oc5ErjVI9lcSCq
3MEF0CJ6r8kcaXoNnMvYFVn2ejU2rz77UhP/GYF5Z8dZB8d9KM2diNkpCOBnQg9b
3IfpBlFxN6evcJ9rIkzJz+oa5N8d5jqn1RAgy6Pz69QSVI9Btc5rPGBP1+l9H0z7
pCf/H5YSQWoRjqDvRCfdsP0jVjBu0WqXBlK6eaOKnIB9kZt2oTgTgoOjAH6KUAID
znU96ISmnNsAOsTfX4MTHxfNmxOL9d3+izmedKYahVuwHhe9jiNFZB2KxqeFnJiL
AiEg1zNU7S2WlTgsYZ0lyfzNaxqkzqjwHqPbiZH/OOqPCLiTEkpWBgxDUH7a6vEh
jjOlRjp+ipN/CjsakgRDIfU49g1mVPIqWIYo4G+oE9UZDeR+AELq1BsxsTM6dKxB
UOjdy3PRiIJL0Ufr7176q9FfvAh9A9RcbZ/ZqMefhs7dpRc8u6ORx0h3TsrplIUw
69wPHKbQHfgE6QGkm10gIxgPhEtA0JJ2A2A9wZfax1j6t4ZXhi7S9g5tTM0wK4Ir
k30QJQqVZ1+121qU68ZNQhRXBRi/Xtqt1eO7UwlY7YsOldPDgqAWYp32RW0TrQ4x
Sw9O6X59Ni0Skg2fe48D5qgXfo9fSZrDyxzkrg+/a/oxrcBeGAiTifVsIyB4Sh/4
YctBu7o8Sr4kbOBe7gECtsIjiEu5utbrZ8cFwAGoHigTa/HhlyJaYJFqh5mHZzFv
zv2fc0nE3zgSbAklR18qN6toY2qFd9UNIiHyH9ACoeBDh+7d+EeT6T70SugD8BCf
APHUeiTGvDrDNCKs4+GGlnc/n4VaO472UmHWeVo52l2d5oQNwyZhoH9Ytcorn0ED
gcBJE69eqeT9vQQrQ9AjRUPTMgn1byUHb7ZZyzy64OLQ/nNKWwqITy9sYA9QTAOi
eicLR9uZ0Y3ufs46tBdRZcJTnty+FRrLjHk5EYv+9ltLrSy/tPn3Ahhi4uXM1n2+
rqTVan+u3fwYRP1xC6QcPkyXUPSmL0gx5WSgb8rNkcNSq4PZMIYml0wyf8XNgPgd
0d4bT72aVuKFNTX01ylmn51Bpo4LA0nXweQd/RVIjO7h3cjhDQoY2bZFd6fGrxjl
G0gt6sUr+y9K1JqmoHYipa1P1ZSREoBnv33mNaUm79CJuwUlSOFYed4obM6zoX4M
ej0W7smSIur1RQ6PP1lCWtEbZmkLAh0u1zBfYDCkY+OZLCPj4/lIe92eja+kLFDP
5AbnRWCC4ViBurFdBKCauI41rZWxb5p+ucqo81C87lx0rnNCS3fEvrz/pom8FrjL
ibSWsIBV65aiJtXM/jWG3OlGK6mSLPsoYjFcEQDU5MfgMtYouo3QeUZXSpZnWP2r
uGIL10aCAHjSAWpyYV0MLXre70PpIIgiSDzgOvm00OCRkTHvuoVqEUC/RzMmg7OW
oe7pBLATRAXknAgdLrG7rRLYCLAUskArSUOLQbASIqUhNsHGoEv+ZlIM6zl/sbHO
yt+etU/h2TF6X8AH6rd3LrPU4zc21C3xTv4NJ/ys62i7ib8bUXtqAgQxirQ2xboF
DhRI/+TpMmtwoGgXMpua1urQ8E+sgZ1j9ZIojwKLYycGYYXB748SyrXa36IFudB5
PBUBU9BfbdbDrqw5Ut5Ktg407sV+UmjyiExiP+Zztff4OUhoB8586ZVUnqzDrueN
UsdUQejqMeldXOx8spivC0cUzVak+DRRjwlxQ0c36UDuGCiL6u+8zRDVtpTdviGc
XGM1zAg6Kp3gkkjnO+FkdkeSCLK5UwpAUqS4edTv5p2QTynvzUoLrUEg7igQXAmE
v2gNAIr/dr8JaSjeY0chU6xyueuhxlVnfkLd8g8QHQrZlcCnqh/7UHZl+nq137as
2e8OFoF9zguerBef3ouvF42spD/M1VZxv2fXrovSWPoFoaEhb2kKtc1yw2tDFv1q
fUVSrisfiUa/W8u1MW5HTJyuzoKL0p0nsbgLW0VI0tpiF2TGXlSI5BgAdJdFqB2S
1d9GuM4Gf2ar5BHStMxX20BU632NX90Ps08zBxp+w7bUKX3jcgY/4ZToMmv5G2gT
hEj0ey8NWnyrS7koBlUa7x+1HeKy0gExAxBT/3wcpPzk71WPB2/AjmVoWG0sJ3u7
9c0ARejfc8NAmhVKTeUI5f8hDIYsQDh+R71Mzya3BAgd7qz4RPUYxe6MUjvusUSC
5fhr8zo3MUadfnbnSVLTahQ6EDQpiI0SxtUKEy+C+nt1zTFUnu6P2KTSEvQcU0l0
8GCIl/PvLu/6qiIAOxQdO8wK4Z6Nm9a3SfGID9bVKNAW+3COAzs7CarTpp4MshF7
9FWWIPp5fsvsm/YERA/zM2USgD2R/tIaFaEEUPjMVG836ILem1y/y09hBNDP+dSx
5EVpr2yjp1KxOueghgw3J1BEu6cVQASRR9IgT6FPjHzOvZwmsP9MKbutYKHaGPwd
460wdHYFWNe2U71vvKjwMSTqTCCUni7dwWzw38XgZECLAQPzykTGVuhVJ8F8/squ
9qHbGyznTQH9ULFkKXKpzai1H54cPAK10PHiEHEiHNxNPw9vBB4Df5WujRS/CarK
Br67P2tTi6o4sJS9EQe7yH37BUWlz+uKODBgYjcAGAk39bra0+wkOV5Xo1NrHBEp
oGuQUwZJsFjsx2wzvKi3qJMVgT4J+irZh8zoFbkNNQ2qkBUA23rXjUzlzdagZb3g
xDQMMLVe24RHau9CMw2Bc59OznELQRchMZPM5uCsnXJRuZuDeTAlMYY1MhMQXJAp
65W7JTZPPd8dEZm8Q7maZToNR91ca4Tm07QDDpSO5kLkcF/7hp/RSsLNTQ5UELRC
5GL8Cpy5VfXsKjr41zhzrFPX4+nwAhImRcNJytyRppi3efrwCeUjVnoui6cMArfv
ZkR5YxWRxU8zGYdOA/mWK23OGAhsmFbixQL+TS3vwGIBmFO1hztnVbr4kQVKF4+L
gCSI2gaJSQGV0MzoPhiKGctxVh1HWwk2RfNG3FzVuXKPPnoadZUe2xI1auQU0jid
95VIUlKmQsrSNUo3oeduST2uz9Zo2Ryp14IbecW08t/YGJOuj+kJlY63/ycv9tNI
DTU1KPH5HpHNr9krbs8/Y9ETfSl3PycxrRh6cJcgLG8ExgOrxDDpVdTUWFrcL+Vl
HCE+9TeaDIdw3dkwdJVb/eKWmENaftRRwVDgcab9iGPKJ6eKU8csTdgYc+eiz/tf
aVLiiWria7xL2oDHq572HkLrjiNTAZD6Px4VeyP3VN/WYOJP31ydGgZejj8clQsK
lMzmZpOV/p4EXLagX8tz7/7B51vTMQ1mUwTr4cB5Lp8M6cUgGhFVn9JM3x5R+oxJ
H6EOr8pAW08Ngnis2K5sVA5q9pwRyF0A7aTBPiDRmM5DyQWTMvodwcuUN1pVSwt0
SIrouZ/LkaMxKlTa0Xvsi36c5R5/ZUJf51IkuSMr+4pf8BLuE9z7W4FOwWqcTqiI
JtGB4nbMK0EuEFfN8dN5/H8IRkLFMBbY+qvywAt4d3+/mMqJR8MGwp4/vRLF73ZC
vWWxrNJwu/0wd61Y/R9zwVEYOSIeQCyRcktp4FyS0iWkuIsTGfI/reS4ZiiInSlh
55qzhA27niZDwyiCM+ClHzjznSOkojuGPTEgKJ8Qlggwm6EAju3EO+o7yBaOxwob
KF1GLCcQygZ7Z37x1pOgggWRdwRYqQmc7WAUYsIxy7fT7NE8gknXzwcIgkZ5koob
y8M/eY9YK1DWxTqHmTUKXIbed5lPB9XzMr3rBTMhSYUte+OukI8v4V9Ao7ivFrKS
OJ/gfJxubhsYZUDib4TE2ju/fowHhPDOS1bPHs7umYHh4rtlvUbi43jVt7+HukdN
Jxyj4TqLNIlJBHAFxrE+gE2p+ryXXJ4TfMf36XRHehV1psZb3ZjrVbiKG/zyr+xp
zOQ4PnLQeARczcyofNfW/gIue32o0Zaw+cgfSwhO6J1JURTC3xweawvWAjz8a6Xw
i82+oN4B3HoxxNUePWVglIYWlCX3uk+WrcEflWm7bxddcAAX+cr0+c88c1y5jXRH
rIsCy+C4WB2vn+aL8nhs2VgcT9H1LfN0Z8kLgiJqo0btc4wU5cVffNT6wG/3xs9J
fGM9Et1649bcPydt0JTvhwNmZhMF+FupgivSvbc6/adxilP/ofaH9ykd6BaQWql8
JILNT+aMv8SzvMi9saFB7xV5pJbW0ExvG2r075ussApqgOsxdySBMaqWBEg3uPwD
n+RLMdsc1aJxn/MYUxi4ii54WfGWCJ2GsiBCv7dfnFttO9zbFDi47Dotg3F3IGaZ
SggLxEpcp90nyYyxJDHEASmnaNCHC/5ZDoWCl88MHkUUFG9VRqKBp/5KNHfF6iwf
ZIT32mB1yyYg6LbV6PBbUzX3GVS1gImQ5wYn94+c1fuVxelI0q8ARtbbX7Yn2IYm
lxSQ32aB0OHf8PDCshKDQX94k6kWZudyXbI21ibyZ0q4bkLEju5si1S4iU2H83r3
YMRzyM6tY0cPj7Vo6jIDGnPKurvZdysDPQMrvsWeZygIHz65u/KvYMasAwTx9ozV
Ce/EVjYL0ANT45ZQWhWfyLMgDl2gT51qoRQmCjI8zck1B8MSgZRNVrjvqDFiE9QR
qxPiJe4OIDnynbq//nGYCQUidD1N8971K67lX2D3IvCvtl4SLSC2qr749R8noA2g
3Ad5NLR398KBjWAvp6iPv0YI7o6UPS+5jWJT0Ryhn+vGz363Rcu1MT54lXpMexzp
Hj1/TVND2TB9egigsgfbn0SLjSC4CKnRpbVXcunR47TSsT0EKVBJI+S+Cz0sui4W
h29/w03w/46bTNLH+L8mLvEkzS3STdZwd+U/LaTChycO1xiDcTyAy6kI9BmZbMRB
ojbx+WeT5L0n2TOphVmjl7XVyCzI0WEWWw2dqs0p0Rs7roOlNTj5j6of1xtKsQE/
87Ttht1UnUri/v5cmKhaVjEqwz7YtstSdO93lT+SeLw65upBgeOium5GH45DyXX1
h2ZTdzpoFNUxyPK7tCG2uTrZUM23Qpk6r0F+gUKTbFuKbFC8BR7Om7EgIMw3CK7P
rNuwsQpxz/JYw63K+SGs78N982nfCHk3/HsrDGqcqkQEhppMpqCTyr6k7TBw9ZX3
kPCQblXlvT3b7yjUmaC2g89AB35ImTh3uXWFQhRgSrGWWkpgj51j6RAC06s5Rntn
NksjNKtLvL4RxNzGY+G3VmcDdozuS9lPJY+Nv2UlBXw8aQaIc46qh4R/LecaEib3
IPJOFg/64XDmUkOtKV5vNJ28vpEypfxaIAhZcyiDwsddZERQaQPBaIC6EtfBO+Rq
9zMv/+0jHYyirKiYtW7R9m9qCKeObEYI58YqSleBXXQiu75Vpxumq/wjUARJynGE
Ty+1UL5tJKUAI5eMfgnbXqPCkvIqM0Rs0yp0IHJKL98qF/FrmYik8PaAOJuI/mRP
texpue+42nkOCSZ79/OUHxSlCWXw6BfBR+jcOY78KY7A3oAPJHxIMYyzvYN0R1Mi
Px36gVSHgWtsirmaI6zF1tFeB/BlRXnWntBDPsoQySbr96MXClRFgJbl5nLe+7Pg
mw4Z25r1h4WYqgpjf/IWGMiOPlORiLpUloCvHSqpR5WPaZ6w5Xjnn/eg+oTpr1GP
VbIDO8B7H1qqGeodyOG1aw6w2NYodAZm0TLVhOSpSVIHlmKFwBXyv2MxVeB031xQ
C7UAHDB1XZWhBwOhbLPwD2jXa3+MjSazoGaoOAstwQ4yg/emHi02587SN08LIDCK
yadVGd5l5xyVfo0ICMFTSERmtgdL1VSlX6klzB0ztreoVq+QnUAXaB8H0lR8WOzq
PnOF3xaHN5Myg+6pHln8MjgcTPUpPEiZVzjLYSG+RiJKegcF4em8YQFPdegQo+9Y
z23gjJuaCD8O1u800D17bGMrjpiKAhWapvZjH0CpcoBI0H4l/5jyDbAHnMMT0JEh
0izqb38nMJBYkEhh1wplYZAeh98pGGnUkiY0AZe98Y46cqja2UM1lpdHU5v1B9Jp
13NSOcqEFVuY623q6yEV1TD3U3J8oIUexbiZzbzq4RWl0RsJxbYrGmyNeQK+JDSQ
JAcBaGBsnv6et6td10Y4xDTgf8L04J9GiO0x+49CjP2Sbrt01VqB+Db6LS/joOiO
RU3A2e0rs0aiqR5qKY0aUNNQ47t7e6pMUH2GaDq6LmUZ3BljZfA+zxTwV7KxXecX
/ki2WZ6bih7jvl+AnqzIxtSYZ4USMZCS70QAN145vibHIc7ElxdvxPeZInt3RcH9
rXC1W/d5cQzM4CQ1oK032zF0webo+2uE+B9JOHZH8FBhoBdxG8wf0V96k0bKMf3O
Wg/LPENxqNHOSic40nwe1nfIh/7c7CsmcCoMsfSzMe0r9wJjTJXtXuHX0qxagZMN
se3EawxPTylAvH9wjkEOT/JkI9ymZFOdA5KicfzuWNyzkk0vLKzi0WhrLMSGxkIf
45/nOlff6p80xw8MFmjNFG4I4FBZCfYWe9Nd6uOJ9+TjCiYVPshOmZs84+h/pTkh
fwEzyL6zE35L6lGcyuHbPiEwLpd85+PyLhNE/Q0YHNXNyICq+lNUOuJg8rpHebFI
Vwy8sm9rX36Sr8v7XOoI26VyBJ/JYGqN/rk2hbkjk/aO0lzbnHdr3xXbymqZS3M6
adTsCvqGbmV4t2gyspDpjkIxdPV5RVOPi6Jp4hrGiH2cNVovN8IxWk99xA/Z/HEm
gi51GGgZhc7mb7DY8oLQkbooGiICYBCGP9yo72XLnj6M/q/EjopzyE9aVO54gaPZ
S8UyyQdcKL3z1TCe3iSNDBkYmdASYwgOPpwuEq+n6zjKpxFfi1a+Bgej0Ky10vLy
MQZHykv4WZE58hz192k33ysPZJnlJ1UibqcFlLbIkbXraogckMqUSZ5gBN4Dl60P
/zbScsFa86s+PY7yGaMlblbtuHTbDdv6GYoiQwIRH7e/pmyLgilHWJvZm4ZAiE3O
5IOmm40KOQF0OwuOp8q9J1TgZGiW/pEpiuhykfVqM6u93QH6jNgwNOkSQW+8L8vs
v2RZJruc0IfBVbFGHPUbyet4+VBaIdsZqmVOfoamQrWHGNODt93X65H8oB7RArQQ
RxOREABWvDyCn6AOruQw8eE2dbKIx7qhbIeRLWnLmfvMZrJqPeYniXftquA3IF0R
WKO/ePGVXtk6IPNKBnaFnj8w4sJOCt5qw9QLx+REEsHLBxpXRBw+/V3YlUDlNK8B
iWVP2KjQkdOCcIaPAp2V7w7AWJfD6J0QOtrWrgR+w/jqot/GgtDmPgLqg+dkXtKC
eAcj2bTr/4i7VLS9YFxqJIu5zw2L5NXBbT8vXX6hMEno80mWLBTtI/EktzonOt4d
chw5+PmWl2sO5gCEQSfXnVqIvNnx9C9fAC5z4JxUUL6NGI/pg/I8iFd6QVC7wPUE
nXk8nTp2pV0pGD95IFquCTfF3XokldTwojkb1cRt/xt5gBR4ldvLpdRtxraljVEh
ItEcLrgsg6O4Yhg7Ja8EVX362TnOVPK2nTyXdmoW3mRI70tITu0yf/02TRHb2Xmn
LBUtwDVXXfLmgqg5Q4aS1nur/pHuMSAhTjfyYkFnRGP4Dw3kOsVottF0ffBayFnt
NUv8p2UtN6JA17ua/34lMLQp+YlkoSNbztPi/setJFUK0a/y8YxGGlwnTNeqKJWX
E14f6pOLSnxvHsrVtpltR2vfbFDgzTRPzgo/7poazVkvF1aB5Y6QXNupBVy7j4N1
YLkU0JU/C9D9/yqvspEI/Y9hpeZAvmUV9J9gbL9BFP5gvC6abbhmqWIDsj3rtFEh
SoM9rW2Tec6X1tYK1n10ldrNwrk+m2/8VoQm2IetMsOWNwCV/BH+3P8UXKuCQXXb
ktBlDOgFsOO7LdzT6//wqGiBRhA+3okbM60K3wCqBTe9OvQGhvo2bzOVwshp09DJ
fZG33g5WUMg189CYlBLwcbONdAAjiDO+qGqNOmlyWZTdBCQs20jRnnyyEAlOl4hL
U2qQavdxb2thei0akbaLfCC6d31HZOtNRQls7KpRcx2pTZFZTxOy7GVUzrGm/vYi
KaEjFL7r4RitSgLL1CJS+l3PyuQVR4eWZhm5rdyXjjgJJeBtt+UcNduScqZqK4ul
4MxywYZgVg8JsEOX/Y5AjzF5G9rQm7pZPzZLIPW1jU2khtUbOu01jE9KtbW9BCl3
59bPzDgRosiGjdcrVho0ocLBRYU24JHEynzcc28WasD0rnvkrVxigWazl0MEOR6d
veN+mkOaKvAJZGFL0sY6C6SkomF/1z1xp5C86r64pxy6Y1FLEMV80KxcULxUfnCD
9rRzxyXRxF0JRNgQEp8ktDuna41X3QBu+5f++xv+TnWfU91rkfhz1E6ULUBYbf/a
3ann3IxJNxnkLbWvhLTlZm5KCnbd+JlkcPhLIz7ZdONix81Smx+yemMSP2sSr9US
yWeGQML+Qqy8VBk53HaypBpdjaQHvSmKk27k+j/zoZbkK4OppXU3XWfU4+TtHz0/
xTXpF//2vtGVGoydl7GXeMTB4XwpgUODwf83eJGy3W246pDuNWgKrPSVj2z7WBG5
HQwKJH2h4FSJzEYUDNefzcbOah69Hs6q3pe7pxngzPLYBuDAkP4vsPD46pj6Br9N
D6ZgZgRGcbKPwm9eNAqTVsqykLtNtvCTWYTWGEV9hp/SjX9GY8ynnPGe5SHHI4xR
ijp4RfPfClDspxVeXMLl7XVUt/hu4VuDePXRSaF28+O44xY/nE+kaEa7X0Zqik9g
+yT7c7WcykN4DYzZvkRGzG8HjGCWK680uQhyO4l80bvQRqnEAxJbzc7h/r8VebW/
PIdGk2f6M9AjTVRX7p4f3eC4Yko4RR6Db1Rh/i3ct0S+M11dswqxRDjB69w24D3o
ZGbYlR29o4WJ/wJgiNvijE5NoeYVACO720sw3/9T/CG+15yF49uqekc26Skl7C3a
IhM7CcL3t1ZD6IfH2fFbOmtI9TD1xxou2U/ZBFp1H2gyZs5SEEUct1rSZEI71EC0
VLHKVw/CzlGKrVGZNyh5Sr4tGye++YT+Cb2IKE08EH4Q44+n7vIWvEX643Ry8cOG
VF0L1Q0UqTNk3xmdTK86aUTcUqypNxbSdFOCvrJ6I4VD+sv0DFBK666PIYc2+THf
rynDN4Lg8+6dk2UHWMf7BZ2TCMdAH+u+vUIKj4uT4Atz32af+2wIiZpu055XZ2rM
1UNUSzVa74frKn7vkEBO1vcHPxDU9ZPruMrUrfZC9sSuo4p5sgsp8DbGNnwDqiWQ
c40rp9Eq5xhWCF0+770q4O+Ufi+mXwyiY306ZWBhcuQSkyvZ8e6Qmc0qDaWNfMIM
u5WwvhjaOwNWfr9fSVWVJyd24AvcmulI04do0U6C3+xN7vDTS60S0dQIZbaRZ7Vn
y91mu0Seq8qf/vhTiWM1BvVWmYQ6AkXVH7FKf+8ANx43/vtBrwik/DjDhhwpvA2g
Oj6iMLEF10Ttwj1yi+l1BQgINAam5JcWL5SZ0x6jLw2ePAOYwuhHXtxHKarDCsj7
jcpuGBknN1dLEzJdFJ8UQRbmA1cXZmVVFSUiRGoHj8T7yyEEobPYRPeMGozMm6K3
tBmFh6J79+qSlWj68apSaSm9P5bpfYAj+WGN9zRVC6hI7TBFhfGVD0A+HlfT8W0t
OZ44bklPc4DVKXWI93HrTFImPRhdk/K1Y7ApPDwy8SHqya3DSMUolRjkepfkvc1c
57+WlQdtLuAxgiXM6BOwNDiaSHFYhps539K9bcZ/RCax6vGfPI7iCiwkT1OenOPI
seixL9d0GqywaG/OLdtczvKBO3q50qa8IrIVQZWC4JH+nE0203ji2sLg6sMM1IIs
Ais7/pjceU8QBskHrBAOoAr1wvXCmDQLfiTMOnpxbzu3LS5r7FKplSkrdsDF8ppL
TFTd+/URBYSKGK2z8LShc2wnG0OUIe6BOifh0ynxxqUEiWhiJkrd+FHdmrwoS9F+
SZnAsPrO4EjGWSkiytUX4/OsdrJYLi5I2GfWvWLUlbp/Wa/EcPmPRMsTXjZPkWKv
0Znv3UX6lKOxvuD+6Nf2cniOjg/rjqk2qoKaHkM7YAN23KePjRY8fDCu5m0mAz+D
ttIpsssxboH6hHEvjlttrtb6pWnkFXNY+ILyub8rEQtBjfqz+zNsTbRhTGP7KFok
TpOzv4oc0YJYGmMoiOrQCJVqrCj+RFq3C/UDv8k0E1Jx5AaEF8nVbhJDM/+qv34g
VjRRU2OzmsCHzNaV0D/VGG+uP0pRTWxJ7D9CxAVIHcK8ffQR2nBAL73YZl83D6rJ
HA22QtewVfLmBkWKYhW6HuSe/hZECRqCxn3ZJLGxrM0o3oCjQv6nvLmg8n5haIgX
W1SwUfrq04caRghfnl/1NzWIEyE5HQ1yMx9JxlHGT/OV+iknOtZ73ZFczoccN54E
seCuo/IrudIRivql+BvDc+ruJGopbKIZH0k1MbBDvDlGa1csCkj687wJKLDJWLVQ
VY/ecVB5wRVaSKYgyQA70eyoSY5C06YUnmcEliEhQqk5xVg78yP2incRWL9hSNCh
v93VX1wODdTNrRuHPY8xvYiM+be1hkk65SYG4ob788GZX8dKKFjBXp+ccKltmbGQ
Y8wWxbUIkWT5yrDf4Lbctxh6RRHpD1RebQQ+5D+NPYl9q0WNs3aglvfqCQrBViu1
BAk7JL4e5BBQSEEimr/H3W1fZQVsz8L2GOBipP7RciISDI7fLqRMejHlOQ2wdX9Z
VAusLjkMm0H7IPJDmFG4J3lVtlFBgSGuD+9lUrluswF/AYTbZGGojj1MSwDV1tLS
06JGhn4wwj3WinFUNYx60t7KSQJvO05Sex+CD1iBarTHmHSRoGmGqM3Wd80gklvx
cpA8f29WAn3XdS+dnwzW5ZZ1o7KNi2KLKDKxWKGYbHBZD5Q7d4MtwKaY16IPo845
6IMqcIA+nOfuiQpNyjlCa6RGX7p2lkMp8CVgb4S96zu9Km/9dyXEU025Rns7aL6M
RFLQTxLnR0Kq+HM5o8kmAHD/bTHGJvBTU9SUhQB9/ab3zZIunsiZqhswzZi3YWla
OTy21p0OLhRaJRSLPgVAQZfB5RtIGu9ekWdAsrHyMPGaVMWW+Er+xn5SUnPFOkJg
xyON1ujNSDgsv1q3kkfTVwRZrK+AgML1m/V6ucuz3zC9RyCtLGhoNfY1rNxev+vF
7Odz02hXaidgPgijdleQF8Q7RRXva5nyuoptbIOhpKR5l9we0pIuSsb84ElmBslD
9QpHe/EQS8VBRlUHGdY+DmZ7MEoye6t4QQtUVm2SfMkYWQS6JeGXsy4qCO3b5JgI
4XagQugd0lFUryshq1fGCEwqlLEcsdncmTdEOEjsoLtcndYSOCse9QdkaRA/4Naf
fzFavhiN4a7Y6/hG/b3dMM3b+IbTaHF/s3gYo3FCAd/GrfbbybxVcTyyGkXjC/Q9
kaDC7KSSwW7V3/B4VNcQdpplSbrlMR4f4A+hA3aYhR1ldG9wpFU2VRjK2MJRP3Xb
IuvdHvoauQo+b3n6Q+kgWZWejuBKpwpYIEesTDbJXdjhCO3Lu+GNu26JoOEHUGBc
a+DVZurbLX+dUe8qJje8vTMNtIwF+y9/4nZduEyAlxW4rLNwey6MbhTf4PIifR7N
eTAu73e6uJTQhZ1QDcdNTlQ5mtEKQprxIY75oJr2/TzkcJAe0jJGeWejhCMjtzUa
S5elTlgi+Ycrvco3QRGMORBHD3THPokYDy4vXmea1y5tDfkmluCaVAYy2LHY6yWU
ygCrjOMFc9EUoNeSlk/H2qs3ZJThd/TCV9ZCiB3D5EObMBhcq/xwH6TPSwK/h5g1
s+vhLWLynoqcHCSuZYSa1G58SAHPhyaJnllxf6VCKgBA7dQtejP3j846b1qqSOff
1RvuztEkTPfYNgYCm2lMw2l5qde5BTdEjg5sYu4zNWJ9SxrOKUO9kDtBYZm9xtKJ
WdaS3Fs8Fh0xijbVRz8FC2vsDNWKAFiqUVcxpwo+NJ7l/IOAOVnzZ62QVfFHogUy
P3rJMN+QrrSUGFPVxwBBsELUfMfv/RE7cZmKSFE2BjJbwKsTOCEAodi/41H1WWWb
XujVCUog8u7IWRFbZTjQiT+EUY4NDthFq63mfTTTZdGcB0At7ZnSukHv0v5qah3W
Sc2oogrL1lQH/wbgGBW4+78mFtseRZg3AE9pJWidSVLm8qsXmZNigkOS9UWyA1kx
LVCEe6He6vDvhM6vrySHbrfEa6GZM4y4nZymP/CirKWMOZTsiY5beRwXaz9vzzcJ
cTF7kntpn5jvwQbe5LFbhsQtsukkdYoE2WcDYHpxHLVwtZPE5MWSoSDQE8q7IaVH
6Cm5sCZ6ldf3NCGkNuLm1ahTlYw01ULGy5h6aIxFvMLvmw40Eq6TiUzGHxaxfnSL
1jFuNDdak/B3gNMHcMCDrLbYxf3oricmX3u46v73f7B5k+8wj6nBZ90LvM5x2BMv
2xlkN5N0JTyfYDYsux1dJ2HuV6D2yrYYMlpAjksFHzg4O2Fhj/iTHYp3RyiXpILz
RgDSlJMGPVcMZOajV4GIwKLJ8P21E2nuqIHe6CTriNb137s79y/hu5fFUAfSEqDx
x/UG48lM+sIZQhRkurmVa7TifZ8rgcSUN7KcDk/KMP1hgIj1NxlRTiqd8jrOBNQH
yzE4/Asxkm1kLzKxzN0395nZnLGmr4BySzb9L/819MRduTZswXbbo8sdITQ0lcIe
TGbbDbS70MByux8RDcXbcWSkDBicMb5Kra/yRjsAB7uOnehTMj1Vphz4Vw0TDUAr
gKoRVpPzx41JKl7cLsUFIKWD/6Kv9kSEjMKbYeCxgxV6ydgjP4KpThAlA1XEuwMd
YHVs9I0kRPejHtpVfj6+j+GMmGMNR3XYYfD4kjlXqI5d2TL/9OEQ2BfAAdf69TiW
xLU5aSmD/gDUUsoN096ES9aLmM0syAMeii3V1kKHEgaXI3dq9uB14TNyMHQhHkjR
v6sDdJEE1PaRNK8QSYr+1aFkWKKDgxwmp6U74pcanXljnN8Byf94eLgNFhf9LBd2
r79omoocCib8I/g1qDG/Hk+YPIC3eD0YXq7ns8XgHtAo6np7uZr6aP9BByZvs4zD
02x2VkyRtA/qemJ4/iE5478G69viGZ6nhzf0YiwFHcKz/dmcX6x5B7+MUap1nCHJ
h9P/Mm/ZL98UAETTyW3n93PU1MoMO/HjqBZsuzz0dLpt29ca+muqLlOwd0MjfuF7
3T3ysrKTmzjVlw4jO3Nor09dZVlxAMe6Lq+5F7raTA3Sw07XfNOGSOf0KWdqlcia
4EWs42BvB/UGud2OvvJ5mhwyfVrn0vtKDuRFZ+hMEH7kcMsI2s1M/2AFeF7JgOQu
SXpDyNhSHOidclc+vFmBY6hrycQD6cD7+wzHjOM6+b1LDjt7j1RwpsDrHLOiSas5
R5swDdPBKkR0HRyhiNE9iscHgvR+aFx9cbMWpByIT69BLRP41uCgGffd6Ov91Deu
LN2pH6poDa70Z5JAatlisnluWAlBPHXSO//kZgCv7mey+YO8BFi9Rrk560NhmoSm
aLxIW640QM6ORR7Aqsk0sxQhi0DCXuVC1DR68QaEHHD/VwnawBy5hr+j7F6EjGQV
S1YPNkhm59eme5kiWjAO7CHy/kObEaiHkLL/C+joWnG07sGdfqX21ffnpFdWdWB1
ROzdyWoAlpdsM2a938wfESN2PHm3pYsGqdLxfi7Rw/yzQhFM2fGKxzTavDwVhbM8
oGAhGGmjUfnGeIWdjQzBUDJFtZbSFIEcaT6mR7uvGae7zbJ6DHDxp/9i2a4Adm1y
lepfu/uZz4rCI1lYTwN/tpVW4IljbSoSXGmvN2QV7J6LsKNnzv85PA/thjn8+K/k
gM1WBVC2NCQoXHnV3Qf7GNjVBcvF42Jou4MlAel8F1MQL4yAFrjztdEcVq1ztg8p
yrrnR/rtltFedLBQYnLbsJFN7dBij1CzGYkks/Wz8jZXtGj6g85KQLcAaTGd/tMH
AHJCadIPOyeVMqubyRWG3lGVnVl/0M5Zvc+a8UwtHI1WuxItKE47CkcqhWYlnUev
tbdSx0j9wpZmlhZZawHMBwHXmgx3rYCqY3LRjr1xbVbX6Zp4dDH5tVRSAIaICNci
5+LcoDbWBkJyhmioymATVP3tKPla2HmEOPp4CM8nsxwRAEFIk9OixXILfapUCKdt
peE9TovJbhs2zyK7MOsSiA6CCPXvyruN2WxI0bHHlcUqHa/eYhTqZoZ9xfvo2X8l
QJU2I6yxKSc0H7zPpYjirLXGToOP9/qLQcFw27di7F71i1rj/dLcopctroF+LWlx
UQeUWMT9x32LzQIsExvq3BvrxXv+4dUVm/0ktfBvntclxi4ECgkdiV2Mw//pW/8e
HKyzvkBzucUfgKUWtZ/XjWAEPh50UYyYtu7+eQY8L+CE+27WY0mcLFZTXPJm0YfI
22SKG/Q2PxdgAgcV0W5OIMTM676sFos/MWBXsrJV6BUVIvccMynmTJAzVy6KC1kk
5KTCZyaBw6fKVyxViCx6YB0og6cEpg6VhjUq+dMhoiGrXUl8lHQPaXUNsJ81yubC
BPvl2hO2buAtOGOf95Qwyr8WaQO98q09crYsnk0zq66lZdnNYdnQ+ksqiQQFIMSj
ejJTm3I7/YlfekPVmjZOfnxZ89tRxAUK+gcDj7weYAu6YHxnYqIb2H4myRLPsWcr
cc/KEQVroTDYe9MUgd2vQn2rp2/3NEgPFtH8txXBqaA2OHDOOAQ1AGWXGSyznw62
OFw4SFRIRx3DzJcp6kEVCOgids2wcDba2fF5M5QYjSgGI31zmasgWL9a2050T5IH
bXxHR2hbGnlNCgxqOLANfTkJZkoHYOpKCSKfXItF8St8vwgQ1qp85tjQf7PXc183
kvnMzcJkHc9+uCLIxko0LKalKhg/XBCK+RwfiGb3/rmWOzUnvgB28f/zO6gSTwwQ
i4rMqsz3W1Otpsv4PwDpPXq+FMLnnNRNS/frF64+xhhB5YrJwSBrZyzkfTJkkMOK
wizWhRKu7etH9qSwTZXv3Zk7JCfulQqruFo9MOnPEEqhZSQt5vasUNjFjx8bQDNm
RUmJbNvlTyyrE46OwyY3rrLYAqI06M2iIhVY0Sz15Lpr7vnyd+egaf1++NpPxcYD
aHCYDnYDfyRHOGw3t9Sf9dnoQ3MJv7YjXnDw/yTCs6Em6hT8jlJFB3Ba9dpgsimZ
ACiOCO6JbMlprDCWMcKoOOeU/VRYdZb7aAkXTNS0T8R8lpkpMs0wxrkO4tCLHCHv
dwqvBVCbSUgBhav2W9iGLF6WVBhPZJqt4E2SzWLrBgiabSOhsrNpb+t/TbcEdvu7
LPEIBHqftSJZcrX7qJbwmzvaozSAyC3YWUHSNwVux+wsbp+tSb0/VBFfCl8Y92LC
9XnclYMhUFA1zAdvwt+jcQpGl99Qdij4+BUZDEhhMRqwSzaQr7wDxTFffH2pmeTf
QvAEuWN88M8Qx3Fr3OGiiZvepJdR/G5OvhT0/u6zQHG7Mbek6pzPgTuOVUCzUVXa
LdDPi57JF1UCxYr1UhPlARe0vwyI3+Xn6hLHwWI9RZY8w8y4Z+AMyH6T1NRgHFc9
dKC5BuA2GFdW/PVRTiWurwe5h6S1w1kkXzKj6NRDZFtZNNoiKsLHX4+1r74Cqu2i
0paD69kJQ9XcikzR/cw6hw2neq3sr8Xne0nA3SneYpxAUGe5XDQ79LHM42w/aYEh
cfgiJiQ/OVAOpOS6X383VKWyv3mY8qn9k6to5m09dzcZSq1P8cfMIMDRNBpO8MMn
aI6slHZtfr5cRparylgMpyX5x1vDuQ8GMUjHXYwDBjL5n9Ma7btqGtjykjfaZOd5
lQrdjkyo9FG40RBNv2wB10MvN6lu1upqYx42Y474T5WSmiFi8Xt+TNUY6uzS+zFn
6iwEHnp99CzdIMRbbYopglpvt6IbGWJ9yvCJ6003CZQsf0BxUIj1h+LwUL4C3tpV
vxrI1i9OduinX1A6RE0C9/U9voLaGBCRLcbLH8dMB9DBBECwtMlAyK9x8+sv8kh+
vpeX0YQho/trUy8LmuvmBeSNpVW6F5+NM1/PH6UpcSHyOfLUqLS6aMZTAFNeEwqN
wvDzSbgT6GuOrMnWtxQ4zDtBWtiMtT/XeQxnrhCu4nc59sFRxeqFVIL4L/+9s3v1
l1R8xW/Dt+ZcA5MfjNG3AAmV07sJ/C74F9im6NQBII+z/5nWaZ0jD+49hhOkbrii
Cy91wSmjn6rk3cJyKGKQURNraKr2x7Mv/tfrY3PutX+Jtj0j3s1iJmw9AYdHFGlI
6x+DCYJDzJe2ElyCjHMa1W2EIYwDkIYE8jTRRRSDQ7xxMn8BsisIZD0ST1ELjkaU
T4OGH0rhsufJmswMitXX+j5mxFNg2IyJC/eNLypPfFuQnG0+7rsKrkDUeA41pbzn
4ckKVwkwE8TsiA3drC+M5AEWkh/IqDrmL/CYVtO9Oz4x2YVI/wIQkOqLFjxGlj/r
c0pjXo6QXbeLuH3OO0RM+lCEaPvZ3EAv96MUw38T78CVNb8N14SHoqVg1pxXjqfl
CWhcU5dwwC8iCbtsmLgCqEts1R9WJ4YfAOE5hwpD+08Y1rJhXyPeR69LiMgB75bW
3jMQRJ1ovc6/mIKtNNwVumuQ/hSaxFA0ouXr2i8i1k16NmaJHPDe6EZnE7sEMl3d
E92YPXaJzRnlJcCAjqdHbWqSJWELO+WetJZabjdt4Bx3mancjeNqVhmt/g8k7pqP
tuw9CjoaVxFnozdYhw2b3xpb2l+uEO3REt3WSqlAlbeSxJyntdasDbc3zZAwnZVA
ne2kCVloRuW+LtVsivy1FL2J4mTdJA5lubjfuTEF/KxL2SSyj9gfP4p69vM8OJFW
GVDqnuMI0ACfBaA8VkBRqjQCFtcpmtTCnsyKY+HVp7GrNwNOQUvV19ZM+MBE2J24
2UKhfOGKmbfyYmKbSdv+OqiLUmZq22ziyBeqvUmoJRovHi/nt30MIdaKv3xyApKi
O1J8KfZDkTLu4RypldJOTpJj17+ZeCT1Be2zuJVPywLP8VK26x9KVNOQSPhlSulA
GcUwJJEf2zUt7kSoh6LSDekm05y8z+epG7uk96jC2E26qwvF4hff2OY3kfeG4zaV
GQODX9jtPt9KAblpYxrnpFpEVvoGN1jqBonKVoRWmNuXvC6uzXL6XL2vSN+koYb0
Xuyk8rDiRODs3iFx75ifhx/gfekmEIEjrDeBVsD9yOz2yCdXvWNHI8l5S8+UFvZX
8lzvyiKYNrzO+SzsEVHfpzuuG5V9PXdg+3LkghHchvwopBiZa1GkSHon6QK4MMQq
45Eg3LJQx916KJh81Kfp+oCyVA/oLyFkA/QvHwNuXEIrEv8Jk28t4g32dCJhYXhg
K0oTPI8XuVtppSGNDhD65i7MEsyFGasK0ySW6cdZFqxffuWmeSLUr5Kj9AhHioaL
wrQdvU1G+A9qXijaRLTYkMjafjLbceP8tQsh4zUlKmCpyfzksjTqFoAWfUmMHf57
IoW2EdYWAFbT5PtglhEJkFfLh1OdiKTVsXNCciMvhjKrUNzUA4LRcuDPEh08csu6
+LYOz/+psebPncHZX7DHt1smSI1M3lhjxAjNZHnMBQZ2kAUufRa31vJXWTkKql3n
hQoFyuvx1jf/RftQtFbtU9vUneIXou0/H9Q+CsoLQKhYEXGbgwf/8Ty8sJpHk/6t
i0/q51xcuHnjbqTXLr9jfyAlDANWP9g8R16+j96adg7hzO8xJ6X3n1R9z2KbNZNg
1XlZjAAIo3B0Bm5W7WphANfy3JLoYCd6ZX6oc4mO1coKTA3v+jxY86HXg0rYrpuY
gqEisCwrYVfj4FJ7CNgBVvinsjTRcYMHiAmA66YeiHJvRgLl0KuQcdM915X4KzpA
Ee/6fks3axuvhZCnw3Mu/pn7aSWJWNu+6mRWllFAfYOJEZdjD4FjZF79BN6QmIFl
Eg7umOnWnYhIcwqXitYbh812XdjNrIYLhGl+ZdhqSqlxGYuBvwgXHouOoRS8d+ou
wIkPXK0O4gcnrnBdiLNjhu/KkohPwWme8XC6MugN1vb76h98OGX7u/Eg3nCTCT/+
5Mqddyd5ebt9KXRIpvtqdogJTEg/c6Jw5uH6FSLK3rUgQhnBlpGpRAB8LOjnLqSu
0CeMFQrC0Woj7hMVameWiyNQiX6ctGlUshRDqPcbq8aiTZhwf3/gDJ0F5nPMH0oa
BQFob6ygnLNqpVyYn1/Ank7bAwY23SEWousURs8OmMdT9D4qGeWEqTfLlbmBo0Ld
uaItnuwavcmwg60yhjQAAtaRYCoAdcXN/BQDwP2rhChXK2Q9EUwu/IWZCL0LzhVO
2wShc05yU4GviVemgKE0aQmVG/q+Q/I/njkJb2Ubr3+1C2kOolKmAa7tfAZ5ctLe
KgW4ZpsCjCsUr1IgqChThuJncnRW7raQqiJIpYy6NzeUTKNzdZ3GPF4U5/rjsG/j
GwrBvQXqop7JSzFM0unKe7UsnSe9ZhX8zbpEXQ90IjnbHghyhMlYzrNofHL+iBat
TyZ7/ekNJBxv9zg3jtPNcLxR0KA053+ba8MqB/kdJnvmutecW7EdWUQA1FEkm3b+
LTuMzA08scb6hmNHc0Ele6JTrM2Td0mM2kfCA2geR4LFj7W5UnL7aXn6KYdIi9OH
x1UEeEHappEavcPlvv8+7HMhFvFuZsy5BLvRwTwpHR9+dtGEGpN8TmheK/xCtoMQ
QvRNjMQsQFDpo7G3MCNTxH+EU3nb069Y/B+xzMLwm2TW8LcMsrfrFAbqczr8r4JG
QZy6u29WoHm+DY3nl+HUuHQgf4IchkpADfb3TbCxIc3OyAaT1l4/Q/DgnIb0G1jH
06mdzEfqFfMQ+907A7T2OnWbziP4eCLghlU6JC0yaWvHuyC/f/1SZJbHQ4ZX6hXt
n2+gQcUz6m0uZH1aguJyXC/Y1S0wDyYUY1N7ovHcJn08OiVZF6YLT+ad78yhzU7S
JqYXZljVP4C3EaJHFFoZde5vW6vucRys+itAOPx4xY1KUdI/RIzVaPLrFe90XZPW
oDFELWj7sg9wLXeRwB9KKct6XAQh+iLPJUxVMc0NRVw9k+Zjr21Zf7CT4Qw+iYJF
tLIE0IkfUAPKVR3M6WnsT2YTwwRPtl1Ufjs8ERT9v33c6xlU1BWenHTPt20Vc+R5
2g5Ip/fsxfaJydzeJamgr58Ft7bRqF5Hx9dt7NLgYClkXGIE4vh6ZhGDlE7LGzRP
WoLYfcmb51vAv4BgcZlC0LT/9xwEijZ8KAIsszT9rmMtfuCDm00ldwZG8PuZ4TOT
+Y4cW+QLnTHoRNHIenruk4wsZ1oLiBZUB7ZL83LHyjB2aDGjOGMIp7TQnJ9dc/zC
7zNnKqLmfi+0BD3exGay04+8I5rlzUHY46R5z5NS7EkwFRwbvxGfyohUKW2yymnD
B8Yf6Vok2T3V8LQon8rn2A+q8lODcZDJzzhaha14gdr5jCcV+8fB0x+uce06cKMo
PHldO1tRi9E0K/JJxM2qVJLEdncopgZbAh5LX/acjHpJRRuGgrPdtR+mejJtjnuJ
ONB0bS3b6wC9NXn9mmShBczMHIM0b74Qwrnn28f4zUGGAdRBVvOgUA8FPVoME2j8
SASBpfRrf+wLwpdNzaGQi8RA225/za8JSf0USNMvCxzaR8Q4cv9CJnVQvgF9AHDJ
wwBmMsb2U1BP6EngotC/3/UQsKfblPnorn8Ize4ARtz67HaeKMHa6C5osftRVHvF
4SIhp8c06PYa2SPF5mQgnaeAaiWzve7R/iIERlB8GGCRtzqLz6nv50kyut3rHnBI
oaFc101RvJtKlESK+7YLnBxQWZ+GOxbju80F/TSmoitcSDUqaFj64u4+fl0hppYP
CD0y4Q4LGg2WphCe53uJnzozGQHXrH9YQdqadjGmkJsVj/Qze0clz/yOx54pr8Sp
c8W5M1ZlEucj5zEP4FsodG55ms71f3rYG85zVU2StgzCuSd1BWPtifEM9B7Knolm
kElj5H9rI0vVFFt4kSjJlWQVXXJ7+emLDz7eB5WFYgSbLK1UohpjxgcGm1ehCNPK
9+wrt1y5cfafnVRhmgqS+A0y5EIDrtsUc+3Qpc5EXu1LttaH/B4kUHpZswQPNl1s
4tpR1tSAzFcjfXQpHzlJb2eT9bW+UL8rfWyXPGaCHsHQWFD8B8TClnxsCSsFbd1A
ilfTuH6akj8qhJ9rcv5JAaZWiYiaXUhdYDDkx6Zd6Eg26dspyDHq8VQy6pOj/W3u
Jt8IJInvo7ThTj/9APbqSx0tyLNjDQy4jhg4esbZy2HhdPWTD/bRZZ14vH+kL7Qp
qaFbsCbxwRfj9ooW2lBee332TIZwKb7I+2bWnqlOpBqL89wv3u/aaCNnM+xuAYh5
ZryXo6rTVeiyl3U89N3kFAyxkRviIuolBiv4gKlTpPZkOQMSAtO2pkkp3kbGugn+
E5yimBNhJW/w14Lv7u69IS1W76IS8VkPcS2t9mJSTgEh06kvUlySnrEMbJhHpAVZ
8O9VzXwQrkCTw56M1DRZIQg3XpkmdmXQLQ9RJEOQ4xKHb5aM1ESAQZzqqSSLHbXF
y3GQrSTzsSwlscAiNylRAgh5jLaU3UxXgSdTCBHfNJqzau1F+xNqFog+fCWYaaDC
l5bnci0946xPCYiJGAuvAGDNWfkRzBHQoaMk5Behc+LagNlYE372PcDzt0LpuLWa
9kTfhAdKLvfosV8mtP5RtmKp4uXloV7DX+vc9LqqEg1F3jtBEF3sPydzoX2C9o6E
+Zh1asfGZ42smrAQgFew9OjnmlKd7rtJWwqPYxZP2NJcF4YNv2gdra/FgGrz6Oxz
2hc1YNvLGi91mNQhs4/Ef6uONx/e+ORCdYaYC7MfE/uh8D24gQwaRAkBitNXvEyY
goTXtDJKR5QQcSgQf8UVK2f0C+tlI8lmfKokOg7jzWLkuR/6Vu9SBQ4syEBKNlsD
H4izGLyKwwWgbBhOYpvtBb++wfuN+6h7tq0rWfTMQ8shV1em4aG+xhD5/WzJP0KA
SOlADs/sLGHUX7k/sEaAtf7WnQLSQXLuv6jpb4zd2LPqF0SCPM6IX3n5sVQQxVVT
0ED5pI8E362yBTOPOjprnE92++qCiHbcct99pu4M3c9sCRrDCoSYFO0Q2jxw4JNn
2pB8oRIudqIUD5gFjYY8NXPNiI8kJTr0cCasAfHhRtR2unRUgW6CfPaEcJMd3JBj
E+89NNbn6whFhr3yZrLlChOecsrWVKivgcq2i3AD77oMV92UczIRNmYB7eBxulh3
Zd3asmxK2STeUVZCGK3UkSwGBUgVg+70w4ZLJM7fXS0hRufoMQoLdfI1lKNshK7R
zdT4ni8Btl4U81Www2jsAJKMRvUU29HC1UecW4KpbEB5rAD5f0hjzYUkdBhw5mhP
bLJmY0oA3rR9yG8vGa7mS9OigzgiJodJ7uB6WHRJ+3Mj7JzkHAfMjqXyjrSnNENX
cqxhLPC62meMeW332dFkBRBhheseBN3teUpPTH930aZZUZ6HtMuE8FZK6+a7dPFe
mZjyfbkWZK/51MZEr+z3XV65hF1gqKFMV7wjKJCDW4XnsmH+u84qVd7QJcdC8uNi
9EQrhCvGGCChhCpBDhAOTDNIITANAf6E2xL2yX3ibm2OYhw1Jzq3iHa56Cy2yByC
OX3vZoIL4bpwOHEdyG0p3RdapSrgcloczGC+14lhnDABctYDqJe5Izj7JdUn9v6n
FeITQG+LaFgHEG1M3w8QexZPu76BaE3IZqNG52Bkf4LQftM6296szWSDSSC2uBSd
f5xHiYFctUhYaS/d6ZLsWYxQjZaxXwRSbAq3dTRk3j0qDyZz21xrlSs7P9YWuDxN
fVw6t8bOBK2zwKlJpfgNKMG0snlKlKw0hkxzUDZhZFoEjojHHyRsEKtg9x6pD49u
YEgj5x3EBR7cP1U8HMuFi20kvF/ttyHYahG1GkhkC017c4m0DfHlMJxEEQAohYmB
vzHGkNvDQUIdNo/CQgVNJSyPvVUpM7Vapcaxp9DXuIckDB+jhrB9TnTc0d71u+gz
IxNowkTHsRwTqIVRssrRSv2SWjquZSowN6St8Wa40ij7iURxDsH8DQ6FJ88eXnLb
aIl6MDCw5PHbLjUQYs7639wqnvPj/zJD8FogkjvbTn5ofd3XhBKhJbIIvR6UkUgm
Eg/AuiUXgq8SLD6D047cLm3DdERagumgdojMv4JNZSLQAA33HQuer+wGg8INqXud
KEl5mK3j5CDnM0gC+8S5M19LMutIFOrIDVP0PA+E+HdDh/LTCo2GKqptkKFZvuCu
SCxygX7u1KpTMLqKTf/JVkEhFU3qkS/8RNEMTpJru8mxMCKEIDvHsURs2BSgGdP0
3K/OGGImq0imAQvzKlTQ14u3LQQOScPbMZ3IKFQSF6P9XcdnlsIu8PNNBQ49w0di
YTsOsiaF8mwSc5/5+E5AuUOepmMsAqiG37wwikhbL1nB/ZYYhb5m9HXuGVfbWF6v
46eKwUMWI+7HxQC8ZhQXqo15WHZDiYXcwik6JtxQxiTY8vx2G+lKIBOhpnFY60P4
RV/xSG2Fwhdd7eBClmh2GAUB4qH9uN7CvPzl8UgChM/ySV3mjV+if1tnsvapF7mt
WEjorjl1thhxbGWWsSKZIu212zna+rOSFHWIIh4q+h5d/jwmMwY9JMgFt8niIdbR
2GAs3ba7IBYtkVAbgm0mxy6MnfByjmMMKZVs3GdQGJjw+Fos9flXlaMzDKyZHZuo
mI+eRYRhJGfM14dH57kCH0NiTp80S0Rl7yH6nFccbWCXYhi29LHfgExIE7CkD4EX
rN2d40IdOfPmyXd/7chGjc6CpCjRCjDYtGO3XXvS91Fr/4z5gnPa8f+XNeYVBP9y
EfwyTH92PXlMlsNPkzGe511jcW7NBkNpdRLrFDqYU33ckKb+M8C9fnV6qEBv+Oic
RZ5mg/h3G7D2FAQXqSaapbaPjD4QwLXfj6wTk2l/zTD51MWRh+cZo+b0pr2xDtIT
5Gd3kgyD5DWtlhMFn82ElCTKWsFNcZ4jQ4z5L6VngSusEPz8n9g0ysCc/25Jtjz0
rBa1jy8z4DtCvzFxBr6qjvM+ZeVSM1p3BEJGbz7p25QvmdgdFtw4fJcnWpB8UQEE
tAuzkiZd5NK+BRCiY9958tYMZ2VOBCN/2ravdqa72Xae1BdqKVIGhheoRUD5yNwW
er1xt4q1CyfKe09UAy2dVfJYguy0jc2zcbAo5vEAV3XrDqTqAkwyTWEt4nNpmBI8
RlsAfofVI+pa2iP6zH7beynyoxOAZH1ZSKC/BB3xngGrHy3Bfi0lT9uAtZ388yuK
qR0hpR0JGZ097YeCMAiA+2vLLEijnn2L6ahY0baTUjh8CjFe36VaohuTpqWZ0JiX
FHd9gIwBpjignBzyLMq8cNtf5QY5Cw52knT4N6geYeEdxfIkhCJiNt4vAjSnQSaL
Cvpl1UvIz9FN5awavFk1ov2IiCeq0gWxmLzLPttr0knCLrsIIBgrmmJRQU/fbNDF
red+A6v79ndpVO1GmRixfccRtz+W3B8D6/DxOppzI8OiUItryRuv6oWKAMwdkNuJ
X2wAljiyss3mD8XczGZmPrExu1yyC0GAp3gklk7m3KXePYeJKrKJzlSpijeD3fdo
n2V1dq+X/9PbPN/VuSkCReL0vXZnKWS0s8+QzPSZAvSfmuwmc4GjoQGGpT92p5xW
uCBR/4gplRSJ3CaXg/BxYeMGjIa8geEy5IjmHUe5A3dwz+keYxQDshr54U0E1Trj
xx5NUq8SaSI26lxOj2XQvsaoL9uJw23EvLR7eO8HJUuwq4HQZu4IisqqEYNm5/tM
GnuzudZHic+r+8d+H0t4AaOhsI/pKeIz846MdMuxzp65v2lrsyhBFivHcqOIJkTs
L3iPY5XWKzApp2y1qYfilwP4ygA+/yCi8QDdtNzbBQiG6NLbsN2SgwWv7eu6bfa3
ETYpkp+xOMLKGOnoNk/kv7/qwoEVzj9gxZ9DrstPOTjshuHQRMYd/5dIIJeZOrj7
TnLB3bUIhme4sf3/eBIlbIXOL5ZtfmleWWerahqYab9YvVy2ZvLqi4uDjG1ljREu
4KT433uHF3D1WOWeI7NI8QGMiHjUBLo4KUHhr1HqWme2PWiuOiPVkfoH/EbMq9C7
l1VGg7KjBBErUBHk3hraAHJTv2nD82etCnNtRjN3HS09t6lQgKETZ42RitzzIdNp
v/2Mutd6Ut9PmNOS8QzSqsDLRpVa3HT7aEJAl1goWOT24M1FruV7vi3a/xPIh6Qm
ZRbULf903l4IQWKDgyCUE/3wzh6dyjuzck5rjB6CIsZ+yrtYNCgkynTsh+SV85Cd
kzWmb1JtmmNwyiW44Gsv3uRSNz7u+44yh8jhlBita17HTvSoPctuUYXc9t1GtU29
vOEs3lLwBOa/O3Tysqfm0eLT23n+tKVJP1VaG2j9yWaFQ9rDiG7wVnCjbRE5icOR
t1GqXTkc0HH2VF3uLSggHqKnx40GuXcmXQYyGHfLIjhUw8YrPOq6Y85i2FgW+B8e
kneMG6r3FeidLaTzWtNORKtw2JCGszmyhSdCWhr6LUp1YSFAy5N0VHX7WgH4Ueys
Sz4Ff70N48jHSEiGoQp2ReMzYJPwZRKgQVSAPKRKzG20v2+zg+ANYwVPwaTofBjl
AesGdAsDbk9G2mUNQ7qfwesPZ3HUC/GNilyKJVFbkIEoF/OcaSwcWGRp+694Igzx
QdbeYHndHLYnI14ExHoQd9Okptwv252B2phNSc6+f6iQTK2ecBeybi1WYLUERm01
1oln3rs1xvDkyxqATzx7B+3T1GYKgTf59nfIkqUl5nimz7pFF3Iz+Neg48e2BGb8
2qsGQ0Z2Mrc6uqxu1Cg0HKHKHtGk1MesUgtlBNuRoutxQIOIjSiMyhiDJDPvFFi4
ZjK3dmQB4YZVfDVf5891V0c5VPbH/EPl/chLTUxXCkndMJPe9whRhREvh389yYpn
AW7c6aIYoBM3gN5vAOPGQ87f7Bu900n7wzQrS968Fq0oqLnmezFENNllxVJzhXzy
cIbFDdWTg6xU6jD4aXSqKyje2QSjFJcNXhhDy7hp6pmSwCieLx8Y418FriC3QyGD
93VY0ItCyk6SX8+Fbt4HQKH64UVnZctIzze65jGrtqMRy0rUf8xrbeyjTY99RuYW
GNP0bLf8wd2U1/+GQKcF97zbTXaJVtVvctCvH3tQhA4cKdUEl70oEweQpyeJ4qAq
MSCHtJmF34jdcFTUxJ29iiBA6+qrn5xR3rOLxHhYKYhyHVxtI2WGc432uC3TpTvC
y0IDAC4OkdAhuEOH90Yvf6wWgDRYlczxFhhJzdq2tNyG4eNIGYL6MN349H0T2Q5g
KC3ZVYn54HFIBHH32vBONtnbZf5H1si+Q5hjkeoUf8YgAZSyGYOlpqe9WhTrWD0r
IZcKVakCHHwsckMF7IixM35j9H4SflCEdP00uAGUrdnYTxbTSEiVJ+kDlb8es+EC
skyReEPC1fWpy7ZJ7A/drCPUZnn2bQK1YOmqt5UoQbx09bls+9tajYnSsg90UVgu
pZMrGUqppJKupgoRsij+DZn7qD5cDSNTkRas6p/uH7+PUyyNqjsDfZlE24SRVNkE
H3yQXcrhnAJu1cnrcwNo+3ICzp46/0bKgrwmsabBdikR3JSb80kkXETd5/eAJdHV
FlNAKD8zYkig7P39rrEt2AgnxOLKlSaqZebQIUZ76oVTfeHdf0mkUhRUJu49a3S7
8a9IxKe4HWqA8UsRohBLYSDzl+EJO+3my0WZqnocB+0qTBcb+44qWkaDQmWhMtPl
lpGW4+taipHb25raQDa2DYcK/Fo7Y4Sk0UiCsrHdD4tWmXnmFD4FTcN6JMcecrdQ
84FJiFDgJnPVrCgfaRzTnz9GwLgXjz8bjdRGBvm0Hc40AbaLIb0XGR1n+bbAPqr5
hduCLVne2g4us2zJOf19mpN2qY3Xwl2Gnl1+8luTtDbfkuMpyaWRoLREeAL5MQvd
RnAwnx52QMpbcBzucf+tUXNT5D2HJDcmlywOqmgZbORZInLuMZ5WrP+x6qeOD+Q+
Sx73SKAqRDXvJK5LT5vMf2M69A4SwtRsWool5el1/VwcMD8HCbwQKAslRutjb8e2
Ljsz4NkiwUn5XvZYMqQVqmZUMk4l1bJcW9atibY3sOVTrdunA8g9/jL5MIdaXmb5
dAqe1qQC4PBzypX7i+Ki3XFYY/Bmk+MTuBGZDTsLuLmfVwXWRBvTvTUErwpzjeY3
vKx/NqpGADfxYGTLANP5b4qvMadAIYGTbU2t7kvhoGx6WSfG+UYraGX/+CdRT9dY
aYeTlGj8PQHDq3NeB8klUHbs0yOfpZygo6gTYTaHwENDnZTrbZO6AwZXx9P5UhuX
SMUp8g7+vFGuI57RILSc91w60/T7G+kGdX3cYN5ekbZLTR6l3/4J8pYWNzQFaxMo
ISKpcTPoIWUe+qKUTAPQZ/nPGZ5+2zh2SBqljOybkp0+BYRfYDBuK8HJc9Lt7Y57
+uGPaBvEFxQ9jibgXZkYiQxfVxAnqm9xMjpzvErrOFdV/gculob/DMdbmpNq3mCL
LRFB5iYP0BGsUmPMygogz6ZW5UX7GtQvs2tLA0+QaLQmckE6UK44qzdY8cP4jPaN
3zgqpngkrK7qOKkSGvMag6qIjT3WNl7L4QOgZgPZqdBIiKnhG0C71Wpumdwu5BNI
x8Jkc6e6YPnv4hsVrQzgiteNGVi7qjX0jFgRPDJYk4+ehya4s2AnBYliTTGoKp+S
HknhSX8fP4Nda7OIYRljutlC7T011MJ9y1qGr4OLm6vfZJBwULZ+M17qE9MBZviR
Sc4cxpuvxH7Qt23jnE6ugwiqIGCng0DkWfCyfJBPOdc1mg3QbPZ58KOljPBizzQ/
dnlGfIjMNpSjFy7SJIsM7ZXSXaYzDK4ZlJBlX/16t5s0bT4DJtAJtqrDb9MBHSXC
5JEgYfbmfA0zLbymmI05xD3jSWDFZ+Sb/RL9rF3LnzgTdfCGWhD9PkhF8f0MV+Ci
Ae+8YKboXcS9yC6UM2EY0hMT09c2sqY7k3UrdZfeE+hDMOx91AE+58WO2fgbofjS
owM5TJRWLcgK+7jrrqx9FUQXystUloUrfdEG5mx6+GRO4ThAP0rfYPnlEd7FwRsQ
F4wBXMMdpdfMw7ii5s21z9CwyNWfhCn1EeQR57RuT7q5Wrc4F+b74kEG/ArDIMPk
AHJ7LVrmyjTR+rpmJtY5WvEzga1O9VQHv6g1H10tcY+c2YM36oIE/mVHE3HxPoqw
0WvCZntIRCS78JXbx3poRAuJncw1RM/utW0kzzAQwW6e+S08ZrFDpzPhwrItyK78
ca4t0REm6q535qdh/zeVMYfSQDADXnfDdSI/QZBhArtCFbdAJSgyqWBtXT0031v4
XEwNNUpFJCujq51lB4MYPYC8THMx4s/Jyd2uN8rsPbRtVuTwwavIUpw3nT3lUr3Y
vRiPDSmCa6Cv+uEs4VQc7ZzUuDQTWuoM6cTMp7ferEHq72mWOt7ymkyrf89AlXvk
Edyed01HfP1P+EPiYy8Gir5nO/aXuCfBaM0Gy8FhZxz3sQfOOmv1T264uQh/X4qL
Vb5p3wCaJkc5ke1wknyAlF4EvxcMygUu1/D/NUv71bU0tqFJCxKjd1A36wjTQM8k
mH4bT0p37K/2ce2e6LzBSFvkM0Kgw7bK4avzBLtET9rzN+K57J6DodB/pcWg9v7M
zk3G/LwA/0nMwEKLw6C7NnYNUcJKq8z1CjBi4Sb0/Yiaf6nijVe69d+R/t8BwU1A
tzNDGT9QNOY6AdgFAnFUbVE2RvFWwFah6yVzr9M73e+TCBa9iVVbqcrrD7rVVl+Z
mEB8G6g9zK/C5JVXCz70edMHQ5cXKBzhi2XmfzyuqIR3ZOQW0s0Ps86TDwmT+q9+
OaeXiuHaCgnEU8tKAsAl1EhjSyzmHNNw2K3AGRNLV8+SZiPfnYasWyu4NImasnlV
8V9vdZ7muhZq28VCV6PFOr1++FQRhuQwlCN0EVxmgq53OCfmaWkbdfHqgTAr2ogT
iVffAmKATNgo8XdhqrqBuvP165X53TtBCtJ3OtU41rQwstk5m1CwX8HdzfziUDj5
1hVLV53hn0fyd98j3mbehXPcewrtL35dKS6RjIsLg/KU6Omqkkgp9fI2XeKH6/bW
pn8dQ+RC4ZsoF1qoou9m9TctSuewawzLGaecg9eWvXV23Q08FWaGL0kvJMU+WO5F
rDGgBmO9sd1xRz6EHoSgaNnV27d/V7uH1nTZkP9jmfw4mSv4SRLd/YP647OrHXmy
6LL3OSki1mLqm3/0HjdBg6IrOJytrPpVzOdeSqQV2DC/vgjqeQLbllD7PwDgl20N
2SrfjeyY0ik/oR3IvvoRm/eyaXZev21y16/Z8alKIlwjRqWSfBaYCnhgJLtvn1UJ
BlJL6q2hFfBIokkERNZo6WdSRSJzN0Sy+a+EzC4KfpxaJ7P7vnEKHceWp/Qp6+Rf
loLMvPYn7bgCZDQOGT2kx7nafpz3ibwLBzopO5FcYTS83yZNMCIYU2kxhGXSvSbU
ziizkAV3ZnniQ01NWY+oiKCII4J8Ba+NZ0lWhC4wgglMn9GeZM2Uyc2JJySm4h8z
uIHpOPhPHnLUzIkvE0+e9X1o5tcAZHprgTUbyL279Cmo8X0jM0rR4UL6dU+ehFSW
WRlSfawWjwH0gWNNtECjfXai1kzQygNpfpI+Q9m1ORYHdpdHoG/DgcOE2U43y+aQ
ngYgbk137ypiR8lUdbZtoqy3+yhdbGP4wX14pXhXwg5WCTR8VpTpKiwuhG5hR92x
GqvP+djXCP2ckj0tbB/vYRhxPHAxBF9TyC3g0eEirt8yNPrkm3CeoRFO1NqOyBFg
aZWud7IPKfvm4HWqECIHKoiAoSzCuZ7XRpBBoBMNPQP/WAWGAOHc3t22hcr3k3+S
JWBD3cVul7Maw3061itd2I9hc1dFs+a6mO/6kWhKKzqtuJky+C3T2rEQSjws/z+s
ZuUps9VXs+lHof8u26TYrfpx98Oj6qMFhmXpd3aqITi51PZgjuNSDnnfVNW9goBY
JJQ6NqS1X127xqq1t8WTdsX3vimIxnKnaTsF3j0222+RzYB8l3K0ecujAnd51yo/
Wpki8lO1RRuF6HlAIccRF8O2l3Jo1EjYK38fUu+qCAw63j3agmVoyArBVmc3us0o
ZH4QdyC1lrYtLNFPDxfMFIi5iLinwYtQGrcDSeGXPC+3BUCVtLrF6X9hI4EHa6gH
ld/dRdIwScbmzstcerztyD9i6bbnU5YNaegXWZhKQfdgjM9G9LHxfDvKvDa1cLZN
qkF0uNq1HyfaJG+YawZKwzQImqX1ob6QCdvD+Y8u33RVWXqnzYKiDORsVOCoy1y6
TvAjyYJHR132Nym/1p+RZuEhxvfjiazs8QFpu5fk//CGU27q0sH7awdpQiawJYYJ
XWKex69mtvkxxp4p1hwMG33Jl3O1AKfYYlNiFqksWTIbeDoMBsIIAdl1rkGbR5tz
ZTag4pG8GsR3raojVLkKiD12cC+BD7aEdngpCTbJzVWhXHGx43fiXOg/NRmJUIYk
B3fXUyu1vXLlSNyCRIQiF6J4KJI+WiKOmLn5Yf61jrEvFRt3uo+mpauUq6y3xaRW
I+K0r02xS6T9XhshXZm19xM1YLv8zQPVTKm12yOG+4+VKyXezGzz3ClKPnnUFv4v
1blaF49KiWufnHBXJuVXZfO92HDk1xzO1f+Gkytsks05QlqG95yXG8vtr7l3uODy
36mDTfsNvcqeRetDO7sv8bXV5KhJPtYZ+seHd09uIxs1GLhuJsZvnNmY+GDgYQ4i
Lx5BOBgJg39Atf3HoQNkcpjodaG+Ouqqf3KDKvwlPNk1WLiXVMICnhfZRcuKr5U0
xzrMAUXPZ9SgjUwWI5G1VoxVkDqh9vH4B9EG6OrbO9eCAKMHZfwJ9Drh1CjeyC84
wV8oC5QwwTG9VS1wfY9EYSmLt1eM5WiqY77NwlEuctQcr4bbIT06/eURRwCIuTvD
eEeFno+SgBMvHOaFfbbGYaGqBFY4HA8i5zkT5pn5jQVrKd1kI1lkTAWNmi9KyOlS
M6nz8kBvPT43XUpi0jR3GZTlYE1/GTFQnw5x3LLkSfSs1NJTQfsbzcjaj/OjhOfR
K/uGo/GbrZyLPupofSDUjZFuqBrsiZ1W6AS6SNJ+og/pwwySP1TIJ+5mnL54w9ie
62Xs7kpV1R4TJVEEoa4YG/BFP374csEMPUnnVpOPHMk63NxHRHFS5sd5mC/U0QIm
BYmwtQfTDwST9TS+S3SebQWdYQRtDN53lRiSaE5Qmm876JlNRxReZi0u7wk0may+
9ndclT/TOiEzeG+Ryrq0AbrxBx4EUX3WywTURQyzrfFVu5P/4UE1KpWmre3YoUtc
bglrNGekPfGCV01385OUIjrhmpgT7DnRFfhLR0WehU0/f6nq+jnJTA9lxblgb+Js
GlNsIjJtyR2eWn6AFzRXy1IkZuJ0DlppHEzBq8bHETazmhsnz7J5i19DRiVmNAb2
Ak8jYOJVKbImGkDOTCpKdR6sr7eYC8tGw/mEPX/PstdE7ZSKY6DTt8fqMfqOpL6x
YWecV8XKCJ62wtE+3mfGBpq9um43jUPtPkKWFpnr1JAM0V1crnqCcq8swn/asq+A
NZpD5ldiExaHMAri5cKGMo/xifQ/3ucF369FCCiAjIjdi46ZdZ5PAX05ahGLmK1T
jjlPOzSxfk9WJWHPlEavDCqq74ZUheQDh35mONtLHDPJLcGTnJqXw1Ojhv83VSnI
VxdR8NnWrB7xdfYlhcybWEGsr0DFvRN4dSVGTfP5LupWW17TSAwW1pZoQmY+M5O5
WKGeG3LykVDmD1mVKrCjeuS5yU4KHjqm0ckjYZltJb6ty1sBFJIpk+16W9OgJhH3
YBk7dnQ2igpCX7r4a5aw6gFoDdr/q0kk/EXcAth6cpZujgBphheAURTx3dd1wLyb
JSEpaaUrRf4LmsBY5sQFeizvse2blV+1kLF3Zo4n+2K9i/n4j84Ixn+h5JrMZHIy
NLiFSz9cR3OlWRcmB4gubZHHpDIJIdHfTqJYpdVSKr8TDSnGAVvvRxsPlfJ10qjg
Gx/3IcIcvrttFLZE2+fVQs+yv+KWUIXvo8wItrNWIDh9YkmU6rcdbwzYOxq6nNOT
+cIk3sxWWQyhJAG8w39L9kzGu8UUApawMt4wRGRfrxypyWYSxCnFG/Q80txe45ZK
Jk6/TdHir/vBEuihfAHiXasggbBqU5RvaC1FnAAwQrgEmkhsJRqDtin2OY+IIcu6
Jr/uIYi29YBL6KTcPmiKJgBr3UnpSyZHp7G5gyYzt9UcQ6m5BJFSS4jwRhqcjrEQ
/9uKTRdRFKYrXELN+jGFJmtXfR9K6inwk/c9v/4qgUJVx9FtGDcjFb5tcG7ofxei
sm71Y+4LBrEEFtYKbdmOuirD3KwlmUC/mRYdhk1aelrLOoq1bgBt2E6t7lIOUhoB
E2rtrF3wNT+u8iZK4my+s2wTCPpnYVwSsqvQrCUWpLBZSfwfeKogSEsYTQZwHh1T
tFOW2os+e8LDrrrYI0aC4/YOGh1gXUO60G+Td0XdQPK0D3G3sk8LHcX/iQ5bO1SX
klDByzu7CeFq+E05T7RRA1Qr/9wAivT5hqrh/aNTRV43D5AWpDsEY5sehy4h7caz
umJLJWeTNd69GQPjLvwKLLf/amBzL4HQuIZBCr4FdJJDgjU2dvcxcqxpe6acH8zc
8b1x3sXhKmsnG9ZIjDSq0ElBhlUfoSwAwkrMoxpSCDmKYgNGcwHMQ6JmDGGZsjoe
usxIF9CXCA5hsano+8pIgbjkxF91mTQhEZrVQ6qKBnNtMFK0X2NhKwFhmy8jFhE8
qowdXSnvvt0sLTTyZMBXiRC6a4jlL5wZ+nD7doAkyJxcKUUuq+hv6nYkmVJ+dmjZ
TLt9Mz9oud/eMCEUAIhWbACRfisCAtZmmu5m1O5qIFIjOc3x6X7MIyfnJ1Rcx3FX
gw2lrXC094UrUTDi8Xam5vJPcrgxWs8NRqi644wyWScwolGfDSLmfH46o/CkxC/C
N4J7kz0f41vgseEQ9t54UllLwsJ69RyM/QeAW+PIDmEGIGtk6fT4/3sYfCO4mLs0
c9jyssbuEmoQ2HDD4wR2HelV3kmahcuKaUI5EwDJIbfkx66FUxleCVCEm6eX40j0
/i5ufZYRZESefMjwNkwpT69NHL1Iwhn2PttVbUWS0PMt6EoLSkDyr6lBKALTlnjr
su4lGyRpApvB4ABnw+IIzAI4qbtBGUFveL1vLj+rc+vGk8lIKXrw9D54/5wIO9uP
eyzeFJDw//0UwlVOB5iKjqhgcwUl3i+3gggNZ5fL+Rx7duIDm7+RYUmA/yMV7xvD
jIsKl6jh5cChmwOZ/v+I/wf1idSzPX4Gli/QXzGxBbxv113484iFYN+5fUMJ/Zud
MMpIboFMyOoih3AZEEFG+7KA/CPWejX7GlQu03bJNCHtGK4wKvqSiXvrf1U4coxf
j95LG7fYCXSl8KVTvipMfoqmOBCVE7xEvP1HWmVZ9awG8OPixa41CnnRoCnVFmeo
5KsTClTb+Y71f4dIXzFz5GpXNqH/HjrGhMaDLHLg9xZ1Z4LH9iaNH6Zxc/BKoNBM
2C8VqB+R+U0Ys6qU9m9AVGz2AVLPaZoRNkYl7yujszzxNrgXdeuDWOcXtwUF1BXB
qzAOCBWH09R2SumtDqOg/OE0a8cYsZzVvSejsmE/RArn59ZD/b85Msoqv8TeoAHc
vlFfPuYMkawAY3X5TTLjmLvqryXlqqO3t+DOUqbi6/U1QtG/aT0Vyv2eXw9mZoxF
cV1cEPSqdwJnIYGMlvR23tnJk9Ia3pibzK1WaZHrKfrisZO5KoPeKT6CtXHjBIE8
5CoUVkGhgd3sg4KVkSETbfrs09qXCRD1r9HazwNdgGevlkLLhYoGkYdyZL9ivwFx
YlUQ/Z6AZKchxY0vK3HUlTpFfgnwQkMGUBPpB6EYO6kHIegFGSkDmE1NBT0Hfbou
isowlBvUYQhfb5wbYc8C0V/+n73a2tFm1Z2MjXRUqwqTmnw/ugZRP067ThCd/acz
224KUGmqTUvCys6RHFvYWEZlluz9xOuag3dUjWjoGTXl2DPsGuiH2AhjOmDa8WQ/
42DRaiedX5+IBOy+Z9xTm3TxymZhNFXxrPRnvsr5qOJtUkTPG+nSdpbkkS8adjT1
27HNEwhzBZDHcW194bwKqvpR4xMVeXb0YQAnavhkwDPNgQl/AqHExpFQccscTfYy
BVqV0Yxzrd3eAmNWxu9PUw1iR7ykvWkqO6A6PrVvryuFd01mbabZ8JHAbOSzc1Vi
Wqhg0ua9af6FhT+YJiIB8MegC83Jj8fEBSlymk4pdgIg1Fr+vv5dVWjmObi/zk8/
gQ+lmee1YFBIwkl/4202k/BR/tWvF0SMpMmDbTFwQj7mq7id6NUKzEONJilJUQMH
0HjlzjoMIxoS7pKWJtdQBQLnZak7tUUGwSm6GdrcIZXTlz+bVQeXo9FkQ2qCrRUI
84lq4SIZq+2Oh6QJ+Kpo6jTHNFovBCv4lGIWEgBCD6r5l1E/zAyXCNfIwt/qfTRt
JNeNVmmGZpPfV2ld8hL1HOdlyd0TvDOhPXiByE51sfiYufptUpeSJkfT/4l44oFO
NF+uCr9SZNwiAFDKRhXdeuTkcOIKBg1AsVH+//1sL35oChW9gWHA9MRrOO38agnU
K3dV0Kc2tEN5EYdZRuz8kBNRhitjQZyV3t1qd5HjPaowlSzH2V3Rgjd3GC6yUcKc
Bahy5CTfSLrdnI0cxEhiTpiIQ9fwtK5LrroSlywxJdDE79KsHVPyQ/DlkjsyR3Xf
dZ5O0x21yk9MtGO/ZQjP7C794a1FDen+THsM0rphJ1CBTbXfJWnk8PkA/Pcunap2
UZnJ73Va+323Y1RwKosoiKOG+7BjHsamAw04RxjwQ5BTVmBrSy3qLbJ8OVS7XzVT
FCSH8BQjhYlrU0f2xvMBGTlIaUpDYWkZwlYpu5kROdcNOrJVcIAckettM2B8aGhd
7b1D6tjRXL9qTMvUJ7vpaTCOn6qGckB+R5AGhBiysxxx0UPp2LzxrbiFeNHPEXuw
KrMunxWCIvPuZOzADnxj/IP9kjVT2K2JUqUtJ3DCmRonOYwdLg5cmnM4gNHO+wjj
mEc2Qo9fualKC2MhWwVWYHX35SCTVuhM5IyauJvCIlOK/OpF4k50cDXjH8COZYRh
1c4Lhyf52RWBgrHeDKJh/TGJQjIEE7THe5Hu6HYNNvDlU8wAEq056ba7XmbIo2Sy
UCrLcA6ApOYTAJ69ZHcVUSJ1vWD4C3apew5xHMh8jUt5+6jDo3mwm7YPW0n4Cmt3
ukgzD9zoorZVrUs26TzCUIGknejB4LkFb/OqL+pJxOglra4LXDf4NxnlEytb/67t
2eEP6Fg2It3XYPme+1tjUFi0ylnFWsHCidTeuKk7+Gu4RN6YUf2801Sb6xK812cA
hcCoIx6SnXaUVbDItu9P/2bUjw3sf/CYVCeu6arOz7Z+2TkpROpzhfcsWuH8v7Vz
sNmA2Yp5n5np1lW5ouSjtHI3TiaGL+P0mVxsCv9O1SUSR3Jw2ddqXHJ3kqZiOo7t
z3Rq7TLTY228Xmc5HGRF59T5dTgVZktfcTXASkkl2b9Y1tZl581RcG54AdwOnwyA
6MM/d5DDmx7aEJSD9NvjjVOL7Zg+2NpSgtuCztPvoT5filG79913eiQ3gCQCQNdq
8CD2gMbSB6DZHLGr6BNoFZ1Ekl0+biCnUyFtBaVz14O+u9sj4NpCSOwO/RB6DJ3z
xs1DzZU368iGYGvJySSUjBhbbA868CtSEFQSpJLO/N93PeVXkS152D9WUX5wCJlc
G1CeFRAfHyYyyn5w2IIQC9riWEx//aUoNsnIoJnJIZ2NRAnIaVBBzehJ+SXkdJ7U
2APQ0m/GITMdAKNSvjt5KBXujcaBEa+n+8zph+MU8GU0xyVqOetLfALYBzTc7+IO
JjTTPIxvZ/sJAIy1/hL3T5bFDGMimXjL5nknYBWQ9C4Gzs0XtbXcD4IVY+TuQFeC
rNGI4PEcJqUaViP+XyqNxPksDrIihdsOvzpeWYOWe8tZc0swNvH3ji7Hf+U0rw1Z
dAJpgjckd5iW688qlLGKpmsvNVVsGeMGQ9AdJWLmEzqHg6UttVMe8wqLHF2ktRp6
7uL3NofCNF7mrK1GGULPhoc5DTWl4OuHawsKNDt08smsD71piGbnZxYc3gEPeMJu
kSxX6mdp3mB08qaY6FCGf0glO76/XNdh7SJCOg6YfW0EJu3i4gbeQovJhWOwoYhC
97cs/2+61/EmQiIIqCleglAV7u6SECAJFpmhMfQ/6axhQJhVeLOrR5XP32ziW7Oi
PCwxetbFVz0RtFGa0yIdr9uZHxV+gFMz9VvLHnmizkWGu/A7YeAKgwIaQspv0+Vw
gPAmQSHqKdzdoJZhqY2AvCHfBBIxdr4RZfTo/AlQ5L5alWmyYBMi8px+fsSj4SAl
lEuB3REjNMj/VfCMBy0XKwQgsb2ZNC16cNi9QD7XPVBTiRmLexvEs8FTZHRCC1He
kaew3WCjvhHgkwZxEOETuLxgXYmsqPIvbvcSdkCZWBJpirzxf5EwMzwhMfwfCP1N
JHuhDmPWiHpMWbeHRegPAowIjlVjFcOOVzN2wpXAPkZUEGUa52PlELKaGZlztYDf
iN4h24wSsHVWaxpzonGEH9AN5rgrGjEXgBGYOcGF9rvzTCv4Z1fZP8pGRNhrsugZ
89n+S4ECvYFz2EGk1ge5iPsNGVHuM6yL0ivu4AARlFqLx7dGKNK0Q9cx4i/kTqaU
a5irN+qH9IO9ubNpUU5OFXW3jFH+VHHBV5odtx48vwZWAJaFe1qMSeCulpuO7h6p
ZXBlJMINT+mu2UOXGyQ+gIrKhdMUYnzzF9Lcfse7hUDlyhM1mmJavj/86dn7ubUW
6vCx0j8TsnKYBYyKtZWenv4zIEyKW0v2ls87c/nV9+eRNBNe4XPZ0SXzeo9Vs7lv
tHZczd8wkMTpWwpyLV+hguG/N/vnctvxY8LhNo8iMv4Hnmjps1oV0C3Nbrm82lfH
zMJhM9m6M6WgV3dJITG6r6s2Y25qnmfzDSSIn3iGn3/UO1wG5Tfn9IX/bdMuwDyd
MFzz80w8JQdPrd8Z/DduZc2znvNyvmiJs74ZOLBQMqvpO5chu42BbSynUsEmAOFt
16bMVIgAitgzzamPMlZFGIpEfVxDop3AaotkOx3H/4rxhBD4nRSYAuKXxoJMJ05F
jY3JnrHhcKK2vCCTiXBIX/8El5OvFfRHm33z7LBcJLXdNSfGcHNJ4XewzmKif1Ir
AraWFYvqTc5AqQm4Vw9JHRiw3kimWKc8ueJS/oHa/tXpOCJqDPHolFkO+ivb6Db6
l4XZiXQVwz6kEoT2DE7uDIncT8snTCebdQG+sJC2mLog037yzgZWXWNmzKHz/ymx
wR3Rm+GDKoQmvPnQeilaBbWnZFD+CKdZu+uopVEttdUahYizarG9JoGnWZxU7pfa
jzUueZMxObJ1dFq8EPuNes88VxsOuZeL8A9g7W9MuFqMe96pQPFwaeLtK8UZM90q
467Hk/VeIKFwP71945Ed1drrINpWXUVWx7NZrtVS/oQq00+4rdifozvjudrByqpa
/4u1fcWTXISg6fC9KlcGjHe4e4hEjMzww4qsNEwDXaHIwltN21hsQckeZuhOA9as
9bqUkdfjd3SkhDVc8QpDNDluN4a2NwcLw7Nhp7kVG+7K9W7f+8kRz4Lyrojax+e2
5L7LMkHE4jAfdKEDez1w63hta7Fsrjz6JytP0/bJ5DQP9UurqaM/Sv0yHJP+QdIS
54Q1rbwEMLRattagDfmiv06xvaZGRREDtHNrfrXrTMkf6j5xAVVRAWG8dWW4yURh
+pHW6ezh1MV8WweEj8/0WE914ENde4Gs3VyK2/HkbilIsVGl3AQ1QH5q/g1nIi0k
Jb0B6Lh7EN7lrg/e+g05NE+KQMDI/tVFoX4D8c37blfhu4uQi/UcTJbwr4x288HV
PqZ2cROD0/rqC26N+zAsNISfbSkyMzt7V8Q7E1u+GSrqG6kpL7QjhurzyKa2eLpb
ajC0s7X/IrSPANVNCqNN+wLazwuWZhRwU5DWx8Y70U+rwnFGyZxWgBvdGk9ZD+Nv
z0fsDVTpSpyJn5ApaqUqDCSH2oR92Yc036u8uzK56NWa1cDzhS5X9McqHtXvTWEZ
whVrVKGie2zB0mjo1pvYhIVWo8wHYy+Zgv12tsbMz3iIxW47wnjWhAPh2abmGl8u
2SchvUBCMXY5OlzdrrjlMubTrFhoY30n2AK/UQ9H8ryCGktEow1ae74PQBDlsby6
JK188z+Qxjzk9mrJhUDDlAn+Z3lwe00U7JVQGDEY3rf3T3BVcnixF752aAOc6wSj
CMSss+7ujzZJfP0IhAi+tIPk9jJC22/npJb+Tf0EgJBcSdmjlfa1tSod6LiYr7Gb
mrAb6tl6KaT/T1pXTfS+MvOCdBIfu2wLb+Bf+wTG3UAOHvP7QY7UfZZlibcoUtQ7
ZB4CcoHveAXWtJ+oNhCaqWOKyswpujwQs9Rts4Pr94iJvihsoZMa7TZHxnlJ2EjM
ysauFEWx5TCEQ1928nmLD7tT9omV8g+og9bOYtWpE+Ng/36atxfkTIFq1JBDISi0
oz0Tbfu7js6UrLTlYbE/mtJCxjN+Emo7M0jUzFxnqy2eggor5XGPltIf0kPcny7P
AoR7pL0KRWeUi0UTgS48+eibRfJgfK3GiL33kM/BAK3R8Z+kbqc2nmLa8RcnYXFc
VWjrMXQAOVsWN/zqpS/D4zQhUCEsrcyhd9Hgjl7syJweONjGmlkHx3bwsYGabjXw
pQjDXERgirfqB2lU5xhmbFfitEF/+vwOROx+sVdQMQ1NG7ttaFpndpoul7uLq3vO
vMiI+3ZcSxgMA2BkCkLZQ3elFrVRdY9+23WN5MKarcxFks8qqIAC8DIARXl3S5HN
az6OU5Ngf3YnDo5qyRq2dUk3hVR+2M9QZCuC1fmadzbu6gtk2PZrIZBVAp/B+3jL
3fKPECT8VpQx03q5LDbzyDRurETOo5PTjXZYZ/bLJXv5o+opfutpMPwV1sljWvN6
LRlC8Rd48nWbQdTUit3c4iiuGhJ3Gf22RFSN5TwtQR6Jpa7Bvg1wtckw7QwWWR4y
NZqScSQckyv62jTV+GdnvSTcaUiitaxLlBzaccFkjzRRsaL/eE1YoNDwsQKfM9rV
Yv+jjAkzS6IVuYJowtbAgo8qZKnz+t8/P4esAkKRTDK5rZxLkLYfGZbsob6ytHWq
UfA+kozq1WiutxudtWVNBJP0iTMRmAlJm4Y/JALqD0Tw2jx71xTApmYJfePaDfwT
W/j6HyadFvm3I3P2+D/PUqoSuLIgQyHB+G35kGpM40zseZ8wLtCISEdIkfH1t/yu
q3gNDF0uWXOmQBWNSlDgsz0Q2kyLKXSOIdvInu4n3A5dsDw6CWI8LzYG52zVIK6o
fYXh4iVc8jAq6igZOWx/9fu+GFsKQ9k32nvTJQXys7AfToy+KkmluwZEKVSvKql+
D6F6Tyh6qx9N2Gu1PtvWwMZ0y2519VaauOJ/hsOiS683gRAqV71ZZfPsGViKneSL
3nW2j4/uBe/JK0rBXd7LUO3++3f/Q9f0xRjy00mflb+Q2R1+/47lA7l+ZIKMdXRY
EwfjIhU+xeCoOoDIA66KgfcC8rOMgQMZKT7sjspxfWU=
`pragma protect end_protected
