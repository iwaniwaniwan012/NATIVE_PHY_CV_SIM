`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HQF9zP7Ep+qkIMg7pbAZhJcVgrI6LMevoOIRl3Cpv58DKhynRP3A+SfEc7dBdD6t
eVqismrvgPbRkp8QdZ3JjO61pV1GiGqO+wUf0QC3+XawUBsMcBVhYDvsnr2CVsPv
IaT1sCGLiRPgKLv8kz8/+QtyJv6lD52oxzaObvcV53Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7536)
wNOS9zbOXUkrCHKivKxPc6z/5MTxTNzU8jPB+9an7rDOVPAZxopFef46pbYKqG2V
pP/xjHeMo0sEDu4bGKsD6Y7utPn8fvc06IuHEUQ1YUVXapkcPNud9YioruIYP5iM
TSswwsjKC1y9jSsviUdPD32FqIfiQmhvjv5wbzM0rqzd6cg91MOXAt/xlth+tIkS
XF4vfB6MP45Og6N0w4bzj3WRkVMym+XwQBTAgmthi8BYjz/hAkA2xFgGd7lahlwh
EMJVPj4GkLhRZYOWXMeFGEGePL72sZWEKOSniqxY9f7GJ8dDPt8Ooxfe8lUrDkQ7
2D8XBN94gnyvh6AYhMnTK6GBLte7mnN4PB5Eq1a1FzUcIf8lYU5pbaSsy7MqOjs0
7mUKyBRhgXv1Cta7JZ5/MIpFDKOLgqE3sNc5GpsU1rFCzGXDIpQRJnxVK+ErBM2A
Y+Nr/n4D9fOQPnrimb3/4zUTLK2dG3IMr+rJ/T306T36ay3UT0aJEB2y2zybG165
oeowl4JpPBcy5mgbCVOCFHvzYzdH+26UkUmwB4ZiUxX2o1Dz7IJZLAdVJnDYs115
rNiwj2C7stH+S3bnR5Qh1jHyAZjHQi25aQj/uGu4bI40swXxUH6892uiQeq9xVj4
wPAq8hTVU9gyq7kdl+ELmZzPNiEIeGt2R/Nveg6nkKMG/iqChnPA4ULhfO+XjrTF
HlpeI7yeTcj0FiX5KshomrjeQTmQLQQvJzU7eebXaFdOPIJmYSLRKT8IocRRQhMy
XNmhjJSbtVOuXRwJp3kByj4cwqIqdCeB3Gf902lP/odNZMuUrkefQYOZnmWb1h4v
6GHtM6pzTkTN5AWD+f+4haZiu66iopIoI0Odon7vaKSDbzGRPAPCJ8m6rIoJmnQr
kIWoLC28DRorsweHQIbNgIcp/dIhUQj8GFAJfZBVtG8S8gfBhopsQ5ijb5pABgv4
oeWGf4kdhgG2hu9R7y+etrW9ZmgCdSXxo1FNVwJj4YHjzpnqhcgnuhOXEa1LBQCz
Mh1aiVdXZgvg8Q8aD8vYYWir078t0/ilPTXO1k/GURacpk1zlmO7jsHHev1W+e4S
a0iBWbtu3Nkv2rmjxrKiSe8BWApfCNPFNb+3JrsqZaRiwbW0+kwmCBPwEdBntxiu
U1YLkzswvcp6WdEP4XJKzzFNuAXlCMgLsa6p4JdMkgtU0y2pP4Cd6HEIi0LPQaQ8
RNThunKOLG5DOCVE21dk+t5Q52D9/BhayZ50q0oSR21n39AK9od2h3EkEkVmT9eB
ke4YBmx0zKPqVbDLPOJ9v5l6kFf/fztw8IIKoK1GyZJyI8+Ta9Q0YKIR3m+Sgo2+
PN1BRUYmL75zDze8y3zAIsQsQHraoQvl+sjo5i3t5IKlqkOdgIrFPrUCMAqLCp2Y
EhPKvNUHLt6hLzJM0S/9T0K6mGyhR9OtTfBWHJ7Y1EO8+jr5sajCt/SOBydNv3UI
99hF/RPJJ1wUmfiofyip2G1e7JPeeLrHagx7JL8Jl2wNRRDeGBlotAQz1ODwL/ml
1WFeJ2bQGIDlg+aPdO93xZEPSQiwt2/UDtsCo6zdxOQZLv9mBojAXBS3ueZTKhpl
rQAVkxlICZJA5fzrSlTkCexs7KZDHk6PiGYGc9GgkuooCcd81YfkLNQOwmLFVOwD
/x1fHpFwBXie/mBpfV5yzV4uqFsQdj46hFOiZ7cgXpeIYAE1FPU5vpBoewXK6FXi
dujzO9VJjqqYMOTgx/JH5p1r3JfLfFRqLvdQ2F9teVep4Tjr2oqsTTjyT6lCYHfH
aYqThFbL9Dqv5TpD5/u/KvY9Eo1eWmObfN8BXA7WCKqxGInoN0RUaUOklXkNKG0A
LgpMdbz3cO7WqUzEGO11K7u3EI29smc6IEQMyhOoqQvtEKJivc6UrRJD8ySJI2IA
WweCMJdL4tYNYCY5RZDpQqkViIOs5UzVpRdputoIwlzocFofY45kgcKl4DfaevOY
+D+jWtBPHBqYhBbeIrWeSYou71NhzKYrKzt3taC4iwcmC0X6QMQyCO0OBIFJxW7j
0LnKtxXktulkMJsVbjNElTGvSiVIgY0Ax5AwX8C/hnY8nftM+rT+fl4B1d7QI5yz
i4+96jt0nT3Bio8VwrVxZXvVlxGcWbPp7BTXWXO4hOKDG6lgoSyjcvOouyHqvOE0
Zlzt006i9RMXCIaLUEpT5SvXkOXgjsE+g1+jJCS+bexnAq015u4hIb2lTLZ6aEZ8
20VPyZ919kyZ7t/PTg8VUQX0OUHwmzZvCZZkv2mI4nrp1Xhd8B+eh1b4T9cdXebu
R29K2bKRAUj/uGHW53dhP3QwYdFin4sWcgo8KACNoK4w9iolOEdu9FxUFBTAslSN
iuXP+xNX/bfy1pfBk19JMF3VsMkUyxaL0HXCxU7Gw1ApFB/aWT5yAMy4u5OhXo64
0Di5t+TkQ5ftdj+hfZT17NfUZmYVnLzqw2AZwGzDjTPPoxI0JvoKtuuoNRz+v7Ul
C9+W9l1bbZ4S58YK1/zeY6JqJObclhIE9hb5MxZs3VnwL6VDdHZ3JaxFphRgUmTG
uSVSkiaTSjVIJVinTEoylDT7LYbaJxeMjt3nqkDcPHumx4YwI09G3O4deeW9fpLO
6ZjUItcnF/7bHgm9KuAFtfOFZMJklIo7NsI725nopjer9yK6w+Kd/ts7AVvaKZLL
lbgGkWFN7aqzvbVFh8AluQIDs/ciqvXDpTFArcD/QKRDNlSN3lavMYnt1ucZ6wrs
uOgzHo2556E9N3vZLxTMXIJYCQwyzq/nqt7PNUCkFvinApniwq8Ly/NFCy1A34Q6
nBjLLyIcy4I9JWS54Avj/j6Y9GvPG/o7UqpcDy/X8LqJdvFBjEoxQGjBNrRYYVzU
DblPXfDBrO1KnXfrv/XnHjDN0VqyC7B93RhhDJJUmlEO61BqBW3rsCOvsMKuJyK2
IyXaTYqrBriUhGEYTH8/zuWqFDOTP2a6wMvBWyX6EaAFT6h/XdApJWFyhC2icMp2
B+zueS+TMI4bih6IlMGU5caKHFkEuMvR5YLTmlpQi6l1uLMOCGSe+9RVefsVysDV
JhrD6HKXatQFKOS8DM9Jf3lTEWf5NYFknA/jpA3lMZxiEVLKRtF3JYPTbRefnoLL
vl3pBqPVn5sdxmSEwA1qAphlebMWQAW+VyPM+xJAUr6UORf75c4Rq1frrUGkIWl0
bIUgZUm2PIImK4CF9OMSIuAgylCHfCmgfgNRDNv3ZS1K19wrJm/Nt09iAdDublHH
CY9jCAkd2g5+bUrEa2+k1AlbLu1inyB2Y7cm75KxB1LTKb0lkjEg0JdX/oGkmsrU
/auVzdHC/XsPWVbYOjBEUgVLG7Rvw0s/cr1K8OIXfsYDn9xs1dAeM4kxziQZi4H0
THlSFek5g9azC14OQ+1zal+Ut3J3PxqlDDcfUgZD5VZRMjqf/jxLczRGC+ic8pW0
hllS0GQoOVegrVYpCP2I+Icsu4G701tNp2NGFU69a54936Vr8WD2XaVamve/1OpZ
qWfPvzv0uCvlZPOy12DsJO4r5m4b6+AfYdgN3R2k2x7nqz+Ya8S0wI3DxNV0+sv+
UYtsHUohaI+abX+eoZ0qkWkccEz+ZDo6OzoTle6w6bpLy/vJ5GmjbGso5A9ZXOk1
HeSeoiK8JMbNPKuA0szyG9JEhZ2yWlhbX+luikskpj12k/ox2YCapClbwSaLstuK
jT2KEdS2P5oAOxxp/IPEA4cY7VSRk93F0MueX+ENPLw6NCJInQjwCn5LRDBfcx1e
p3iqO26CQHNtuySfr2+O5RLTLCT69WhxmtMrd2iyx3s3MdynPsHKmEFjM5rkpQWX
ic1Wbxt9docH5MbNjyaUsZ/df47LaJXm3lKJGXyGwQxWIjWGeqUr0JOhGsxT4xQV
oy5roPCYTrZwVUTc80c6UBP6Ko82olDp0giF9nW1uOuwj9eS9u41LpfoB4Y24YaB
dTZIzfMcYLB0Iaq6SAGXP2SHZNiuArXvKmwcEjUmAWMgQo5ZCWdraZClGB24XZpb
Txl7EHzA2qI9JdQErScLb991pNLEeLDyyWDjbJX+M7cQaF4Kx1xV5g03pHX2wnQX
qoSa8+YmcT0Zu/mwpVu14QZ6CKjH3hMaquGS5x1i7ggiLkJ7E0hYLA6SL8sH0RVU
FdWbGBxTj7WRFPY2u/AiVMrBT2EeNUiuL92IZNlTwebnHQ+5qtWUiOQqOV2FjwRl
ASWwu/K96zdpgodrrDCaNj1qG2jJVW4v3oHKBNfr6H3ez99fqEKWcIe0EoIEFezd
iLCCY2FDd6D8t0bcoAWUTYe1wBpPVw0ogTKYX+tzcXE7BemegLe7OxBR8bflVHja
TwoZbe6nOpsUM4Gal6QXIb0+zq/x00sbg1K+Ff8yEQ1dNjrxrSpYlZs1Z3Fjl98a
EdUIexLGfVCZafb61t0xbmmthZCxxlk0I6kLnxSxoKlyQTCUVvH86eopg5MXMBkg
JFsZ7K8c75N5iE6MKyqVGO4OzAdASSkgtrlAvjavvyL+Uix4QPqmxAyNxPVmVSuJ
oVUXKoSzr4YxokPDWoZHmEIAvS1bvGC5roIsVaB7qSQU+hlgx3IfqKn1YHc5kpWw
lO/FHU4JJaYGZMFyfBGrc06XyGBuHoHugUujf942UpAkNUHY7Gb3zbDsWaXVUhPt
EfNNLGnJ2gH3entSpf6FBFrNpMWGYRYA922vQd3W8IJieA5DyOJdCzqGOnQ6e7Kd
hEy1XYw1Wcu9VJRYwOqv89JSIJ/qme6T+fmNxwmlKkaWOTd9LZqnztjd/lxlBESq
gC6JghhWINPta/HOgNhiw2vIKc8Ui6oI3RT0TaU3Qt7BvW5clu+E0trAsl0KHpdd
EkcdjAYkaT6p54d0KX76cQOoWvs1nD2lofrGLYjZ9fcsxdLlmsfq21xEdWrZKy01
VK/wvbYjAy6cMWRmHRHymNvKLGHaLLdC5BO6zls8+FXWzjl0nrsAbBRsuxmNrQgv
XJG1JI+AgMmsu134xC3RN1CIxcJxzq7oTbHfWX0uZBRm3qy7woqBTqoUtwsGDjWT
EHHpjaSh9CxuHBSK5XDN6p3N3+g+xwz4X6OwuJb0qKDVXuMPtdKLQUoEwqMM2wzx
lQJqaXxq4zDR6B1DOymKwg7s7dKlR37o+JZFdq42xht29Y4Y4hRZfmUM7RDpfLcs
lb+eb/6Sx4xg/ymn9WvGcJC4n1aYR+XVRZxk/qbrKyJlatzhYefmNrIAhpgJCnLv
3FWrHRgmpKhKpYxWhQsTjpaSjgpJNYrzwOngYvPcbS11WYY4qSoIxtFr85/CjW+C
b7gonq3MhaLih5zUI3STqSvPcZlyH4k0ie6AjsDNv9N0FYzQcfpu7YMkrc/pA4v2
LBmpfnb8VhZ1j8rTSR99zWp5NQmZuNjOtS7olyyIsfZzF9U2GQo/x+iF05GNyzyU
Z6QILk2nSxf6pMGszcVsL1pG3Q5QNLPsaDn3FR141JyFTIUhmKZxA/1/vt/504PS
N8bcKj8fUpTIZZ0woMDcbI1O7fAJpAmBIsUcPsloNYMk5J0dOve6oNqEW1xKHruf
dU41pXLcNjhkkQSTOw/rNpIzeroxe73gx1Dn1Rsf/ns25UAKD6X4/nOfWpyDtwOF
AREYDVjW6wq3Xtd+t4A13ove/jckQfvHykEq5g/zRDFZ+Q4CxHluRwsZZ4a37IY5
4iIO1OrU2O3RruqDn8M76poorxGcAgbL90dVE1rOA74MXo/WLxiQgbaYDGha2Umd
xSynZaT7q685UNiTId2XIz2kk68mdHNBw/wFu8nUuckB4Kv56uiOuan6FyRuotL4
KYvQ52qnruveQAXxb/SuxymcByRc2Q7J82KPfr/sk32RwXoifddl7Y9vHdresd/C
643j/isYGYKvxdTbymqNQUcNmE59xy1JQI/mNjHsEqqLCZWpsBTaZh1w7BuWZbcO
ShSc6eu9GILQr7DibWt0KXH7xfCFI1SoIwdzhXvqmi3ZMkVQe851CHO+le/x6QOq
BNVn4co6Uoiem86cwkLpUgqFiB1Nk+2Sfubb/Imq8Kad6HJTSYxNOQeQJlpZzKCo
8P3tmZjRmgpfFgji39rTbivUTkXznTHGeD+D8D8bEWalv81mdx+blG2FqMj+TNX/
wdWpPKsNvwkR73l3GpiVmCFu9CEy9WpIlq3rbXVgS5K/xn3wEI2rDZ/Fis+EHvH1
uB1IJ7zBgAzgHUur7SM3pp9r9HSNFr/7ShPJcC82F7Ksozkca7DOMQIHGrv/aHVb
dwoa+GvZ+sDunooM0RRJpwRc9JNbUim4Gx1p3pkeTIUrNQniKNNHv0Ra/eu/MU6e
JNf31af2b35zLPFSFAMsYCmESQ6xiXEYPF3UPERBnrR7S485rR9foypGYVCTZHFS
oopEORk+C5pwjpcdrLYF7wtxs7uY+HetOA0Sy2ZDxbWfAeQRSZlEtEBefdwHniGp
JY5ae2jKVSqf6kQ04Sw0kgS/A9IRBsdoDwz44+hr8o9ZNw2+2b+Sz2tHSVKVJIJv
NbNjYEpFH3UAiObSWkVOII/alU3Lu5eXH23FTBbWhR+IwlSKJTR5GEKqjk9WCEIE
XU0kcrVZVvp6UPAoRBsjVtaocKf4Ui6762ibpO+D664sWSOy0Hvs++tqqSkvTghN
arC+7kPbG916EvasTZSDoD9pqr7BL5tEnONj8lPzEvT1zHgQfKR8/pmCBnXuengv
2IHN9Yyb6OC37+/2Bv3JS7uavNwr7gNntWbQmzqAwPQOX4TzYiTsHiMnQY852lvn
7sjZPRG1sXYBeaX5UrETZNkNRuBJhErdqOVQG3YKc5pejpdDzbcVunzKo8APlEXW
K+t2NA9lprg3sLm0RkCwnhe3jcqD+1H2FwlqiFSdvKUTazLUan8l+X23JxoBH1aZ
Ns+CsmGhvSY4eeIs388XUi3WOXy1qGQ6yRYSLiTwR3p4SNPtZNqDmuQErSpR9jMK
6mnEjggGwocaKRTqnnNFVeK5CQ4ZTTO/BNiq7fJnvBesSsn4o0Ye6NF79QJRXM/+
O0SQG+Pi494l1SZnB4o5exTVlsYAONORbgTCfIcmhWjTvi5eJrcBX+FHZZouYlDU
rE9odWHjKndyM8j8s3CLz1flUExgMTf5iHyAR0WUFvkvPpIXqwrNv/hsK6F6R54U
DAflar3VouUxOLVPfhafyVEKlsjP0sB2HuXHJ8/a0QiQDJbU6ks9qCBErhbtB0vw
cTKL51yt/fgT4fLJJmFeXmjUFmdEnlZG76QGN796tneaPCxXs6Be5VQU+VSjPmhP
MN0YYDFShmxlc9Alm+sX9s8/1PruR1mT8vcpWgAjnZFPzbcLDZCb0iyHbUUk8PqY
KP0sQobDc/j9rgbJslFRVblOyqyKvUXhOK/IhFvTnIB3dRDoIepAqeWx9nCAZf7v
oXiDwVltWBPLfKZySuQFH8OP8kyim2r4JBUJRsCKOAOkJ2YkANwDJHag6+VlK7z0
PLYAD4HgodcBNQuQfidO7pg3C3is+fwT0Zb/d3rQtWrYsmNl6kv9SbDql3S4dRHW
VbrievSLzbZmylprUJr4m8SZFAVnEOxV186RPAZ8tuiB9v6IaK3E3X4tMTFIZ1Oz
GUYh3oRyl8GjC4czV40erK5725WBry/nt7wEMFg1TPEgEEmRjE0QCkCxYzzVTFO6
K8kxJZVc5PHnyWJUOcKOhbLVsBGEwwAqh5O8Lo9XlD6MDt01Y5tCFTIhg1GHhrzp
rQkbFmQC3y6Dkoap8PruK+IJ3NmKsHyaHiDQEQqmQ4m6Klonmexo/rUvVTt+lSV6
Phz+J2owxpDTHW9oB6HOaDvMDxZLQaFeLuJjzsXW499bM/XtM1OU0ILapy4UKFXI
HkKl6M49Q58kgVpOMPekwEh2yf9ZPGRDJm3nEdAA4pFCWkkZfvhyvXXCkPSX7rlY
ejE7wmU3AwTH4jbmz66PRFDybz+bp5siI/UJsqIrmUzv5rzyHB9qK1ju3ALFe3Lw
tYbczAZlwBuwi0fQfYJmQNFBJcHFjrCu76GHo+hboEL11Ug8oWjmLmzNaeYeiF+G
iYRrwGSkVPaZb2JcTRtNWPUmGuXxd9SfHPUCal1zVglW90jBlJ9xZ0YDle7irr4T
9KIDCNEWyx12Po/R8bZbLwcdMc8o7Zzc+RawVsXexzVYWutSRGHZT/GdSvYR6+Rf
BshEreVEJv5DbK6esTGOp2BeBxgQ/5exKIwn/fegIoDTwteXI9xtGJNETzQa8Bz9
Z5EUPe/XHWM31WRwcXgqRAlTMSkWWVslx5iGoJ1xEEg64KV6jl9kK0VGqCe1z56y
AQjCU3aVgnL5/skNUb4W6b6o7fwjmOvGiUXm9ooHauHlVUeCh+YhDH4ANRs5aK1m
eDP4EzZ5G25GJK1Jvog3HX0Zsm6BcMlMaj0sBfacD2nq0fOiIh8wdsey5zz905R0
rO8+7ON0/6F/vTKlb92aA/x+08N1QKRvnhvUhzrFRRoRYq4rGcagtZezKe/7O9iW
4rYfVqKmVS0C5qogtlkRXW0B6A+prk6y4UM+zGotttUOPXT3nI3Co2DYBz5NPTPT
+M9zmcT7doE7eSQ8kuKAH+lwG7KR1DQxZYKgyxzH4ENmAQwLu4qct1kNgJ5w1OYx
PRYw3N+Hg6NcyTYieqYmRXRSU42p/G5DlFgANZ0txS9anwgAlDMVlXxOlQgfzJdc
KIZtR30B/UHfmO9/c4zIgSbRBqAWz/Gn40ci3UA0sX63Y3JsT/4/oIpAiK8kaVmx
vO3pdDeUx/hSW65SpvrhhA64SCwNemRDpovSZ31CmcHOlbXxE6f3OBRxPmVTJPHt
ehikfcTGdAKk3A46BM9GBARKGCQ2xPrESOzcGVXbvTYCdRVigcsx2ZEL/zFtgvY3
Lpv+pByJ9BfUB+aU8PZ6nlZMYz9Fl+Jf8ikLa8MNoiz2gT8glUqEGpl+4f8ci2+j
ZX/hqHFs21/0+3/mHreA5TIpPpc6CwrVRJ/EnRnF4AQg68LDgjoXJblPdHKzdQnx
kr7LMgo6i9jWM1h4Uvb5fptEVb4XsCgMQ/EU7UqqjGOb7SY7yV/PTuTZP3zbbRXB
gFOS7pawbIO6ftBy8HhNWs7MosIvQ3Kvinmzs+8vyvkomO/caLp50SrV7aww7UG8
L1dF3QpV8Ao2BetixvAWzHW5913NNM4XjOJU7BpEplh4t2d4m1ABbX1rEXuvxQKC
C1fPZAJiwXXiRAG2jOE9QWyoAVGC22G/BCJk8Kqg0X5A6AXUoVmRgcd3Q4M/8xGX
755M9wxgmKfXKDA3U8NS+vKuR7soqeeejdwg/fmod7XOUjmOh9f/hqiVkTt9gtXU
bM+WTMk9PYkUrvPo+aUN0dxvKsfI6zwYTpBg46YLMYbklMT4j56CcEsgv0ha2B5j
PnX4sWUv9wX+tsUEzAOHt423kSVoYw6ySiTKyfi+8VKOrW+yZ+GGHyI782hek3wO
EvgECP5d65GH0uJln8FATDZ3hDPNiNNdycIIg4poOxHnMtF84FDEX8uS8hUn+3/I
fsQSkQ1TdX0dXCpLMc0eGYzyN6TL38J3Jq71aOaROH7M4HVD9URT1TZ0QekM1Vsq
zXsY3rxAeyJMbSoLl0crufzhZ0J8ivV4WOea62I1mUBphGSJKKNikz3yEdKriOhV
WkwqbKkLPc27tNh35LT6R0IEdyALNkrvAlqP5V2XMVlY19DaLDWoyKfMm9BrKG4M
E/BFIV86686HA16Nzm7FwrWZ+3CL+bSQ76N86rf2S/2UjeDjs2xG6o+llDiKWJ+u
rQ41gKK/yjG7VK27Xrt+/F8KM1/cn4+dGkNsmDt0EfnZY3yVjlMsori3MlP6RyGb
pOrAht0vaw1W5V3QXosJPywA1CPZIhEhHkYBjiQwETnzQKbqRcjHE2w8I+kNLopL
8Ynnq7bF3eq0DNavdJEBVvmCzCA9kHLC2ROiKursK3P/nHXMtJM1srEMnms7d84k
YkGPdvsjrhE+IiS7hdxDKHXpwi0/TLbtZMy/ZPmhYV7puRmkpyo8FyUPEV3LnKnA
`pragma protect end_protected
