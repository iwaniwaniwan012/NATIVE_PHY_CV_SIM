`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
O3jRh6ONPB+8D4pYByQCBdxszunxnq9I7OzJrUulYNeeTzHdA/hmADpXKvBKmVsW
uckPRDJ1qH0+x3Ti4uE9LvqCrwbnlsC6mP9YXbriiq7De0Jy32CoHMTtpMC74g5N
Fe7EEbXZBvXvnh4WYs2FqlDV4p9xcLoqVXWGsHJoRvQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9632)
Mkh8YxHWZ3inc6nQI2DQ1q4AU+0ac61MKh2CQ8mII1smz6q16gWlDm5eSGlbAwjd
oEYzqzBVXthU1issgbakrhIq3a/J3G0xlGaIunZErWGKRKJwjJ9TdKMRQNK4ckCq
THIDCvRUa83E2YF0BS8gXpQw144Y2WCIdRLOpIQK96msYbQ78JHiS/q6L/P20eWP
EwMMRY641gxSWPPyVVqvCH7tzqJN/TbLp5rMi2rNaE39gyLCG+uk1m5RTjMk1ciV
eNNhrnE4pYUfnCFWAludmt6boWdAn+jpN7juUiBH1l80hOIlBVaW5ahr5/kfXNHh
63N0seMKFQOjJiy/PL+cb5jhvWttOrJDBYo7g2acrdWeDw1ANrOcsr0CKsBDznnl
VnC4B0vgk9jw9tKb9PnovAo7Y4IvxoTGVXwPlQ19Yq6d+OqQss1Y8cNY4LCWyxS3
H3zAmnA2h6gpvuC0Ur/zgifEh4ymfchAlQmS5XLktgMTUTzwiFq84ezY4kAn2FTg
nBXBvadbbHtLeKglpajhA2Ytoo3bzCqTVISJ5rjK8qlxpoZBvtMSFWEvnkArudD3
eUmT5NeFeeGSjM76DVwWjUe0GLtrLxxo0OD01UXaXvIa8+TOYTF8MxOfQeTVQ6EA
9SxAcehxOyI6Lhi1N9pFu1fTtmwrpcEAdhkrkbRxsSUsDPpidsbrsIc1YVn6NgVh
uSZNwh0hJy7vFGeUBVfli4+jYQTPeH9q9a7dtEgwhBkqmgFM1mYREfYzalVPzRFo
imnxEoIm20BexcaHtIKwyVkLjIoSiFNibjFJYC4dmQC1x2lToCHHRiFFCb/GeAw5
DtTBZIaV1FbjNdDR9Ckgobw8XufziCZg3NJJSMwcuIWLJIFKy8kqJBTfXLbojr6U
64GnKmuHywRFPYT26DcaCkVYJcUzoY9Bp1CH2IhvEn/BxAnEZDdX5R2Ka/PfidgW
2Fb118XIcNsH59P/9kbhCwtX9x5/U+7ha0zp3PrpZkUC/C9VGy59T37D+L0yodFD
mL/92pkooSIXEAlfZtSBkXEWYk78R3ssh3OLxK7CeR7HY5uy1owgCCcmb13c77Mq
xWv+KTtAzy9TIDRhmLWLGRGmx9fwyF4c9vVewP0I7qLcNOrrTuQMBpPXbaVRYgSs
i5prYZnMQPB0f9SpyY+vL5f8ipJqpYYVttbTSIJRKasbdztuP6WF7QrWO0b/bkcv
gXH5unRk6/9rQ8VHNetYEQ6nFvCH7GOQ9tTq8SYty8cf/i9DZDvLx+E9TWSdr2j9
OtzDpAYk2M0xvfNdptsH2HqvdhetrlOBRakJknQElS8D3NZvf71rgq7vZQQEbiU8
Jnry81DviWcv3V5tqS/gqGF2F7q4VCk7WIGadw/Cf0fbAokvIxtoVs2hgJoJmnvx
MwtjXgl6a1WERGo6zHkZrkW8sNKLACCdT+7EAxwdOYWH/QmEyvIt9eT8Ve49Ynhi
/HJRf0tJsggLCiG+f8qj/0hTeslI+eCjv18Jr9gjuKcQEgNQNksAve7EEykg+ckV
M7Kc+xjvAfJYkQ+37dKnWL3H64+n3olGCbeFlzvTFDAF4i4xTq2ijB6lenS8USGI
RtLt4Ys/CcA2x7EmMeIrUMeUABoM44w4J9EjlF179C+sssC6YqX7Z3AY2UxQ9A6E
ziWMFnu0VuVdyw+CbaaFi0uEu5lzzPWq5qOBcdesrLRN3H1RGnjk0HCQ86ooCg0s
y8iWlE/U0hS5a9xTSlOFBOzIl2QGu64MAWZ64k4DxLlynr53gzo2szqxT9QYi9uD
ZsNxulzQWNLWOl71POMoYQv8j9AamNglo1vszIxmL1lB0Fu6zLhtMfEbiyzQ5cdX
92sIwozG0f6WQ1OKpY5Km/Zz4vOSdjlyKiK8lOgqR5WitWoIss98lHbuFHYVIYYq
YSm17HCL+G526B5fXQF/gOYpJ4o4H51+xFaaRX1l1ROzsLyw+kXMSazUn4UoXI1E
EBQxlRAedH2kPOVFHpSQ0C2NXisIVdpjjMfDbC9aeCYu651/NYrBtykZSiVQ1BRg
b6aPCYlBxTSh/tM6XgNx/W47sLEilhZYp3llZ8/Pl0kNY07JXEDl02RmDT4z5SqJ
ra1lCpB1bZ3akhPt31sRBNqp22kgcbKyjNLu3jqsBrmyRLlSfkwNujg4MznVIapC
UdJl9Y4n6RgWWH1T7QXjnqWGhaCqfip6QO4sNlyR6w2hNdz+8D/wJKF8hxBRslCl
AhexjiYbAP2DIlgB0DAHc7qTP5eQRw8WTMjkJN2jaoMu/pC2GYzt7GwmYWGNUJ0i
zXgLp+/eaucCgG85tJTQu0mZBoPO0qfrQJQ3KL1GrPJdZ9BeYqpf1CRHxoltIbtc
lvhKjQdju5Szyv3w7vUl0Hp3eKXjsL9Q1zZhPNA0Ywf6hWeTiJwBv6BLzqUo4JoF
LlyT3P1wO+4sCLGDonifqd/to/Wq1aRoHpsbq4ZM1Y9+Y7+JVdLqUFKapqkFjHYh
mX6QIDvr8FJyhEr1HKNZ7bh93s0GpRXrzfS01tBuvHNb/BKpoUQcUYV/TMzHyEal
npRVyKZ1FDYMQQLvaGhVt5ZBrqEtcyGSlGH/TWwmukeoY52hNOiFn+ByicnMF6BP
t8iaY46rX5f1YI4Y4DzNZ6KFUcGlE1w5BHcn/4VzOYCuOPmoRWChcfipZwHfQr0a
RwOHuc8fC7OlTYCL7y42GUr1LTmTbt0rYCFqymOQ7fEu79563bOiRX/VYz0y/k1V
Snvx7Je/hjsp9lfWUlEXqvvRBe8wcluRRM7upMh3CFMDmQC4egog2AXz0fZkNsPR
41pC4Jpdee+Xnj0NAmtT3EdX/a8ane8QjE5XSYIOO6arZ/bTUAYEKtMGUsgQjnIl
Zz5PsRFA/7nUi2zCsgtC2mG/z5kR4/gyS28EewzdovW+0pnLp7uG2DUwugGDkZ0u
lIWXsn3vyT3261+6AI5tqP0UVeR90res7RNk5Hz54v9+c0AgDbxuiRHnv2xQwk5P
4LwIEAuqBQrTUR/RuNU9hQYGigjsySHjTEzizI8kgNwlsgdOu64Eyb4+FjMeJM+U
uOES/R1reTmxjoadKJMe4KwcZo26f+zcLhyVXBgXmuVe6OZ8cwF/HwMjSXKRbKb6
B/Fe3HafHgwGHsuTqBRXBp8N+gsi2vBUsMqROnywlpU60DzbEWV8/klK7wYVGc/x
Mjx0QDpOBWrSMj+YnBccaPaBhIcEZBQPnFnva5g074O83v9FkU5ElYcj8hDL+0Pm
r6Yol4OwKIoR4ISRJu1v7NNFylI4PQh7AtGuckn07NliFCWqsiC74I5w4I1Aquqn
1XyiO2LtFsF+dtfr11+SI/4tIX5i9LsfEuwOUGe5D8Lb9dPv/6Ofmn8w/kn4d9GH
9bKJqdUKFMP1TuXdxMSiUNKwUlMVZr3yLilM/qg4fwMxL+D9irlb5SgaXDuIltXJ
pIJNHx9jk9l9u6vpT3SRfBBSIU9Yd2HSNfwlN2C1EbFUXwsT9HujzGSKcZwM3FC9
ETRM4OjAgYXU8NIrGTCf26NRfTRFY81purLgcWa6SwCX6uZ6NXIiJv9ED3hQEEXx
uWLZRDQWNBrMQ0c5vS9bKoRYEjbvH8vsl/38ufK/C5NTeLo8ABcnA07mukGT9VSo
zL0ibHug2SnXGi5tTYnlakN9MBR2I2RN0LtL+wqh74NdAZWbpphABJtzQbuHy+Lb
Dzsg7Y1h918B+lAqkOKwWhStS6IC6XnxP7piCoKbn5pQnQuwcfiM1XhWNRjDOIDo
gJHUnR7Ja+n1h2R9DVSOpLCTJkZziLX76ZlP9IQMYvRY9Kjxz7lgtYcR+fbJMmx/
B+zo949As/tfcXypLvkwcjW926xDcZklfiSTmyJLkRtUUtFyb41qBaHhRM7cTCPm
/6DNprBhbWWWoMXwmGBXvnSWgiJkxcrxxbu0RkQkxEDpxDj2FoSD+wV0MAJfNw1J
TlrjBuXcVaNDZ4lY6PYtGgt/RcG58w0notpbaljSTS2XFD9HMaBw+16IiuUjlFyC
ER6GR8uAO1wlmk19XCayKhQtpuwUm2edBmNzCA8F5D+8EIJ1WucvvZ8BzaXww5kw
UgqPLwdb2BCVX5pqKnFXNw3oKFp2KSEAvZ54bIofDa32j73lIAOjkt/2m6jc4xKH
xOcMQoTu88PvT3TlyxcbbULlwWIelQUETqvVjYrcAnE7ot0mpKwH+LkTpXQ3D3GX
VqbvGn/NCiXwk+REUlhBPd4L7nykC0nK9L1TClZBU2g2e+Gm7dNXstEwwKn4c0DJ
QVbcEsG9alCViN9fAkpj57RWIiAcFuQt5eTFgarIAc17i4YePrNnDfmhaoryGtHm
kihiTBlLpXo1M0gxp/ZN339iTsu0TP2DExS6vwFhvYyxSapKUNrqk2KIPoCuCYK9
3RSuFpPthQu2lkgKg/5rLjppbOdmCT6x5v3DbxL2NEELzOspYTnJ8KNWKfhhqYxc
MzQAB7Y1ZW7ZOFhYc9oiyrIuwtNyJ7d3SNAgpotEjCyNHFzB1zVYQXy4Xx7Al2sS
jw0HGRepKTCN1kJk9FQWSmrnRpQyHfzDamkjVMtCXqk4WwD7kYk2D6b3Mn8eCLTn
kC1l0Sx24EQf8uNy80wpA9DDHDJUlx0OU2yHl9lBUW1m4x/2s9MfNNkjUSwxoSRP
ysA8cCiFc3VMCnkMkGpRySQrw1issTxgbtPOdXRXlitCojdEvexi34O1GMDKswcW
mkG0wZ3W/ItJEHFBB6lVrRkhV1Ap2SGvkwInfkMg8ogR9t+B48bfS8Yq/7SxhLhv
YqxGyK+fvr0BioAqwfax/PPY2mfdzaa/qK7Aoee3FaMJXa/tiakbljhFXUPEQftj
goGn4cxRnC6ckUFrcA2JCb/Fufh6E7Rxa6dD8dkHG1W1MZQpqoSEfAME3m774Kbo
rV3KBMmZ4SJNJpwfims+yy9aQFFbV3abRMG8FmiNbKn7MP3AIOZnH1J5tL/egk+P
5yWOn4dsJHsabb1bCkQnkp29Jnh0ow2AWlIkrkG3mHoTp6/uFkCpWRuwzpGVp8om
gvlDmK87aWGbANoyTxrO7ME52VbijSj9vFR7fH6koXohUxKzpxXMSD6HTRoIOiZP
HFE0mQajuZR4SLswHBLekKdVneYn/ur2Dz7AHm0Kue2m6rRa8pxSQvgSVqTORIYV
Gs3jMHQgIP8InBeEILBjw/KXxBkWx+6HXBYo9fvojOFpmxyt96Fmim7bWgs7n8JF
3YyIB+6+Sf/BDWhr6fDtN30OQckLl3zsgA8hzQOHLTkNGiE0zvCeZs+9LWAdg+Il
9iZNGy//i8OrSrSuYvf7/q/YRANOhvyj5ovRU++Or3S/uIhsA++HHzlA3OHQh9Ed
9SyuLs1lFCfK0LybmM9ZkzaRUf2xnmQ/wNDmHfH1CO1xQ/DUQPfvpHCBjCSmhMAN
EKuZtnTHpjr+IuYivcz+B7nvsNUPDPB5ooqBX6OZw5hlCUg0ugdwqw9ey6kdoTm1
VDFnJS0oK66gImi65xIj4/VNfaSCHx7XQZTGs8xDkVa0Ot7sJ8CDGeBkEEyIE6/q
GuKSG3sjArO29mhkQK9rNq8RTK4CSphJwk3AZNF/E2ekJidl31cySsWMW7dZvIfn
7odwQhFTpU++ZfW/WoWQXU1eiQkhSUjc44/TAweYHMGO21oOPx5EKuXeMqA0fMZ+
fk5AlpKwQFB4aWWmFe4OT63bB9QHPmD4nUFg3Paz1yQEskHetrd9N/iSeJn9mqJg
VJJlgV2g46QQmpGi+OOwTDWCuMFbLh26NzxHDTSvV2mkuo+3QuQsdzYJe0A/TTPc
AkI1n8HBWAwB3YXSII8Wr7EVEzApLj8OS/8y6uJ7wU46p/IymLsefwkSsLsmB+f/
hKatkxr2NZ4EtJcWADUSP1hXt5YDX096GU5pOZRKbz/rz+55eLwOgZC/v+KfJHMe
EW7W1rux04VkyaCkf8hAvi35uhboGYL8e3jGFJTXcxmnx0HMfGBt0vMKKU5sDPrA
8sYnlUTG8HQEy15rhICgC+eKsOdPXrPatEVKFfBJT09whpsoZ/GJdGO1MKC2wj/M
2k4KjU0zPIN7iIPMbhbC7ce7drDeBLk9MzHXsxTXCKEV1SM0vOaE6FBvkIHXjUHf
WDGYgYFGXTGLFFf6RU+8BPG8wmMlBf6bNDsaqRD6LoKR951JQrh3VV0DOdLMekhA
K2mkz6RJ+ZyKLOqAyfvJMniBwVC3ZeSRYrvi8kVdShVQw8lzwIzwDKvMBfVH1mVV
0jiat68MFFfH9r3SF9bfJMnHShktEkuzq5ICX+yYGb0V/r1lRTD5O1kO5HG7aTf/
bsK6JyMYZHe9nUjtKSUEG5Li8Vo33Zq0T+wY8B6moEtXULPtv4cIfEJ2MK434XC/
S1p744gJiO2N9s+jjSEGZOto75dlAT84vvPd/1us8rpgAsoWzuBb5FDSPsOfp6dL
eQK5Og8xkBazULIeL3jYu2mqwIyRJ55UkrGAfzzpPmNfZGWV9hdYkyhkQo5F4/ES
SAYIUHeEyYmSXjHIsrSdBOYkww05uIpAPAL5x+ODsgxcAPX7BAwr35bTWS4gm5Sj
XdiJ6aRhZt5v7ay60PnFC9Qv/FLTsgn2x1/ti7DFDVlccLOoA3oEgtKbw8CDYcyA
QnQfHX5oQEoSmCQDswfqPWVOku7btcgNDEY65F0tgf9FEaVhPs5uPKrolBVYM33S
Dip1wG1orbuKkfGxm6trEiV1AwGpUFsXzFxHFDGOSAQ/loolEko4DGHuQgGSdwF/
cMpShsORZx8rGpz1alU27uAQdQK0sZ1EDccLh48pDvYYwVdz1KqqO63cppSP2B1v
j2nVC4qslJpZARncNWJRTtYfdwtuNItoDXDG+y184kNbM3Rey71NZhA3k/c8rozZ
ta8AjdxoP+BnU8sfVXaHDDInhh/bvfozk6hzqLWBH1hYhWBnBJ5JIkfwe2q9ARtO
twwt6h3t+p0qsruP01UMHn738RyE8IlWhizk+flsz4SuXwdN8qFc/sOhn/lJ/4nx
imtoghcAMQ6kDvXF6M70Gn0SB1lwC+3HCdCP0w0K0Xx3eD3WCNgGchmgxqb4riAN
MN/3lmqpFJ2R+7Wj1C8FjXqmQF+WcVA7hs0AcJkKH/JlfiIcSu7soxI9Ezgjxd8v
4b8BlWvPKdgl/d9sA+z3UdUoOOhtPg0pBqMJoM1w4Ot6H1OM7VfX9Ropjdn7srB6
SU17vvvunFU9Cl6zL/kqQ27HXjyPzCvBAV/0oXALkiD3LXjGIc3fAp72kOCIrUvS
z6hD1ZeZn4kVMc+nxtJ4gOtPyoPLQutfP5SESNuZjYIfrEqol9N0uP4JgRgEi63z
AsposIIsNRxl/VWfiAObPN/Lef8JaiMmVoCxiXBSg9fbbuPTtUt8R+MezYISFr0V
34dParMZzN+KHiK1Ggb395z39hq8NoZypmBbDAhuVfHvSorLRvPA2zKhMG1eCpo5
e/qcEEVfO8OipruaeXNWel9XhPrtopTRYAPM4EkaZbIbVkTXy86PoTo9v0/T6ISH
dG31PfU8hCmcIAfrwpYULVL8X1s5LEVuHH+6WBiXhVVY1hI/+KvTVuEck23qfOls
HGttF4UqOIezX1QxyYrgTCLa110WC0ZObjSNNkRIqlHs7iW4xJwz0oAwUi1M97D7
yE5d2MSGo1SRs0KNs8CtmZCtDMOngu4l2YvJ/Hs00XsZTaKiFothw5vRb68rPxzt
TaBOAcoE3FPmD7cj5vjUvTtfppzC8ziB/3jdXUnOa4zg0CEm8cXEibizBOglc/5D
n++cK+IdIruuKYfHqKB3z/Kd8xLrAyBXhywgZ9a0NrDZa/jawyv+o87Q67mCPe6E
2nlqi57N9W4zqQD1hfJ9QYp4UOv2qwD6WZykI/0k/Zab7bRo/vbfRk/kHt/vL8bb
4mvT5bIrUx2UUS3bxgrNlMCX35aFxObyrZajIw7nXTdb7Qw0EIyaKmyEQ1NHWShS
JQyKG2cwXJVeDMVnVWMgt5BLtEAttUqU/s/hZX+vTPrDCTcZ7PhyYyCsgzLJKZ45
fqWbiO/c9/FZ6tsG8Lhst71lrxv6sL/q8Xu9YEao2IjI6g0hSOH4RZ/bzGo70D/O
0yXbEwAfuSO00Mm9jjzHMo5g0z+NpfeAOfpadHANgYYWjGAU81ycUHUOieawhOM3
rYlA2BGMG0vhkdYgGRjI6lesijt605ra11CJM+7aWvb7dwnmYb49V6UU1DhSxhSi
1tsYMP86Ng56KAQlTXsIytBiJY7Ilo1+ML+IDgsiIlLzVnPrqSzQTx2drJ/GPm8e
iIormzcctAxllu62/EWm3iE0QaO7X8jtOW1FXICqullTElr5FNGnoT72g7EQt2Jc
otDjhoL68gpnUi4vF92u4erV0cnSZ0sqq30YYZQNGVQSaz2jEym40RSiWwtmENUv
+0WBbFwj5UvYK1YiDpDwZqQM7m0c/BL41rwrQkvyHBnHBQ19fT6vrCt7MsX0yMqa
RBenQX5YCkGLVwc9IS1i83RV5IPuVxT6VT68IA1MNIwkaNTbkmWKLe37my6i5Rob
9RSYU4mpGwbRBAbczfODMqjrfJldyIsO8cAtg9nOLLeMZp2nbekPVjAs09/oF8dt
JOAxMJ4NIl5af6v++SGsnmlHm86oQiW/JcGFGuNnymtL5m+uXDLPQK6PtxIO44PY
zM/cjnSTQBUQ+3UFjthmP8oYnkkLVxE3lK44ulJ3dowab/6SU3NjB1+YNRrcykjd
nDeBd5iDL36HIA1Qu2RWQ6U2gZrSRrvGrvcD8mesi3UvxOGVMzYuayCXPk5Zt1Ds
syoGaQ5LBeMaTcYucUgZ/ug/Kf7k96niFDlaoZQn07o3917pPVEbvbFswCIZfiik
El7TNTsOUAeD0RrKe6Qy4vn87Y9r+Z4fxMCD9tgZ56JhS3eR/W3irz74SdXo3Owb
+w1+2c+HudRHqJI9tumwqN3wUfI2dxYFDP3yh8TIHC7iAiwtMS7/8jHF8ol87N5n
ZfWrHEe7UOgJ/2TXYHFgdDX1PqOuY0pX/01h+oDLzAYDJrm44zY3e4dveHdXFFfv
25C5B13Oaa5jXMdChtlMJRAJWv2MGg8uv3HqFdilNP/BMYDJ/sQ+2Vbk64sQBbsT
lWHJArnHAcS3wnUaP2h7+MUZKw60VneQUAHK7CvG6zfsg5xUzzKcih4NrrqxC41A
134FQ0PgewAOmNgAvsjIuaDpRapV8XvbgAXmgRsGFveqq/Ovc/iqw6JppXCG8xw4
A9E14NuIMshlQqS0+bsj4n6r2XdCt2sXjEtumXcDVt+ARy4sEkyW4BLyg0p1FTvX
Qgu41VT0Z/lBlrRg0lr5orTlCYL/a0nWIA1OxbxL8f4jqOs78MEVJ6gorsyMgWdL
jtAvo05pQEJ44BrzbmwFFfID1SYAY/n3DdHu1ntntLQYGJwCkaSrSHUUge95RHRD
aKyTiDrhMURBwK/Or0MftFnhM/F5BmxNrnFpysIYz6cmfAABGDeYRB83MBQK4fmA
V7FnyuZ5ZVcxiurdVij8Qv+tzSY/2iDc79bfarry0xAKYkjhvzC9F9apVJ3ixTJS
JsnI2GwnaRIikVFmf3EDD+o3J+/6eD/U9aVRYdaydalgi8f7Kj6QK/WT0RdEy6Nz
f92jmCQTtOL8QnQjL7n4EC+eHfSdV3I1YxObUZZ0UErwu0F2YXT3YugSyADyaEgx
xYVPMVehVKXjVXabq2IC8Tc1sgOQa4rJI3zHtUE2c5Way8lFbER1UgSkjud4BJms
brYaqJnpP/3ySqfg3vCvMTIlQPOeov2fAtQPLe1+B2Ark9+TyX9wWgIOhw55Sqs2
JpqUCivLriLvGpJY7+Xueb1hZB8JeeriLVDaUkQBRTA1A6R+YVAFPdB+oFqFOlZH
CRtSfNanBg2JJloW8KGp0CGHcaFbE0s/msDS3WXvzxHN3ovivbyQi0cdIiNE7pOG
XN29gfoDxpme6FLPDHqGb4Xyj1k09JXx8tqh2QRoKN4x/Pd3BrMxQAeZ8aOfPkF5
CDcA2GYA290IczwlCBdLq2gR8+RvAD3d149tLQ8iKR/aY1h+8d3Hyisht9GptonP
RTDqQ7u8tK6heizc4ICV7pRk+ofGSbD8pMQq/PscHMp3EcwT4Y/GbN8EYfcAb5m5
vaE07WI5sMGEUErxE0atiKO+u3fNL2IJxSGOvuQM6FZxQF6fVki+snEiaS581n32
XwxQkmg4Yn/yNni0jO7RHva9DcNmDJTdsweFXCwE5BFql36uthjW/uoPanBceARm
1hlpFMHkKGC2WDpniPxjt9DLFfBFdbhT1fSbHGgOlp/XedO3DVVZOjlBmxWvoGFv
ITcpCsHTn86940/mSI4E9EX5eWO7uKrEkD4rQII9tJksME9ILFLQ8qn9S1XytAWi
7CS5zHbQYdU2Ax5fIVCtO7ufHmKShc87wbTM3vLgPZvdbOjSci61guDNSHmkQnMk
hB3POJh6LeDSWctJzZVB6iRhsaCWP6K2fsL6F3IS6K/jqZNT1wWuVh7eYISgKWMA
C3bvgkqdaOe7U+nqvwTBt+VmwTpTtHrCLHINcgTLu8cV6An3bgdl06J6dAwUTZ0j
A8hgoCCbi2qOODE9UIXZWF4Lp9xQiV4LN7NrR/YFsn8nQzdKNXLOM/pZGv+suZ4v
vouGRwrauilYpDq1AqCBXUv6F0ZoknyPvTCTI1VRgZuUxQqlxvH+1h4jAo4C5uxy
5iFxMs3/ODbGco+O6ROFtrNreVnYVh72hffiPecAPqeUdIO3otGarQHwTZKbwVyk
3pCPEdn/qSzHcWM0UzqzJbw/2LkxODbv6A8qbETwW9tfogG2lXRGjse5nAWx0Mvo
Nux9V+5lBmUOo1M8AT7XtzmWwucgUI+hhzDYBC6SvE7NYMaQu/EEL3k63spHD6O6
ZG6E1n7fUKqBPphuLq5OJ1kbgu7RM79AV/Y6tb84rykhK6uzsb1HLUjFmMYx4gWO
aXqeZAAnAN6CRrmtpwZKGXzoA7xoM6vsvTkVl33PtOIJHXx+J9Jm4EUIY+C1T2x9
L9C3ip8UMNiOtjS6+Fwp2RBfMXi3kCkEVhmGtcV6wwXj9050HhnBGqQ/Acuip40X
fb6cKbfmFaUJva66h5bv38VNJWpipP7VAC3ywx0PDk9kRnhk26j8qVVdWTixlvsu
g4YaT9Kj7esh+JyxsDfdkHdrerR8JwHOdAZnQvnGp5SHZPGXyQJ5BUKsmXF5+/xl
cH269fTxTOIAbn/2YInKKHwa9iaWhH+Vw5TTUmNTcthDSbO5MDamqyJ1K2oig8x1
QbloaLf/LXC2r/2QXDUi1CE/O61N+VCoOOMa6Mda2Jj3Qly6ZVzGl7IN8wfrYray
63i2ncW5/UuyFnUXUIIQGGE4NY9jNbVhefFio8xEWFCxjaBWTutA3gti4UxHdL64
OIjqELgTRNObZOoUmY8VolY9VkLX2/RwUcK1k/oHfnDkgCvIF0g46kX4gFaEZfqI
2GwzJK1XXSht2obc81Lv/bo08WWpvrwFamdWKr/91uS3wbRaIe9XmFC5V+MHcBjz
WRd2QhC/GTmZUTtl+JVehZqrOlCQKRhj8ENDBP80aBBr1R+rwMwcOVUKNpLE/6IC
mVuuPLRL7L9VtfLINL02N+3qzF+VF7g1jZv63fu8VSZPbpombgpyow5STsxWVRDO
30L0o6n+8ymo1PBc/nNt/dalh83otzwlAAgFj1uQ9tqFrvd4JpXZdSdl/jMm78Vk
mFLYk3srnB8ovg+RkPJdsmbDouIye0FxeQlK7UfOF15X6np8voRyoStnklgXPk8m
osNO+ZxodCCJW97j+u15cVL68j2T22TAMzlsxJlfp23r0HfWfLG/xAaWO+Ogph/T
RsfAR9HP5dZ5JjQOE5rJsjjvToRDQxltTERnSINOIuFSyGm8VKgLlw40ThsbQyUV
J9EaO2o0Fj7lzfkaV1RdBdLouTca1uG1vG+gMgHj6WJQnkOgMio9WUhORzkr11M/
E92XwPsyUGUGM219paHtdIORX6MFNu/jQ0jBh80Z0hE6mUgF3xsg8xOHxXBc/X8D
imyFgcePElrQiG3D+15E7D1cIS+6M9Kwnum9YbLcrq6ngXSqZw35RnNJ7pplJCwg
LsInaxKwkNACBSx151/KUiclkvtnZdeX1s4hDRxuhWGTIGaRq0caNk/H7Rqt/buS
cGf5sMgF9Q8kNTinpwJjXxULG7VAKOHi1g85jZnXHDjfP3WO7aN5m5CJE/qlF1/2
9dQTo7BX8LszbUbdImehf6virlNrHrTE9HyJ+u50Z3BvY5K8uBlgDJ6B+VxrGSGY
VV5nr4Y5fQaWt0hzpmmLI2ig/mJATBeX7tLhoAwlV6e3Lru3YwIiHV2jONOthe7D
aBKtml+FZgw3+W/m7UzEgDHKf4xF8xYhH5AVrkp0DCKTkgPiK6z4dxbbbYIKb6PE
9x1JObkjs/l86DPJx1omqUc+VVhOs8RcrgA26EvszYFEjK6A2z8J/xwgZNHGWy8r
QcMoSpgGbumg50vHw6hTfFe2yDh0hxarSCLZ2l770eLlBOE4RptHv2SRmLOjWJGf
wbaUmxRHLp0mF+PWqB2jLTQ8zIq1l4c+uT1vUCesJohd3DSLU03nfSyaFUM++m2u
DAtZKcwQMoHPEm/w78Pkvm8tLA3lFMG5nz339YUZ8p85NR1YhaTYdD/wpsjdX5bk
mbqxNSTCkppHm3XIcZq0zUJxUOp4hUoviqJwvA2Wy7PhTF0KX+NlCEk+m7F4X8lk
BXaXQWGTTIh4ECxIxg6AGerGM1CA6Te2nqDG6j3aWtk=
`pragma protect end_protected
