`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cQYQHKOOFjr/q1b/Omvz6HQ+PjbPtNRPCVfadvj7bwoV1H0azNEZa/6YY7Wxjy7c
oIy87EP3OlVLCze9OV9fJ2Hmtr9LGyrm2bo2T5gHxkpzNDrisIyrBySn/qxzg5/w
bsPD28z5vEOLYBAZ3de07rCp+qn43/co7CxQZfVvrtg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2288)
KK4pGhuVbrlUky0yGZMasti0VzEgdOaJQwNU+oQDT56MGkwgZh14XuIPkarGs6/k
4/Da5WUuFiNUrRsnnIf+MbkK/rvGX0GbL03vhOlVUDtLj6qUR2UuJ4ky9UMyq4Lb
mDuElU4q9hHHRseoIF6hKPPEf8mLflYrdYuBfC3/46B0lFYKCQ6cKcTubHEBF4lI
RDhSAHBb/PfkDqeXvBg/cEg6AJ83h90useTbTkSVROHPlgii3KHUKNWmPwDQEJZ9
HhsMyFfBDlRPIIqjHuo6M3gS88vbxE/O1vsc30WHvSUovXWTmqtUV1urfX4g3DyY
b12mfN/3+jnO/ufysMnE6+az9/nvX4BrrX8/Y3p0ETWCGA+ZRN7KMgDbOhdul5D/
1gjUXvwc0uQrotHph9Ly+Aw+HwVAMdiSbjc98nGy7soOL4ZuedwY5brk2Q4KJL9V
xorqGsF4lBg784uAn4tb+xQP4zSy3seRBqdCrZzRf8+Bv/5XJpDHlY2X4Z7lwo2j
GS6xKTEWhXywciNu1BSC4we5KDgvzT5PKahLEEWSYncZgOL5jcqOrzQaLJw4qsQV
ilmsE0fxdADQp+cmtXM4dLjNCBr7qWYGoZd5J7b4aRadt2rU211bPHWoIyz9KSTO
gvaWzqBg6r6aqHsehy79/4bOpXHFWVreDhIRHH02MgiydkdYktN/JWDHpzT7UMfx
KDWc84lCPUiRA46+NeDWPZ+7MwDnUJVEESFOzc2X1PtzSiPN5N1d2/y2aRMFRFNK
4Wv71SQQ9ZIA5wH4RTibxL0qJpp5RT0cnwFROcV5+tgr0bDCRswI0qBf/p7wZcS4
Ctz1k1IosdQ7krTrO60MD6+uAnqytaYUMO6sSDAboK4fIinm20Di/p9eC56KWzow
Q/U1ve59izzCJIb8SFhPeOk/pduZjuJvmO0tD0xNVXDbtt1ZGYTK8tHZXeG6UGlf
4IKDXRvRbxgCMeSq6Ka4VMX3cpsQmzcq3Ss9wg/yDi+P4WptL/eWbaP5bjkL0Zgu
ZkqgZ4rciPZv0FzzllrMDjcFPrK2o79Hq6Hlc+iqcubB7B4skxeDZULv53UqoRSP
QNUULQ2W28jjBNpcEuFSIuBo3abiOdDJoYGK1xswa/LXRrtmYJxupoWxQUTpKHQq
opzKTmacgA+kuaSHi5AHncvMA0IUEZx4NcbwSNjxHrdvjoyRGWjucDeGqcTAWFSj
0Fkq6yqDY9fnFB4VAk6japlYBrRS3bkYMV1oLkTtps/e7hF8OfC2LpejePsEzf9+
K9HYQy2S4KZGTuDm8CowG5X2ojqpK5nA0Ga9tO73rYwSAzt3SDRyX2FnoPVGcP7I
+bvxwe4HLm9WfllEb/Y6BiMvY6GVRNv33SkgHvbQNDfel6dgHg4l8K97FkQmB6Qc
gt5wIh19/X5WVjy92OTdWsQXiVwpD5D6i91MjVLSjMwwfufp/VqiLTdt/9Is/num
6wzn/S1yQbj28Ipn4ZBe8kCufjjU86oJpqcHItGlfxP/fBsdN1u2+bwWyLXvNZQA
O3EHxEPajrFVAurVTozOebs6GSRQ9zSt3yFVdR4CLTcgvyevt2aB+1kSe3l8djFz
GpFb3i10S5xuA8a61xF7GTq2qXf9/oiG89ukjawd1qfAO2n8n5+tq9a++X64+pra
fqqQtefYzWUHuVbC6M6HnGNsX2R6XRGb+SiVxk1B39LURtpykynU43Kgtl9ADTUi
LIgbau4BJFQrU9n1DBsHAfBm2UzUxeQRGUoD+ZDbTXUd54yVk8NqtBv1uzgsjkve
Mf0XlfwG4+/EB1lplmNaNA5uXTbzfmnLfn6D94OC6D6kZaPbOZPwWWmp4Xiemhao
ncdoIV7lV/E7UdHbnVBQbYR3C+ZS75Y3Zqf3+gifkc+Z4aEGVrL94OZe4iJM4h6j
OXd2SzTDKQuMakggreZj49FjHqUAPclA5Hz1irg6bSy0BJI2HfNeRCRG4CtPhIwI
61v5i1pa3/1TWX0t/0YD020NZONJf7vINFh7ox14jl9tf/ZRO1sRVjDvoD9L1ooI
LgEdCYj51Neve8Ga+EFdoQGM/riOalGikBN2likYhUFi+0ncYtgoG03iLRdg/WWm
ujC4lJFQl9ga55hbKwbLADHpAcumxvAkcXRKbFZC0Feh8e39q6kFBQpTix3GpVXE
aEFrXPoghKSyxtCz340KfjlHeRyz5/59oboasqtE4pyvidXcImsLR6xePwp1XGb4
ucOmONpOIUeJO7nNO8fnkDaH7mG9OFWAno4OejvhHqIk9nhl0wCCHBeJMfWnXVGb
9ZG0Ot7tLMWnhy6ogX+UzZTfV6DE5UpZt8yZaG7KjLwAijSAEbwZ0Pa9OIgm4OQ6
CCXEfGs3w39gUtOdVN+AgRXj3ugH1dkvBEmjLXp6iOOAUxoJMdBgqrnDTmf1rZBA
3R728bF+ZwsmeHP6VuynsHQihNmSrpVkyuEKmh6Fl9YoLSRrVYunUoFfFgYeotIO
K2xCk2SUiEyeXB8eu/5ruIRkWfGo/3jPEBwte3joNh3vf2eF6JXMtPHaOVKBRqgC
P4CR9T9zk73NMlZRJePOMKrgMpIkxrL6oy49JZ0DWX3ookrEIpPtHM6qxBw/7t5I
0ThV22QjZ0a/lRHuiP9cQe3URFx0hsA50H5yGQg1Kh3LOHJ29VQN+bR3r804qytn
Gi6vy6P+Jc4bA6VbaPqB2iIChcHyV8AyEen2oToG40x8bjj6Sl86vFzaSdSQJh1D
cOEKnPxkxBN7ujXmkp9+dJSmWZesGIhkHEanuzwTIA1Nnim7gWVYkmB0Blr4WV5j
IUYpq61xdhlB0/o4Dpf6VGdNzLG6b6klThWOCoYru3jMG/T6+3ftb7Guxy/0eX8h
ecjAHPwaOyLEyQFEMoq7d1DOgGkv1BTdvfcKdBz1mAF+z5hs193y/XdkVSIXntZN
RC0aNbu9LRjBEzW4CUF4b0sL0Ryo4h+2aKlAqXIYbyrvibbEp4XB3gGfMinovsSs
wnvdTc6mFlGHgefAqNflBJtMjHchXmUDZD4ktQLj8sg=
`pragma protect end_protected
