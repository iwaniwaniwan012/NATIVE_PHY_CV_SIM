`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UrDOP4/L6iVQti7hoJoQz+7kJ+B/48Nu4GGsNdZIudRoMj3kHuHFIl+vkFP676Fu
X7womWsvV+yE5Yg3ie6INzRF11S4QqY5VAolIAJhOuzUdZmsQHz28PYM5QA+3+6P
EMun0ZibZ4mOarhRiU5t9wkCy3BypDR2o9lvz/DjrGo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1728)
memCgFSB1owRqMDQYYvkyDxwsOJhhi/qu8exBh7aT8SqlAk18hafvFqzce1VLwh2
8ObpzfflM5NpGOZHau4Gv1v4p6hm6rfnuGigXluh7MSB0S1BuR9iD/RmcEdusjeq
tWe9tetiNISZjqRwFH7/a2jKRYd43jicWr0WnvxG4cCwRi+gs0GKwlebx+0sW0uq
Kfiwxdm0d1FG5eY5cpOsAXylQ3ZJXVK/LOa8XeREs/QZiXYnlI7dzltK1n8nLXlC
KIGrnDFeoZ5l2rZn/S6v5Oo98Z3jUt2g1tOQr9mykqk4X4wg1O2rgTXS0jGk0RCv
JS/AY/TnDbDETd/kopEyrs0rrARwuwqcaVrMy7Cqmi7Je6oOdozT8H90UhL4eVNR
jjCzijDOac188ot9ezjnN3Mlf8L13T8iDoSx6JwHS4AkFaTP2ffP7Qc2dKpK6Udy
VqP8y6+1OyGWBCzHhIqgh4HZ25RVDLGlz4I5WwHMQvqPw4z+NpNEUoOFCKk9i/EG
YdIPzV6IRVT+16xI7KoNzHhFykbl63+pfsPv9JGiApa+M9sZ8tewRJOZwfVr5DQy
bbK8eb6yKGzgKJypJXmtzmmC5VzvEzZTmssaa6zdzaa6z3c2nNsIJ6rjcu7ucUni
Mm1b0EWmcmXaY0n5AvDJI/mbODsH03zONa1yguw+pglLUWoC528+IzYWCHa9ImRS
knd9dtzxWr9+lBkZKqLHyLVOzeWQS36XmX2KF7j6dATPTnL4w4mbJD5coTa9uWXi
oLKIN1EsnaRlxtLgD3naqC46Yn/2PfzDebi0kdtGza9GcycVR+IxT20xO2J7FFn2
mDsTG8GknVHd0bQp0AdyLV0tHgX8Hhagl3iT61S725Yez5YF+zECQMMzW8E6LhZo
QVoz+Vuy43foXhhiegTaJDaV8LUZvQ1RsNQ6ZWffj4RBGhE7DfvQJdyL42Ui+7tV
Zyb7ClUclG0xNaTsBEQ+PRy5UXCdEIdDli/l4C3/dg9caSlrfKmbbj7txUpYMpLr
IN4WB85K2Zet2dnp2f4i30wvv7K1RhVVw7TwFK1HMl1p1B5wdG1L5Aoc+Yvz8MKw
ffvNaeHKWloJrTrq/lTHVJXF++8H1X+APp0ab0mt0Q+eJaBPfyCenZgkGFJYYxup
NBcme8wkeIWK426VTaseSSJKmNLBE2i3jB4rnvxMT1V4l+8GVBtppK8FSiEb1s81
Qb2E6i1OOt7EChR5RT97EnEHhtk1ICyiuYnrzOv5myJdHobNA34mCzwHCJE/z+I8
0TY9O08pUC/92Imdk+1mhPlopqZ6GyJtskrj2wuS9YMu5OFFYKX5qiwKijFdS3k0
3y+i2i7uhoiQu0y2WOYnt9InNTnsv/Eb9L6IU83mF8T+6n1gGLNaAts2/2DxfBTz
8p6w9VheDD1s8qRIMODxRJlnTHj3U3aR9p0RBFJqLlYUjtAKL/VL25K9VrcgKzDn
fNx4Q49CjSrZI1CKoCHSVa5ignUD93hsq7LBEEp43GrPXcGKn6SO2oIbU1enLygt
vhnNaGuZnp6Icff7UboP3Ho8lI5rWBTeUqHUfYtzi/ILSFU0TjuB1JB3FYveqT9i
cRFpvDS4lOO1/kLsiV9M2gR4PqARrN9E6pqGIX0ZckxtBqgmRT38wbQEddTfqKdo
bZkZeEN0NGPyr8KE9vqyFrSWjUjf4mCvUYZAgGIVf/krj/WGSEfxXJ/lB8iV2RHm
PLkOsTfJ+8p1/ckXEx2lsa+DENEOVZxVB4E4UubZKIOy8LuH3VzqRYBpf1CBLLjs
f9KxnHgCWZNL+hfMeHb5c+cTvRcUZefryidpwt/fj/l3jnvH59tpgp0ugMmu3Qv8
aU2Lg5UjWuoYtmlLu9NZNonJ30b6Hdftr8g5x/VhRSqLmSCgAq1lONYkKA/M2egi
uiKeSzIv4LaKiOHfk8CDRCpVYNu+RyRi9K5KMtnqQ9FxqeIfzcX7NIUqKIr/2NFg
6aEHi6ZgcIVbUHTud+VulhuBAcYtP4rKaWgOsP4plmfHkqcPpfIBEwlrppprUS59
jW92rRK6ID5F2Aj/AwCGvbB0kPT2ISjE8L+BsB2bshiYHnQv7z6JW1EU8JrPuz0e
iNu0WbKziUX3XTqwJw5Y6H0sS61DzI1A+rCQ2kFBUiMILMiLhTOK/IiScPWApbJ3
lGxz2z2bSPDJ0lPs85aUdSEg3Aw9VlwYsssoTNZo/61F2W5uBkcN6JySKjj4JTBl
4s5icETq8kJ6g9VRLyOQ8fAYi2TGYNYkyzQv+N46Zw7U/DsI4XtfdORQnkNLRe3z
`pragma protect end_protected
