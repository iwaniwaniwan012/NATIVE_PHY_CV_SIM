`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZUDcJ+8AY9+vA8d3qh+IjKwLodpyr4nVVbOcHjBs9so8YPkUS1cuwkKCwsEequws
nwZ+tzvxgGQ8YZGfHTmVstPpqQ3V4BWzfsrVq06RcbMTARx1zoYqOHeY7LBXVL4n
JW7eTBFpTo6Tip0omHQwVJpjgwSTRsRjpHKCFjNB/ic=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16704)
5/JS3Y2AiKjo1ohvts5p/VucJD6N+w6KPv4PokLE8DiUWHc2paZiWeGhzyn2dJgh
dAv9MZ4gaBKDPqvFFiX7Nwi6dqPTKF1BJrc3+EarpnmMj+N0Th07j2Kzy9WA+ZKy
gMD6KCqhbCklKO4EUhwgONQzTOcMNJ+woUYJSHTGoj0T1G9d7FTKF1l/Bfh1V8d/
5uFdwEUP7+IGU7ryJBLPVXFEiEE6tM6LS1AxvEN6LeQiOknPuFkw3BKQTxzAi/Ix
/cjLNxfV67TjabGMKThDzbxsUXpVjHzs427a0zxMrS9yJ9TpZ/CS+XZ4E4HTpWoQ
McMoE7Ifo+ma/auSgJBMwggNGmUoUuTOkuSIapb4fLpY6Na56sKehHwvIZ+rsuYx
mk7El6OJDFwRZKNHyU4ui5RVwJyKmsJXj5XzMP60q6ILe4jC60X+fyJ8RVrR0che
dr0RqMx3jeAsj9F7i+eFctBVruEaRKRl0FD1xggtYXAuttx5zKIlgI2M1ZUdEBkA
0RhiNVGWKI3c5jkMphu0R7wVnJ5whCeDQJ2GakL3mP5miasElsCYFGtLsk9I9jg2
t1JN9RCiE41fIpTp4maUnnoNjR57cFi0FGpd6tgzoT4WejignZIOJoo3ySWDJE4c
gWLaw9epa77FZ8n9Nf2Yxxq5xGGxS0nMPK/xDwGMSES2QwLlSvOlXI6yRTxe3Vxb
bwIn91RxUlSwRW4xMY5YI6KvMucT4U+U3nvTparXId1AF7g9lsIT6GHVCONnMWGl
Co5g54dwaa2Ey8V3kf1zHhiW75rGy/mHZZu9MI1eL6ZxZu0j4EUukShv+X8VWywm
692JOeWS/011s+lHjmkM19g8gAmNqUxzHTHTjHwiYy5LrgbBpr1mDNm05E93mOVi
QpLRAjWPT3+zhjEvQDzd29g8yzXa+ETabl6X5KyKr1K28ChknR0huOzRxdsok9z4
9X9tJvWT+Q6n8M7d0VKSEnyjqx5FcmYQyBmyYQ35TdPemeRyq8ugf8STs8nmG846
8FtIAFRVR7/SR/I0IGEUsDGVNvKpxZP5OqR31dW264zkNqayEhIG3bOeSHagHmfb
mZFJanuCJ6wqZBDWgxBORavHmm8DzOmkPeAq7X64X6nl0GDSIdpN5+N3DY29pCXV
yHWL3jKV+YW2/p7jIIiph9zqQRYtGJ4zDeN9+5ztUrEdVfvyXiFaJvRUxm/jay16
kfPooBg+kSfKN7GKp3pYDZHaWBqLCmJYsk7LqTQrzhGAZ1mmQCe8uSpRTfoBH5Fs
LXx3MbYVIo/l3+VwtYaPv6v/Nb09XJsczdC6uBa4KEgMyqyFROtosODMfivPH34n
gjt7Sj/Oinuvy8hVF5RsONPI97YgHRwDAoKwmxdrTxpmIbsJEQoRio2KSjljQr9e
2Yi2wupdp3tT3udmCXY7LxgbuxqjEsoYe3pCrNuavvOm5HOZezcE0AAZTI3Scf1d
hSPww9wMW02QUZgSd86dmTZOjGvD5+VfmqmPqZwOU+3hHRcXLVgmLDa0mExvc+LR
kM1a7AWPf1h/BvI8QMp5Hk2DDdq7ni0WURtbxREtS2V28usAhhJPHcWf+LAobo04
/zRo8Kc8EWdxca/RMItmZhhfx76sAyobzospNBZtvBfR11WKq9Ewc3Qfb5sD6Bm6
vlPEeLmMnvUsIMgby9zuX289Kthb82qG39Ks5kMjgMJAzmZdfpZ/z9PwanTurhu3
HKv/RdX+gDxkhSQ58k1Xm3tWFv8ndxOqu7VhgitptvGDbtTJGYx3ak6xsKKJ9NQG
vZ4nChHQBoSNTI8Y4GzSsCE9lms0W3L4m5EZq8FbriUqS8l8NhhXD44FMcXrtAWm
e9iKgHPeVhpq4MzAbxq+IAvz37+1g+O0NgDN5qKw9D03KuufX37FnKAZl6wjmDOH
yGSlQaivZxqC/t/FepFI+yBtt9DMKyOpyWpPLxItrVh9B7um+Fn0sezFQBTAs2XC
3qSqEr6aXVMsoY+8DbLqhXrkfmb+owDULMuhqJHY6VD7/rQuLKj94cppkNp0564c
ddJV6BSNitKXE+N0o7h7XCAmv3jG+oy9Qidod2g3RaOdvEALTmsdtAfJQovmTbpH
AqRdnczxng6rfR5rjaTMoCajsgYGkYO5s0oAwYZiDznXS9VjucQJiQBFXPuMt9Wl
wvwxMYvIieifMqKQOMThKEfcvryamjx4OJAjtuLl1+up8RNakJTqjqLec43lKiTD
lkRNnFXGrh5b8uCNluRkAm+VlYRc1Q+OmeMiBOR3gUWzar+QNlM8HnuxfCG7iE45
u6RJ+myteA+pxAm97etwOn/MYTjS1GyRi26uZc2Q8m3oadS2fYS3/C+9/Ft2eYRf
fMj3EDwgEvJuV/F5zG9Ec2WBn5dZP4Tj1zImaeBYdnbalsUixs7qalTQFqlH6+wY
bAnpnC3a/d+HMCOKMaeXQrmyBSNp0mciO1NvoXwDsU2vlullH7fcSBPIchmEboYt
Y+XkLp95aOOlcZoY9RuY6xEOE6D/IDH0Aso9sOIuq/N9DAJgTQR8QcVU9r6dBXba
apEiuElPpvQEWJg3nvaG9FvpVZpmlvVAUUoA4/Gup5D6lBw0GAaVWiobS5MDzb9/
hJN/jwpngoDcvSQx4Bus/Ijl+8YPfYxztbw31IyQja5v5YTAIZ8nveZmOofl0bv5
x99oNJTbDnev6y3t5zFIon0rmJhozLCjtyTAaNt1gugsFz9IA5/US4qN0y+vtsj9
YUVrHN12oSYO/5F5Jaaos2R62wHoP3SWYcMbrQsxwfSL09Nk+OJlT1ka7g8bPGFG
168JONPuAbqTDcVSySk2a902qfS3sBFIF1rY89CBK4tYkjskl0zYoqtCkQsgfVzH
PUwnvXc9WvZffrzKBQJsNM552Y3fm0wcU79Y4haxeVp0iJSxCd9Xjcn6csZ5Uzm6
5u+4B4zSBOzNem56YupxKrvCG6PuQrX+pdfJNljcF5VxABAcKEfnj4Q42M+HkQlf
/OuYXlnAnoZ7pzadNI4ocAMJ3flNqr6EHmkHAm1nbE8Z86LqK3UqAQTZLcBIUkDO
hTzy68aSSQ65gdDVd5MWo1MWrRTqXmxTAMoogK2mf5j/lSmq5eFRhbpaVRVHpJD6
TZIbYf8ra+z/tj4w1/wcunt57KPvGY64c84rGXN+PsWTW+GpAiwHeaRQNhs/8asw
XVEHkymQjoKPuNPT00IATIyLnWp26ftzoQp9WUgeRbxdbauhJKEuBWrW6SRrCK0P
2c7dt1DlggAkG+ct85mQNLH5M4x/Uq9muOPpWiSjmmThR23Ck2ZcYa6HzCBVKfBD
njDIZNbFM5DWLT2xo4lKgP+JrDeDfzCuWtW6Z+PKpV8MIznxir1KLLNIykLf+D3g
q24eaR6dwypoeokPh7EH5qnyLEHo+3hPm6Y+vBDdU9x6CDVJksk6ZxiohSTnx2m3
vw0NZJmKGg8M5EII6ihe1RgTjcr7s0eesk0RwQAbT7ZqLfverWpm6DvGDR8i6dUR
NdHduGCUmGbPcUHhtpv+OsCBp7W6JhHysHg7HI7qsmEK74RxLoNfHx8TX8cF+Ubl
DYha/lkaPpzCbD1r7XFwm3Z+XE0xOkd1/4sb3Hu+RX0c2WfNqMFlfDVglT5dT5wf
J++1qyZr39OdDSV+TgSIWpLtoTlhek/RZDLeYMdq3EfBd94zcGmG76IpOLqWQ4ae
emJHAdiDet+vTYAECEq/WQ7FidUakCupdbZyuIRQRHoOdB8s/tkuEr0j0ylU5e3H
Xrre/7qGnhky2Igo06crFkdVXIlvL9Qe5v9zaBSDBfWxvRjnnk79Bk6WnNtEoDCu
djs25ij0Ypyu0k2D3IicoifyJaqz/4RoORyiw96TvWL5lIgusQH6Wyo51SZE4U1B
IY72nuM2DWh8cYAXuGdp54YTbFVvUpv9bfDseGnUSJlamnoZRYyW3MHLAjoZ4lKj
iquJ6A+hG+YDPl7GJMzYce/qOEkrmp3DQyeCXHj5GRhiZQaf7+03c0GSiwWraYWg
vgG58h1S1mv/mFbvWiNlcYy7sDoprm/diRukseKdBDDmv4P+tRY0mX4URHo6VID2
iW75BycFs3jy+PX8YltyEQihNeccQaEE5V8djyjxj4ezm9c5GpsoDX8ZtbLER38o
G/FhtSQEpfzZwMuroroBKX0aE/QHZKH0B9BVmhxrLAer4bMh41FS4HjERflEyKh2
i1rjNz4VfvNEqhFEEmcJQZ7sc1zDcLltdscPdvzkD4Z9upcc1FWtOp+u3iUFetRY
cNw0TtrvNV+t1Nna92AApkbYBqusJ4b30oh2LTw9rsm42wzGbZM4sdjb4H/77RC2
QcqLl97Y+9ajSsz5UuxavHX2ikYq7DhfTZzVwoEr46tBXnytI3V9X6BjQ+iGQg+a
FLZkdoQEneJO2oeXSYxL3mqfwhhUfSPY1L+kdVdGgpQ9t92OqO8WFO1m995CgsLZ
Juhg4hhDMtgHZ0j4FwVv33XLs3+MDxovE2NF6wt3JNihDvqrOXGBlS8HCiQfahw0
p9LT/c2G7slGRYs1Rmns/vpocdz1tLfFjsNM+HWno12E9owEusB5ZoK1bz9ndRkb
DFSVouqFNLL2yRcI/cryhX16XVweekzxPpVIz1JD926yNgJxb77eWnsYuqNCmxqK
0uwtsN7etZHKcs6q1E92X9ObfZQIF8U9onGJHf3h9y3rw1fSmpAm12S0+6BaYhVx
0WsH3pyr+8mcjRso0JcinRT0oUHbRWN1cO4s13bCL5tDMBNtVRNJc90SFrrNCcXu
zEkwZO3dLsZ+/JENZZkTQNs8dfebEK8vaI7uHQS7Epp/U/nljscvq2qJ5yE0cYJK
c/GP712w+E7SZ33YsWX0RaOVsPhzsJM3A37hN8dp+wG6Stz51gVZCZHKt5KteLCR
0LkD2n60Uf20H18Kma8eHZyyQ7J7tzLofOeBi/zU1sEOk2nO5X7LAGVtKEEYfC/P
XkeyfpwJ+o6fhPl4Vk2Rja7hyDPiG1Tim3+YJtjwF2RxD9GfEuaVrKwS+Y/DP1/r
omFZivLRQglsbrVFZSu4A35w+RkaZVPL0Y3+LgbBc0DK91GoQ1ufP63GndhAABsb
Sj2LHX14sDSldou2YJ2X3AwHfqp7z7UoLf4Fa0FjH9MQrRX9AdBMBAuZtz+B4wI+
ANKxq3ioAd4NK34JiVvSTNKX7RmQAPbLsewv/v38vuEX3BY1G2Vse+34a7YfjhLs
7r7kS5JoESI5HM9677ypBqbdbdAj2v1KxR6TKpVVwB0wrMiYfv1CLALRn8JFclzf
QC4E5bg0FXlx3U/hf9E3A5+2U2jXAPqL0dQ6rmb07t+MwYgdxPGFY3YrB0Ii2/Yv
5MCKvNV1VJ+qDmo5vXp+rVRjDMDPzx3cGYnVeO1bk+Da3aFJIwtX1KrD1PYcryzj
Ep1ZwVcQGOVFXvLMtRzKT9IfRsUW+Ubrq1eHyFnnmcHAqYsOCWyulmxkKUF0uuaU
GAgXF7pGtQCLMEhPV8CIFcsP0PGkONDq9rwi+Qp7iU5PWwPCwCm1EurbcF3sor7A
zPSR00+FUaWJTDD/UhqKPAGjTsTrt69vTG2TcpzCl7mt0VMZwYwmvRr/3C7S60yQ
eTlqU9vJyMkAzYZ5yeUm4jxJfWdX+a25W8aihx1QaiGaYIg0up4ZiHVZ0GYFHoie
7fSEh6rZcb68EIJKKLsQXs5VBO8UFHEmnfgE4ic/B2CFN8i+i3eDDDesqyAMvdN1
l5NgGS00kTrcW8yOD60RWB9S6Zxfphh53+f07vUaL8AhDPue8HIV90zc/hr87Ytc
ekvz214bCn6jbQx/cL0FpZPNihxQ8rAcKgeRJ9heWv6B4K9SW1ve60xII85xiL5N
wqjuTyUI842rEVTOjUxkY3cdCkH1oQ6xgCR+OWXtWOe4llCJM6uPQfuyIHJKmIuI
z8lvrAyvGcQ5lHfAZWODwgpwtV8clrWxyYVznGDGGGfxMfWTdJr1XpLaN0v8STA1
C738ob5X7/wbpq5JUHYrS+H6YbTHIHu3d1cqhmuTdCxRU+whOR3XKMFoA6P7eXSf
pDLow+J92vy+X5CVbaEFh/kLdLsHrq0joqAWLSUujawWg7O0L17YDn4T/azrn4iU
YQATfnKxGr3kNepMjRKWx1wUzI68ez3RF0MGEyJ/bRCEQ0VnOQyqy0ei6QlllnHZ
WaXy+JJ4Wz9/I9v8yh2NMW5oHXsO9l+g1DIlJv4t41f6smrYhlEy/ce2L7sCNprB
DDp07PG5gHW10vnCDt7TLkAXVKLEgT4aOqeTTaEIErfCkJKTIAK4v2TiGwZiO0IF
Vogv+04rADa+7nBMkqLtEBTftoFYxHpNRiNc7LCRiVOXGoSV3XxKBvgssz9bQs5f
c5qrZUKZ4Oth4u0NlwyoJrn7LQGKShp+phD5AoIg44m2lmnCvCb7NI4d1sBqckYp
oQ+cesGQTw8OYMxWSScHwzOSEpkYLcTKEEfwlnooh4Rb2DFbvxvS7B4/8ZYfREuk
WBKSV+zX5bUzmSgIT+aPf5HOU6VidIWFkx2pxCWtcNTC87hP1SDWkauqiv4+n2MS
3CfFzuH/YDETRKh4EQlEil3BknF4uBNfttYRjW9oQmHo7fOHbgREprfFGJTxWvl+
Fb6NvXjDrSjwLTURZgsgSbxCqfbZ/5J+LCEVltUR4OXay+ZT6eT9/k1MS/pEPOFi
nEJ+/+xLnwf4aD5M3dtorfepyDF1WC87E3yWDx3fE8468g6KdMsh8E8s0mkY4CP0
fKgghIk6nQFEgqyG9QNDjnpmZygX55EdOkc/FKTEd9HL27zOWUkblGxXAskqVi9K
RiamScNDOz2+PagF6gKwHmtQTZTFoY+t87xIT793NhHn4SXPbmbEa4nwKx6hppBb
LjqvfIZR4PUBBXpmaP1p0wIEPOyRixlYd+i2AWtb6HkwzbFfuvb8h9SR3ZIVAgMt
wIuNUN82QZGmscveP6YPdnIu9+5VBNinQyZseRcmgXWZdm4MiqIU9ZcLYEy+zwnN
0ZrfOFr8WNxzgv24MKoqc6+UnlNNGg3lrKPhYC2XqWpFZIZWO20zQvAZXr71chGK
a3meV2+C0R53JEGXG4LhHqkyEY757QBsrOcu1+tsc676SeF0hzACiPtkORqVvRVW
yWTWht6GwQBH/YQ9ju4hbXMZifc+Mutyuojcz+NQ1p7FHYUOswZ+/4lH70UAr7T1
/K5PgOUVLONLkfskaAQ0CtZ7h05PbxS3Q3lPgqEUxJY5+ahn3lTDMRalHfSpQlT7
0VZKwpH9dSzbncUWaRVOVzXy5PxG99WvYoGVfV6anv/S6dNWDVCicchHsj7bAE5U
gqRpsSaA8kFJ4wFxPB2yqMkDJcWa1dp2ed1pE6P/zW8ZVJ95ASGwIBTsEdI+Y1el
qBlRwXHelfP3pIVNswqzCRHnA5taa2T1GTp3+0aslEzyqmzVDBddUnmYL8eVpOGL
c1/tPtu1MdNFVFnC2sMQNAh1sjFroCBbExcDNyy/yaWzgHHMqCypx8OzyULW5HPg
Nt+qN8jJ13qDqYLBpB/9JxBABiwb5+7JkhQpAjYfWATga81AdCYr8SU+zy3SBFhl
fIt4Fs7Ogj89O5qrQ+3jMe1tASJeW4NCJahF9c7phKHT+4jd9WOkk+ld1Y4UOwRw
CzbdfEmiME+TzE16/P5ujgAZAIYrBSw+1jpHM5soIT+pbiSwXad30p5fjhRh40uq
hGyYaBmpeM+A6hvwMuQsstEPATL6sSkNpv8IAEhlAjg0KUXCU7+kw6p7j24UmPNh
7y3iOlY8In5udZbhsXO//i/6ghR8D46jXKxbrw233nbmYzhn7nA4XLcQIHx/EpQN
LfIyoKvoGAklzmsAHde71cxQNNDl0Tfr6GDS24G6sRgc8f6mwBe9ER5JHjfoUiR6
xtln5pmltCvLfYaCxpJ9JFXwXY8ohXeDYUMK5XcmMWyKmEMVrA8ClsKxI7KrmczZ
e1B7sYR3nl4wBIzUaoHw2IRtOx8AOU8aCJtPc6S+rtnMSopMTfTEjp/vdgmFQz+B
TXwLREGKbEEmiC7NviNZuFhn8JrhYMY54YhvkStQU4H5gCCAZU+Qi4dfeJ7/PWOV
7C5EJvKAjRSsB2lkC7abE4pkxAzusU1kgQOTeR7Se4U+82SMg6YOq2CxMmaP+40k
kfCKGEisThtAAp8EaDz6dnhLw4odoIKfPLksMbPzFEZOUv+7a6a1NvARp25tgHZw
RDN7VbNm9CgN42/BGOOFu7fnLKGC/eMTMUupq+KOyTcQX2tDJMiDeuUTmfhyM3Hc
BoeL27rN786DafB9CxrwnGSCELiN+aoZj8PBLk93oY1nn8/WJCYEOhZrbr3bYH7X
P0vcWPO2rnglVImVIalqoYazOHXVOl3ytohdYTiqVJU5ZDFID5HbV56eVt6/TJO7
/8PJ83YNtzOWCYBLXepM+JrjmSTEmwV3fjdZ5O5FCa7w1JVBVJZKoYZRmm1iTKA9
VgfNoERsLmlbA/2944EofcM3V8DzcomkULhQWO8zyZWDccO4BQGFeuKnDdS3Pe43
GLoclxb1uWOplyhCJBFCNEQhk93a/sNSGR9p4UeMKauExCEjLTOMj6g/qQnql3Ti
j2seS+4NNf2jgjWnCut68deJW4myUK/8/h/yhT8uNM11SSHdXI76GCkJmM2fk8AQ
u2kraiAvkXX+e0eOueF5FBVQrjY/DpYdzJN70lI/eVcXzsMeGFddVZ4V7wr56cfd
YtpJkq50JBObaHWeUhcq1M2wUbm2hm/m96Oaj3f0tS0tF1W8ZBpHZ8sXCNRD+3OO
cygw/IVG/8nzQ0RO5rFzV8NG7hMhgWvKDic3dViPyvTB3QQVdyYdD22krJhSzuoq
k15NY22VVn8bd0KG/wTnwE/uK2WVTufTV3Jx80PZTVNPtW0p+HwRXWUt4vC46Ynv
NOsWAkmk9QcbTm1ososf59xoITkrmBApqlm34jPffsL2wnXWicuM3yThHKcoBeJo
YKoVRTaOTt6lnLVkJ36UT09o3ho6uJ0zsWLd1SdFX3nmWyaH7lY0ATUFXF3ctROb
0RGU6HPj4ag0pgoAxZbj/bT4oKRvEtEAoy3UXkvcTZXCOdGiW+/WEfJFj6Nju6E6
AYXW1M/QM4XoF7NrLG3mVaelWU7ozQwWK4mdZ4EWLX/4cYYtqcH4D1LbyYmTIDi6
e0muMQZtIvM6+lIpmN2BoZJLMIvDyt+fcLTFuqMbldrLEQlUS8givtKwisn7rtMO
xIJ4gy+0MkZLaW4BL+URy2csKJRaJA9zKhisSOXwqLSvx8gSasNNOQZq8RQXY2Ej
HExHEz14NsVAs/BpB43s1SZTJOMJ/YMmHZI++mI00hxFZOalKb7sEK5WH3PX8Dab
weNkbC15OnKVqsG8ajwxOLeabsmAsbsXj5x0A51wIFoapwncRP3PECfZc3mp52Hg
3TAqwp+XgXgOcfUTnPZpZcXjMMxDKlX29mGyi6BkV+k1UlvE1T/51CXz4BmElHj5
WvEwI03OKmHM92yilpwEx/Fly9gEOh+3vP3HFR4jachsI3jI9S0O/46x5FHWoUES
wbXfVirey15KwfAj+JEepb26/UC4wDwSZc32kbOniKn1GTmCwh5gTOrB7/QGp3WQ
PL8ao7H2oL6XT8bmAy5bMN9hN9YQ9RGSvurLNhXaoLpNMzvXGzEWiH5UEJnkVq83
cFgY/afwTSzVNYcLzz6zi+8gUrJoXwqeRzUSNjw2QIb6mcRX0JmTF2GAjKmkkvwX
bL2tiMjvoSql7wg7nwrLWcNu59rbThSE7aPcIMsgpim/62r9J36TWrqSa9vLE+6y
EPe5IC2eZ+kDBZe+BLoC7odk+p4MCypZMdCUwhgz5uymoE8FRlPY6YcZ8xRIZ8Sq
IRBMv0jZTCpIabaOwlWD7b4FIRgnQwO0FVfn+gnwYB0IdUbn3s0n69h+FuFkOzI7
PVKJrbVEsr0j5Roox6ygjZ6kEuRFVEkwufez4WL5vrb1WQdTGINZoAYkZdod2DMX
Pd7zCoePOW2XsWnUgh0HZV8SYpMoe0WAFD1fcSjXBC/NKDFafygfDqH20rbI16aQ
+DkdXdYDxMdcu11oqm35SfZ90AL4y0L2e/kT3sJQYadyLjDjasBdXVFx96Ke0rGR
k7xGdz8fV9RXOwrysLid59zKvqH8fQJFF5hT3k7ST0r1g65lyWUko0k8s6UJjVH+
8dRIK2zEv6L1a834/unzCqAx4x/Eja6+V9lE0TPiDJe5u2uXJSHAgikmmL4rxeU5
sSCaLgmNUzfDbCT0dHi7OvtyORaoNQaS40dD7upYFxQ7gVBbciSHyIy0Uu3WGDho
1QfP6ocoXusOmT7t85wYBEeICc/0z5+b5UhZBABdkWh8FfDBkxaWZOxByTgWg0AM
Uy8/BjYTHuTmyRpVK0dc/Ys4oa8HMU2vnZvWoQhDXdiITxEqplC2AdHEYhhbb1Uh
1+vKx6vkQEL61DyHI3p0fI8mEpv+FWhqTGuMciCVGgjhJr6Oo19OzTkb0MvfgTPq
YV7PoC++JWdO8mDmtqyFf7FinGuwyaUH1RwVaW3/yAK6C+oDYKI/DDUmjbVuBXpU
XqSWeLyAVa2JLICFUmt2DH8VvmyIB6/mejlhUCAYNrjc2P9MNsiuG36LMe10u8UQ
QC17SqETdm4fc8jb+NTEfQqbpgIUcIx0bGqnI4MA7qpXBvVwzp0RowxfKeOkZZft
t+J3VEPopvM3GCxqCT8rNy/2+/txA9/XygUv5iNSdv7yUFnaOmjJgM2ZzVHmOfi5
LIhn/8RHDeUSeSwX1fbQJVcFLxHyq7AnCM//MvDh/rC0vJEMAQfautl4sOQ57qWX
sMyHPL+guZNzDaCHGIEfooVBlVOH3Pz2/WFzsqHCE0OjfzEKjtgcrECYYgvUHXgT
8ki7UUY1jcyBXUTYMq2ol5/7ZXLbRH+jdx0F4dbi5DiPlqlXYUms1oDhQSxtO4/y
fpytEiMPkSDLgmyUYbTNGdB5SPXlTctRMjlHqLzxCAozXfz9f1o0djRoSjicU9pW
2gHRAjNwipVVFrq6Ch5TMOaiDrUTqTyQyMMzksJyxInu10mjbCS+NB/uniYSkchf
p8/MtRNYwE2hLnOKQnh9TH4NLJRSCp9RZ4lC8DNHNOcn8YHxSCeD9BXVWYPHBACL
dU8wbxHImNuz0v5siifv/UwLoEi/rvW6ztOGGI+VcGtIT0oSO8B2vhW3n6DdqsXG
BiAxyyIk/OsfQT/wLrP+XlP/aDJ5+HGpKQjV3hEkQQu1WNqkEbH8T65TsyK+UIUg
2lzkt6vyvArKaQeFwJEMuIc4VZk6qLxouVToNnM/sslWj44KFJ6xDk2yF934A/aH
nkMdknDErbi40x5k0djJUUoxlEzRhaZYbKwBA/BtRKkiYqkALZFGMQ5g+1y/ibwO
PeYgTrzZT7Wrx883c3tT0luSZFtreHrOEnEMuN5blWXTjWABNUkMAXS4ktPazGgU
AkgC1iOhbszFSDVmIp14ZDQYop7wPTRrrhkH3J2hjnwBwVyVxx+nJ5/YstBU7VeF
+7l8r5OP7BorsumJxj1KHLcCGvUQzGDS46UONoa5zDNrjQiihV+VBPfeN5NGKQnr
JjkdnA8CGLu71KHDxgiZc9gDL5VqxejdNNJFf8SETnzdc2p9sakUztGE3IH5rXP4
Jh52fPWJax98zdckpiiLhW9NqMZgJkAfGs4+m4U/Sc085KUx/HfELXuBKmanhRdn
x8oOqv2Jc3ixgyA/bAa4SmAOx8FRt58/kXlDAwTndOvT+xK62kJtQctJgAUoisXM
DEFAGSPTSqqvKau9uruA+muelHGxzXpT42dzZaEdEdxJscSZJNpL1W55R+ELzoSr
FHHbfzUbQq+AcMH0e/Iy4AFe/iGzTriN7Rx7pjgnkJUmTVSrLwzKYD0X82ctYg5Q
jwf8fRsu3VB4g83B2qwDsO0B13GwD+eato9YVLMyyMEHlbeI6yNWHLGxzMVehUul
Q7PEup6UqraAcUcmBBgldMYq1e1ssY1n0bLnvqhzEShMTCdJaXk3vYx+bCr7s51G
P0z6SMUoay58DPJ5sY7AaI1h3je9pPlyI05ENPsYarQwlnoS38uAH8C0Dko5zwxj
KSof891vQFhksrQG9RJPyqMbdABV4SE+2NQScT4gTsQFmlHxZYHp2am849vl3xRp
CU2omqoWjKCwS9vTHXNz4+ifv6h0d/1JQ6rCuTsAlEpF9FT496ssA/O6zG4euJi5
kqsowraLf8ODDy+k30+Hu8TtGK/xNbmwJlDz11iI8jazHoXHmE379V4kBU8+ehMa
iIPvLsuo22xGnMVL9WTFBLKol2dNmIXUUlFqABHiRv4TdBsGWXekvV5KukYX+m5v
3dbnnlEhUJ4/LVkZI6/0sRZ2RFs3hWy/n0BpogziSfJN6ALvsgUJ/EtvnlM4/1I7
BcVbDc1teJ8S2IMSRc1yMhqpNMe/prSa2eoEy3BBa2uVgiCf/DzRyq4MKJt57KVc
5FO05E6fHXbbFVotsQH5ZSkh0muCHgzsyBCUzVKegDl5uOgbWe6R4kXTDWzehgRc
GDOfzCZ8g+jVmxhyL0/3F2d8dnB7Y+mPRiWng0DBtRaaQ+SKAzyvJlTBk/msKm25
eOvg9Fjg1AWz0i4lEoL4H8KxCuTmANL7CH++Y37EZ2UJfUvs1pEr6AJKOIu7tPjf
ofnQmXDezYQVG5EguOgFwzVM7RYSEVnmNzS/X82XHnHvxfP5tr/us4OWPQxukunB
dQ0fWy6KZQCymdD6/BFb7XmyfscslGuJUm6jsGQM3zycbr+agO7bQ0JZXlMXyrdP
TaoDYhEFZieELBOh29XqUV8kXm149FhcLJuq/XVElqrqI6GW5aTEChogS37MEYcQ
TnvW+rw1wsfimrDBos1O2mp3L0YrQSIFU/5SnW6+YAcIDXcB9zt6An39irknUq2d
mKTLL5toCXoFL8e4Ir96W9Mh7zLC5cMTur4rrHNVtp8SHO0/EKdydSnyxRcad/nd
P9FLbpJTxMP8/vUYjFpVUgFSx+W+2BYehJ1vcPNZHR4+E98OYGiLzQj4bA6DL4IK
XCETokQQTeQL9/IIh5UJX4nZkyRroN4N3OaHJdz/AdYF1Hzksojb4+3vrEi0/E3B
GgB9iHwJCnpkqQtqGSS5VyyBOvJ0SNLcyvz5OZ0jh9RG/bRrwmDe1mAR+LhOIH/5
nj0KLJJa+Co0JF6KJNf1tsq0kQ/sRtMcO26UJbs0pMEiSxm4jIgSpdatqXAdYSny
9H9bZkPulg4nM6TY87ZZmEprqW4rR1AQe7GV1M/+WrDBKYifXJPJ20YegoBGTXaS
cmgUqe3dglwG9LbFosC/H+Tv7AI3dgLGaAxfOowUkDo9OyRS7UZxudVpipEiYGEZ
ke+yAWfGpObqoK8uIm0xFIL6ZkA+VxPviwqDAwbnbfTpueN8aGcds1hOic2x46PG
AyYifczLKL56Qgl04PcuBZAb8Mn7rUptXDaBHFhEc0uF1g4aQqp33CRCs2vs9xd7
rFGk70DdDvuDMNRJRbjM66uGs2vYGHJjQjKHCVcPMwQ4jhyE0MVhXxybOBCEVb0+
l8V3428IMvIVSQwTUq9acmY3KJ9d3I7UhJNkPdp6QU7ogcc7cEykeny5CiYytG8Z
ez3cMnCVlFbKtOu0mrrU/fiAGNk2R0F0Xw6p+iuFAPdVAIeYNkhuw0fm8fnY23Yt
KY6/+/4KN4JoM0vP1RTpdDf9MJowIoHSpto8OgqI/Wc6Q7W700oF2DznG8veqkLF
ffqUk6lZIz6/aCtQVXvkqGJqN3mKHzlNE2sDFdV5/S7NdNl+OvRk6B3biy5zxa6u
8wfgyoAAdlSzMjjuNyDAuquYE/4cH2hgl6yTfyH9qYraWSv91CUaLXn1Xdr9v+eS
xzjeJ9Q0EB5m0h9Ty4xpNzxlvnbO2gEo0dxSayjScFtcSg+Cp/041GcimQxpgs+p
8FPFr2betFUcQ8mycaKTUx8/4ra/tpErIbjFMVnIKtw66Q+1lRkwb+qxi2u1ev5J
pmUcds/qncJYgYv+u9uh2uRbsbBFtVZUTh81DzCRaGHdmWP2hR9Fhk3NqYY7zSnC
qtF0mdmONM6rl1tk6MMyYYY+DApnL0xZYxemzDu14MTfCAW16wYN7xAWn7TqWjpM
pQ/qA/q+xJPBscGJ4ugozsbtgUkjgLk8sNzQs2gkFSxCzSF60qQeIw0ZHltahJws
yx7lFWovTgP95G2XwelUbIDA066KD6haHIq4SetZQEv6gtkqM/gq0tZGuRfgl2lm
nAEHxyDlFPvGrvcpKYqiYaXSqMv9tE20Kv+DGQ123EKa5QIFhLmJzRppYqhYJ4tK
6rppXrMvtdk7gNDpqC1x5eUfGaeY8PiXwE9gQeEWJskwoEBdf+wc/DA7DRcFDtXw
GJw8o5duv0xPfVFPadwMi/AwC308up9OjHJMevaXj8+C/UutIZ8NOLU2M5g4m68r
Br5s3mZllGRZnxLD9UpRlQDy4EF3ck/QRb7m95XxlN6at2c9c33iein+tLOxVHD7
ZcZFgGUux+8MWAlcsHoME2LvVQTPRqfWh6Pz7XsslwF1ZXByD0qjdAA6JtKm/9U8
oGosGAcWEHboAo3/cuRcVuhkWejitnBRlu6qMTVZGw1fV6DyuWfLe1TkWVVLmW6e
WlC9eXC5iPH6/LdjRYh7F627SOcQkNJ35sL1Er5NrmmHkvtSxq3RrkmqWurCptdu
NZKIKbnwudlBzxJUuLrSD98wTx69BHdT0cu2c1Z2sP+IK0X7w2rZu4Zea/zqZ/RV
b/U8WLvx5N8z4syR4Qak89McQa2qwgToJmCn0OMiATOeCEGyLi38WZlk+GPsUBgr
/XjqsXTTYlAdVcALepU3bs7bPIqrvVF8UTn8o20l7IXx7LxfWcaJOHgUIA3wm4Du
evuKgUv63uvEy74DLMp0GHqlBW1J7rd8Bph6+GDBM+yC4wcBPDhMB9rec8The/+9
mC5jT2+5mKyVJ59Bg4LxLyT1IqqeXnAIjFpaYUZlNdQ/sib7Ja3D8pYeg9MtB/6N
IS/qGjc3a9cmq7wOBmGbXby1EI/r59caYAX0CsOb5LKXHhsG67u823oeFVhIrYz3
8ibK2R1k9j18yazcNXzsJKiOq6z7QaTUY7gJtTn7teXFQKQ5mDYz7Ij9y+0ZraO7
WBtKL1OFFZA4ozo3CXKFnF4n+GSNnR66sUo5TLXD460MyWvysUEPX9PCgZSq1Pda
6BbmMAVJpDOqqRpHN5QaCzjhghNpcBpI44XiiTUGlO1XItNRP1pBNKRLSluqyPJE
Nv7dJwDg1ADEX40ZF8jqst/LLc78i4Oec4aFsTL33u0QIOiecUWdSfkKqkkGiTiw
j1FDbADeBDb57wDtkdSkp8XDzXBY+gflTDjyolewEyWY3ZGChHeeWTY9NX+j2YbN
Utgf6vcatth4ZaHcmKRX9qBHhF2ok695UV3SmGrxSg5UIHhnXca6kZccclxnF19z
9lPhVeykwJ1+GE8qZ1vhJLs0JNhh8I21c6ikD08uzBuh13kfU0WhPVC1TzQk8naJ
waE9C8oOCuOcQg+K4elPpbeD19KPW5ofWrJam2hqWoX5CFNXDqGtL7BC5ePYPbpK
UjeuzOYOxqexa9SijNbl1BAU71JJLVWYyDP5sgAXKc8Ggsm2tddl9C5Yqjrp7aV8
sEGpcu4/rf39j+gCE6RP4XwlRqXrjIv71QO5KQWJb0K0IWOoQdD4VVMEP/aSolYT
+sjQvOKgPpgGsF4J93XpFjggJQo1RJzFPpCCOCmaGWAMwUSVOVf152F6m1I4YYUb
x5/Y5b3OCs+bTwLl44oabXimGZEnVurzZIFhq6082b9RHY/eWyG6jK02/nrNCsIi
RawjpE49eUIEp5ACd9JOzF97oodbmbICOBx5Azya0OylFOBwzMHeX5HPWC1P2qaE
NHPWqMaR6pXfIeOBzTS4Y9JD5uSa/BZQbUI4p9pdZ1HtG7voNgDB9DLKLK/10pFY
oPLlB2urHv7QYIqZl3JUmjL9ugnsWCdGXW7L+HOlzmNAVGYwL2rQPzZOOIfk6/Sg
+gj/0pqLGSXTaJxl6UvXUbTflmmLDGp2T7r3o7hWFxrxVh5wDcrF7EJ9OwLhAZjx
J4DvZJrubETi0T/r0kaAEvQUpflYhcANbPw218SsWI2Jac6O7CLTOQLAulTrDpdZ
neOi6zrBdALkhzPtsyaoVdPMXFn0IsNSt9bykdrpnG4bZXCQ8RAncqpAWHovo4o1
ys2c33hxLp2+zlhOa9tWcyJvqN9Gsz5jDBIYb9BLj4byYRVGp1Ci0vXShNcjkMZB
bl7UCybyq77e6ukhhaWkgNIAVEbRpFNQmUL1iR2pOfmTf6Wr1DyHuS0LK40rjh3i
LpYoEYjbPcPIZ4KfQ54f6Nx2ZWqlvdt+v+oYT0vE2Sf+Ogs3vBdx6JHjc4YSOwDk
WAHpgb3knNm4XOxXGclzNEnfyOpD4QjIZG400O+zqERz0DzpOjPggY8y7Eskurei
amTnF1AlR1uH1RKQyZKjA78Udu9Ti2jqZPNN/vt/GfWJL/BZd2F7RuCzGWJytYEt
zC1BY2F//4fBGTIRdB2XzZetfXg8IwlEEPfU7kz0qfiMFzH3uTLiwTuNRVx3hhKM
rbtOrBrRLQo2Ju1B0c6VGUAvPvgMkvwkaILr18TGYsMt7Acr4YFlDyJPbedf03to
FVMFN/DBeF3kW1UMZ5D7ROebZngDfZf6d5kjOnpHmfJ6Hp6Och2ujVDoYuUgZpuS
1uz4N2kVH210lQwotWXqVsri77TpdWALw7NyuSiDddE4kNMCJoP5hyEfv8zGjVTW
nhQjAV8fwqkJPyf0CEJh1PJ3sWSgjDfjRVyTd6I5ZlFcEE/xoNKNynjCl7gOhrRH
6v+5z0LEsT8p67Cz1Ruc/kVLf+vEZZUkPLZqIMZwVPuI8ifHKR2s6mz1aAK32+tl
M6vzx/M3JRF486tVkBWLgHStb4b114Qv4iDk+94kYTVXdyDeO441OJCDapGU3vOk
6FzFftndE/Zag1YBxkDbXeaEvnteXQ/OYp8dL2Q4r6bC3E+s0m4HakyyS9ZA6fET
gKW1Gqch2T6mX6p0qsVTcW6J6pdRZRKQIkYVo/pVbmO5FxMn1aCskQVwjncgScMn
P0B5SjWcc/bK3UdTaHApVuHKKHPjOTG4n+ElnPLPNGlhRfT6xTZjCqcQI5UzQYmc
IK4wFQmeoJXSf69G4BVJM85M2zPKYHHojqRLzv8iwCM4y6i66PFvqrX7t19GCCiF
OiwXMDshAGyPWGe/0WOM6p4vtztwJ70cwxxIJWb+eFzuei/fv4uQ35IEadqi7GE0
8b7c9EDwHUM3NwOJM0a2INS8upIyGe8a60A+dT2nsniGcah9DeMDrLpfAifFGSZA
giWVuwQSTkLiZzaPG7/SH0h3z9aCRNuWUSM3Ta1QhE/WWWnBzJxwY9clqZ7Y/dQk
ei+87zEICQFomQ8O0AYToHWd+j2c3eZIscJiOtyN22aeSf8YvnxgH/X0M8gvD+fm
e/NoQr8aecxKxko8W1xFj9XHP1RmZSPbNrxhcjRythGHwjxhivBdUe1sW+alXANI
MtM5TDlvrdVTqLQlPGjxEzcoq/b3gE2ZXzMytQeVmCDDhlAPVXp5t/4nbyM/fM2d
s7ydRChLH+UWvKtrNGgliKOHO4AsoQ1mqWfFbqxP2KjNr/J9Ghz7DSgSoTRswlRU
owsa209UKT/3kXWqzF7b/defzpefedStG9botWka3Ot3bPIcRRS6lABtCuRq4pvT
ptp02XocyyMjqV1aU7msIpmcO3Tnzz/5MQailV6SViDu93JP/XcZSUFemuqxzR4D
TWqntyH7vYGAEd4TaYQz5mC+UHwWiLsxP/c5T/2MR3dsymwP/eY0jaShgEwJRG/Q
n176/QDziXkrgnKwhU2BL0uKjARAcTtCe+4BfTSqefl6YxGa9zaoSnMOlGKytflJ
eKJ/+KTBz7q6uuhUP8w/1+E2/3/YsDmCZAGycvLQbzP3gy8Aazd8AXcS8GtJWQPg
ZFUuGfwIhOrXb/BmXNjIvabO8koPaMfAykQnTzuyZPdTR+TV1Lr3Qs5f7UromsPm
LCcyZU0bRrzIFO0DoZLoe6HJalbrYaV3i1+PlCvcuHOPy51+mtnQrw3CT4X3grem
EmK903wX9Megci4DOxOsm2MoRKWoHfq4eThDZ8fQRm/6+ZhcY//cMP/qdnkKVJ+n
IwHiClLFAvIkKLAKPDeL61fw89YEIAhZhxQeKpLrdkf68UkpFwBThep1/o9H4Xt8
6RIv8nDyEr9Tp8vA/3pVSJNKWyUzMV3GO/KRGbo8TIOdOIvpoLuS5NkHQrdJUUTl
l6g6m1x96YlXnK4flVD+HNQMK+95I62vdkzfid31H5LxYpqVcpGxm1U5YqaOfspF
cLlf2tF/xQ5u+FepofPhPXNgRfJuqBFUhDkn8gVzuXsvlpQFXfLb5kD1mpb0M+eW
e+28yMzI3JlyS4THhh4JbHpYqJBxH/wD5m34gdOSh7L7LX6d5CnH8txnPUemd9Xh
gIrN7YRz+X4ZEvEKtb0MmAoMhWKt8GnoOH5wak2jYKWNZzgf/k6cVzG3bu/8x3EA
qbWiyxBKSxeB+iakvlwv6SAvOMRzBmiBdiWsPBUKMpWzA6FU1Ld3g5+JME3GXi3G
AegUCdHTm74bLNXdRI4YyepofgaxtkC40kPeeK4AjJCz6uIRvtb5BlWcwtbJnLei
2qcOPZhXb/JZfkbfZcsefOdaKbLjuiQYMJuAd5R+ZZAcZNwJ/Vx5gL/IVgttUhQ7
UHlAc6q6zT04sDNfznTBdZ9wq8jJyM8F3W9/nFh+OaE//Dg7Oye+bYTuZOUF6ovf
AcWppVIQrgJKRnc9FjpuNmmDbVfvV037ot9VgRnryHpLQNGV84WJDPsANM2ilIwR
63Mlka3rxwtK7FPtVduhtku5DZQF/BT9FJmHizDAft+zK5YBIgGuP3wl/vzr4KMO
MNtsfZIR2rWKKO/gn6GgO0ey1Jg82zyipKiNV8F/SdbqtXNMKotjkdGdbYpQweZr
JPEhm641dfC/ongmbDppRfdboKsWw6x1OUAxRFWXKwQnBczZDGPKxm7DP3e7jvYV
WZ44n61DtzKGTCs7O7kw2twqf4l8LttiYvD4Tzp0F/2tBOgNdf8FX8L+ACKLAnvX
c+FYfmSoLgpobuGYMa2ZTLNh2wudwJUMDBGxeyonrGk1b0qWO8hantg6SUZGTdEO
foIoWRn6/1N+42xWBfDa4Jw0OvAjhfy9IPlPU4y59v4j0F3qiI4UmtdV6LDVwkfr
bvQZTHYLaMsRgufYqkgMBko1vgbAz/yHdXxF9d5NVQTUpVX/qC2hL1ms3fVuud30
N+TECgMUDOUJZPfXR+tSeJit8DpCJA6EEn80jwqQRx4ZFC2NHqaf7uf7wn5rhP+z
AWIRAll7V6qc7TVxU227mdpfYfknmAo7Df6gW+0htCk+w1tQbvGHlNsWOLfHUm6H
+iWp6Fgb0BIdOibLRBx01MWhNqZ2ElkT5x9qS5AvwqG1mZpUerDsi/iAJOGXVNJd
GBWlg0uHBBbf0teVp1gQDGXbVUIt/ic+1UvizcmwUMgG1Ob4ckehEmbFucMxlm9/
ba/0AbCmrTcz4s9LxgAFwnH/z3LbqHsV073pGh1usapBVAkA/Nomu8C+txSsi/T2
CTUsrCpQ4vnPnjc76+5vDU+QDJSPzKiNiP3xwcg75OA9dXVRK04DSB0q6PJcoLbp
1UARZ0c9eIy8gxbLv1TCf+j0+OOMN6UDF9XtRh+ytglSQsmRWIR3Qsgw+CZfKPKh
7suIIfq3kOEIJzuazhLhqIvXOlMyqy+u5X8OnF0GYYGcqu/JusB/J+E1FRm2tfmP
saTEzf3jFUOvD4MCfYEBx/5Q/tBG6R9p8kFeIaO2JiDNdRT3GV7zKQxTnAIAy/M7
lfQpBAPVMFh0PhxWWh+3w8PBeYqN8esPNwI7N02100i/N2AkIeGqUb0A1YBOgwNv
FZQI4Rl0VaGzT/GqDLlQEXCxpgbcAtxdxU7Swto+POJqIXm196GHKz/zKFJUDRDS
8N5Mk33vBOuTRZsmDbX4D8sYNB6/52t20eV1R5iUNsMSKJQIT7Jh3TSBIIhcOA7p
nnTIeVUHNK5Z7kKIqayYlAhZSOjX1yFf1caY5QzOrrmm0smsmsvwZ4Ezui3kS6h3
LTGB5N/5la5dlkiZ0ghpL0+rLP1jL4uVM14cYg4MCH7MCyS5soh5pI6wt+dSuC2+
WS9O0YEsdQRvIGLJI0uytrHcS4ZI5cxV8BthsdMgk683D3XWYsWbVPhxkwRY5nj+
felkHn/b/5yE1y9GK9vKDZGLrVQfDnyDbzdZlsYh1YZ3nPQacjrszRqbmVmWRSWf
Fj2qidkqvZXcmgJy9/mlKTZC27rFoMotsbP7chw3kcY2kO8ZWMV3dlt5f0uM9PfF
in3WJ12++ZFsV/nwQcN9beOpwuwAvnLkV+LUTzF72NVA4QjtaCpdOBgUXwei93OJ
qECs+IKbgVdxCwfyhyhwBbKilJ+2TqdcVky51/xrO6l1NHJz2RIlvB4k3OmgPNsC
C4ESqtH1N2w34wMZ1IoohRMqxABrw2henJc1eCw2UYtSGtmGGGy4a0Pf2QwRFc/J
ajmljbZdFjddCxgz4CB54L+AVS21y5+GPuJx7zA4OmXKRoKUeyLjl3PtSobkSa0Y
//V+o/ic7STpeid7cdjIdZ6ZaVAkv6iGCajLfAB8Ca2kX3gl43GHb6T5skCcSsYQ
+FL2IaomSNebk4kN/JIKSi89tZKfL3FvfyTfFdYGxuCe7gmhz5vO0vTEdY25SKAG
J5RwZ/naKb+6xikdSmfIXPCFHtl5H6aa7X4bFJFbR7evQ0oS5exvpmbIVH/ahrRF
7WWS9YpaD0a805EO1GlgIUsUm6bpmu3VICnZzAFqkwFsFOW5AmWHtY0RAQZRbaza
Q328PxdSPEEA8YsrjdgicpxBhjO9bkTYBTKifr9jP2tz229NX0F0W8mejUJHHlJB
S8QOQ3XplSDogA6zfqJ2afTRTunWt6aHfncKwA/QXVXabBzCoqgnwiJheGDgz/rk
OI1n9EtmnX4AWpiTFqh0OFXGbQ0dwtxHOy+wxhyIWGNSP4VKfIeEAMo3wGXcLu6z
bd3mOa6Aj3lTuVCeBiB8FcnKwDPVngqX6UGMNMCU727GtfgBcDVKVvXyT3kD6Gyb
3+rP9j+JcxuZO6vtaTbOC39lsDqK2oEsGpBVUsRN/KuRCgCDjSytwzaJLmQ74ot/
e3x73PAOfqYLbSyTE510gpycuZZhDwE8CnAdDePU6nxkMenIT5fajGmDPUVDKssY
IGrTiNUJtsAWqkhoXK+ri08Cu5Cbge9jKmBulIKG9JYKTsn5zWk7uapiGL9B7LFG
jVb8syW2Ty9gFwopjhyf0zNvGGPClBTSGQI85cb2bJGLRh6nvUTT/HIxwM1HLiR4
K7J4VET9q390aZI+T7JIiscUz/pkdpUDNsWPWjGSrOuLFgxYkr0xC8nmMPu1PpPh
NmrfWc70yXX1kUiSVRLBRhuRF8IhEdPUrGSxbS7XAU8yR3ezjq/NiF7Q4WAeg+va
CRpJNu8IUXJ78VMQa4Du51UfGX7PmEU4ZCqqLoC/rrtL4JTOiXn/uyZPjfwxusNU
bBkYZfD2iFIdDwMgwgv8mVHR3zxuLWwG3gC5iIUtSFwcjhvkIdMWcx41/v79GcRT
BOJxlVo2ufVJKPmKLNHIltZ1IDLrxiVn44EPyQsfOgLww4Tr6sj5X8vPHxs1XFtV
GxQhJYg1F2C6Ey8iUFXmXDfxFjUPAIJzCYEktJ0+WcJlxwZgqWgianb0DGPc7Jr2
p1wF462Q3HbOBjYA4wT6cuQYA0cxpqcc2OIb1IdUdTL/K9Su/SzzEDxrLJ4Wbtcv
B37+uqGu3APEJWr8WQCoomDm2O05LDlDvi4U+f7XZKVXkoa+2H4HTfTN8+zGcSlv
pC28I4U/HqnIwLU0aEArujmyrPYhbG0GssxyY558d1Gvcr3wmiY/4t2lDahEVG3o
KyR/rIne7404FjHdXQvMaewWS6+nKbewQiD6R9PTzoZ/rYWpxOaTuoFrC/WSCITg
iH5m5PbY/1vsQvFiB+78STYxKvJ340XHDWwbuD0PSwosPJyJbZ+A6DAiE3xz2hoY
`pragma protect end_protected
