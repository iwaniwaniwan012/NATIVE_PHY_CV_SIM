`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
K0uT2tuP2DMOJ+1+4Vqoemzm8QPsi8FMo1OJABmeY8ewjEkcKG0rEgbuLx9Gcg/t
JDhl4jkTo2m8z/FGqM7DtIVSrXyH/DBbNtbV3uH4wNlLHiA2m/60tnAt7hYmrSSC
q7aVkuZasI8lfJXflGhuFRGXaIPHdCMAjmGG3eq9/n8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32976)
IP7GDrFjNG1DKLHAFtovRhs34m0mzJFs1VDqAGqAbMFGrnyTjcXpeaM4gUMV4vR4
BgGN5X/RY+qcAqasmiz4Xa6eAwiOV0w7knxGZ76LbE7GYRf3C5r+SMLtyOn5+v4t
/BMW618ZH0G3meaK8Y2oiJK349L7SqYWVf2SUgSbE1VmYDkCIOaphWw9lpPoU8KX
hsdhfaIdqRqEvfUkcABPrpVBWnn20LblIL1TxsUVicS1A5pzBOXC+jOuiYYMudpw
o2IeYL1i/tXH/YvWQvlAwQEgqw7k5LEaoMM4vUhVyWsxfKLT3FJkq8FNQQh7l+70
OMtqRSLIkNbiDFEY+hil/eB7K0/yY2TyWdKsFFb6jf4QJ6jBHwAeutOif9L3m40Z
fbrmvlhEjiDQhVQ6kSbNzQ+MLWd9OyhSuU4NSzHUVSrTpylkiGScktBIfFc9rZ83
X48+TrttTv7t05QGFZ6mDnCNqFEzemew7JEAfofW867jT17O6YqHcG3Nyw38LGbT
Y5iWW4bcCimBdNMHLDC617M+4qZYrwca2YRQEADYwxdIyuMcb81sDa36UD1SMOpz
oPJb52gqcBGAjWDzjNitxtpy7SZovLE65Rw23UWIvN4mXiOJX3lpUfVafz/ui0XX
/X270U1aapSF1ml4B2DyJ1Wad09NKwiJIw7EdIMjAqxF+ucP1cjI3m/qgMWRw+EP
iol7A7RD//viF36qVm6PnB++Rxq/pRyhe/BjO07KKzzlt8lp44BsyqpXOYgQ+l6P
dH/3RFw+bQuDpvIqWjlHjMyJZjyHowgaPRfAwpRI4cfQT42FpqckYqUlpywjmFCq
mw1mav6IUW4dNMeHtx1YCf8uEr+Zd/GAdjU7fLwOadrvNm0wa9MnCwpVW6b7Uq2l
wmVgp7O4DVprh//jg+csX5IURdnKgeiPMSMPIyg1u6j5bQti0Sc5l8NglA8eN/2P
X0co8viQL+3iic+RSkznV+N7n8GdBW4lO4+hevF1YKnHs7FMHVH2dK1RE10AtMRW
GT2YJkFdWt5K03/LzC0VvhafmxKvo6ux/5/pVUNu0HiWHFE+kRbyj7l8GgWW1viu
TqtcyG7a+LvH++QD9lvnvu9P4o1hCqncs8nxL6jfRwwgKGu9CrHBZrulWQmTIu7m
sL4l1CMchHmuKn8HG4Bvk4aC4G0PYBeS6TrLxMhMNSobAJ3tIDds6CmBFdJJxl97
MuPeOtEdtoDJVjtFo856y5/SPDYJg9j736z1aMOxR/Zv831icyI4Q08mYuhKNY4K
izj2i9TtJ6EVrqVK/41S4kISepPB3OhLJSukEmJwgNPA5GG6+Fo7ubMtoZi9m+7Y
iAE7YGG86SeXwevh7FT+pz2uBtizjIdPZf/3Y6IUG3AEUNLHwPS5HoXpl9nxNGc/
VDtCVyKf1w8HR6+ea2Y5DHbwZxzN08+xfN9SV6WuxygSIAhof4Copj8bL7bcdEds
9LRA5mOBmoRfXIoAScDOlSGXK83tkID0xpNOAZsxkVbdjMiwph6DSzyede1j9DF6
RldJFBArqXLi+WhhxMw1RlKUDUAKe1PRBiuXvC7an/zpS6aJWdiGUSRJWxAv53wD
0DINV0PthNE13hXrbzFCMhY0GitKaASbdx2/jzQaF28CbCcw2jvuw+iQExarQe/+
pDUkFc41AsVxU0gG1F2KdRgCwtibbuiUp0PfQGziiZJun8PO09vp3oEKam74NT19
YteTBVGWIL8+oRAttElC5gm8H6QBBfeXf89pnxuOJ+a0HoulEtt/vEwyGCZOw9NP
GJqgH/OSgDJEJvXAStaAKhSZlb4ASSgEpmYesNekXAAoS1vL5YfedGYL0/rUoYev
dP0S8roGaQnZIAv3M0EcWg++/0OCP/QrGpnCHYkuJbAu8VwP8qwJTnwiGi2SJfbb
l9blJnE129V3dbSCeeeUpyArHpo1tdQjR4vuoFXMeGg8oouFtymm9D0ayoLPTZRW
KQDQRSf7U1HItsDxXA++pqzVNeH8U7q24aJ5kjQWb4GknxTTwYvMCt/1fF3wiX3c
VadJ4xk8/obb91tSguyPOTUyXu1AwDTD95DDTuz0XAzJCFzwZmM/TIFZlzolFgOw
rGUxYsNNtS3JhwtNxC48V4Sf5wpWsIpclBMQIZunjMq7R5J8jG+eSySdlFmQ25vX
4I+iw9b7QUf4EdrEkGGokdEql7d8UyXPah3gLOV8vg/xc5OA2zLMV4xtYG391QXS
hECIffFHRP4Xz3eIb6KhOSJTDXsThSYWQVKkL9+O3l2lIktTfRnuEFm9i7wFQtTb
ErUTzYeQQmkv6LvzicEM4JnA9MDoPaQSSp0QulnLgVd9bxi7gJjOd/5GhqsBBPo7
BHtZWP90pggAZaRxsK2bOqBol0Y2BLDkwdFCRL5yujXE2SCUWGJggVDmSWchlepn
cXhJqO3PZg1KwXp0Sux2OGoGNEpWZfavlEWWvaB50HybCRqMl8iLPxzkbMSWGtbM
40HCUVAWAfXlUjtZIICuwoRwm+Aaob4KzYayPjA1Yj6GWYAb3JqIpeLibW6E4Snz
mfGmVO5h7aCR2H88yQKHp2DLUAcl58vnQifOpA6q6INBe+mA+VZGKiG/qaNp7OcG
L5YXre3T5DUd6FOT+BDXESdHG6od28M6pB/ccqwU/NXxrNOmftw3Qm17E/jev3Ld
IHd7bhYt3wB2f5N2YEaJ0Ed+ThFX1zcF3CfWiqpMeIeRsrhABwYSFAdu8hRVSJnX
wALPRnbEt8gbqo+PwP8eFdHe80y74wcScKpfF+qoxavrY9ugPAuBgn5LRIOinFAQ
bWTXXK/95/X2H5u468i4WD+I2+kq7sYb/wig6l+yEJo84zRJ7zj6abbanV+3MdFq
RelZ77hh5xCphuIXiMA9xMkPki8KW8hUsjejWUbcUE/xgOb/VE9+05WNFcl03Eq9
paOh9Yvd7lYOPLCSJ1vfZvZxSJ9wUgF24TfVahfP7q2YqJxuw+am2ld1e+FuU0Cs
C22aSH5bpAL9dboBHehAXyZvT+25MUp/tkmTj2ehFqK05A0/JBo2sQAA2LPx8tON
fC36fVBeI6KiCI2ZpoPvChREA3xFyK1Gxb20bo2wdYMonGuKgQbxjpN0g0tkJMwF
qI1AuvPEdPQi/CsDr+hUCoH9+7vMUPm9BgsHUHCYA58RdvMa4zcQFxabjht7J9JX
w0SGSg1Daa1YlrfMuFPEVvUTLeArwWgQyZjo5vfp0qIUZtqfVJV0JlRvOPZNInOv
+wCzfe3OwxGVUiPZfAmNOjECEFCTtXtusPikn1guiTzHsSKptsHRSQK7FqJfkBcR
on8VLBxQ3/nqFlctkIqtyY58Kd6OwMUnLUAYbEe0h8W3YaLshL1qjSxAh1kU1svU
vqdRKjsBB649gDNxPaL97N0hjPWy4nicgTIxDR1pweiHK1p5j/RxGe8C8Hkjb4Go
yQ6b/nXF84821NTokqJcKm28glW78mLDwF/vMDkk11T4VjtfV2MsOHq58taXsdpX
fpR++hKhoL/tSroHbreV07zY/1+wC9bEzQlvT8dyBaSZNVkcC0hQGYh7WzChOY77
rdpT1CEK/mtkZthwNQ8KX9TVFlTNs+Paoqr1gDzYGuZ4V31iKCW70U7N67rzIi2z
NtPSBHiccR1LWO1oHnbAmfFX1/edgA33zNuBpI2eGOVfReK62ViecnMqcBJrUns6
cca3Cv23vSQRpM8MI3paXaw9fFxAVeM+zhtN/PagN+MSouX5HPv5I/kSCpGnf1mt
KH+lSPuqwGeOTk/rqs1KlJe9PhL6m5wTUQtENVdiw8QUkZzu0ep2L7w8+OjTDLut
0MyZW+03jZAKw3AqDB+mhAR4pYhrVT7D62brqm0aWW2DyXFsun4i/ow+8OOBJBbq
TTpms4+kdtqQu2Tu9K1TeftddAXUzMVgKKfTCTXTB9/+wCjq8PzwKV44ZYXsBHE2
Jb0U5lBJ/BlIIOKmq+Iagg7eg5ybMvtbfD6TE6rUvAQX/cs+fLSxrBUu/tNNNkij
FJGINjGSCLhEhkDX1cUBcRTeiTXFT0iEEnqzynzevLQ/GMgxwFDL++4lkgRBSKSO
vltaNNW+JHezGoBPwXNdna61unDcLfwKffLdymK4AU/fkIdxy4F+ruLP1knPtnGJ
IAYwnmfKkvKuN5fST9SvjwO02i1J0lvvOIcnLN4vGsIW1l5DjJ5pySRAUjIu0cxt
XgE8C2J83dluO6qpEQMgG2UhZX420jpA4Z9giG/KFDCUp0f3WFqevv5dohVmFIM1
3+orbkV24SKM9423Mzws/Gh3FjgnkACbCsaUg+J2Wn28XdtcOMzsPVYVq5+O2/fx
jOM5o1KSytLVmBjbF1nMnJLYQBicYCL8WSM8EJ+QlmcRlild5MILzJOdVJrIuP7o
SwQagOTeXpUTkZnCep16gMKCj5r+3Po176NWEuK/MJPj62wTQawnxUhnsB2sl6s1
BL2VzkMG+H4aB6omLDMhWoLw7A07ChdM1/7Mky3KP2TVAjDLUK71/VazRRIgeI/7
nZ3KyvCJ9pzc0tSUBQJx1MGnUNpI+1rrMS2LHEvOIP+zbT+gk2lgIO+cGmsgQCLb
+rH8greDczT6MTnH/FvPBLtFZqK/oFK+xVoPgWnz/oLsABgx1hfPC0AOwg1BOk0v
VnRDoRhfRhv5+Sy/HsJvOORaHfTrWcPKy2URilJesG/Sh5WoDJ8QWHbEaIzFNXMr
J2iAJfvZ5yocnU+AEg6UKFuLnQ8p0NgEYonzEEjQkv8Kedl8SOgRDafhvzL0e+La
kqODJW4RIQie7rho0SVhbLOKknCCLCbdw0Sn4ovSRLJ4dFscafy2dVpGHVbBrBfg
xFlqse0TEo61CeTi6P3CuFNLV7YgMDGW/v4PinRzwPHLivYJbXAJBMlYWQOCQ5bO
P8rJ/ub2Ql3ZNoJnTvjM8aLTqTgJ9WM7evKVDfpp/EHZKsLI7Ob9OAI1NQmgqOSQ
qVG6kAUhTO0B/lBDMiB2DTrlAIx0yUdmVwfJLMNDGYHuUqXQy4jR2+i9rQkSRynI
AisyndGJbuY0bLIiDocyydD0KVHm/mVAPZbMlYs1lqQA/lgvYBa61adMZSsySSXB
Kfwtv01QqMqasmhi1GW/rD9cqN+ME2jJuWMYefyQ2q8cbKWnltsT6j6p/20MSXu0
EtQ996feQef0+dSif+A/qhJ60QxmDtA64boh0gH2nmTBrFpuzgKGN7momA1JZGBz
2pGhImRg8Eh4Din8PY4IihHwP8fGpuEQMrXZZV3E0eGdTS6/AAK6MSgSuW4Z6SMD
B724LLBRzmrNG1B9TTrwrs1cKInDpZ2TpYhiW3jttgj0GlzxlF/qcEQgvTEQLTlP
NmJLCuEXM1Qhs05wk93FKdItLosUtobX1uEK27PmhQz/FY2cmmrBQurdilnf1drB
SPRcUoqRyeecIoucaiMYOeBoIO9AcRVTGYFll6OSzsM6N7tO2BMbCcaFbcx81DzB
q2nQAW+kFDzRmMZOHoLPb5hjQskJE4sXmRjh3lhgpQ7cIt2dJSlZ6scDQqZDCzAu
e8pQn0EgV7HmRQYFD3cPhGdyW6MbGatkIlXpIITmGkn2mDhCuZqqkuQ6H0BuZg2Z
swEy5wFHx7JrABKIjwmHsYhXpqpGl+HpNydK/D6nA6GTYxAkDo4zv99/BGM6yx87
qmv9/n349gUXppk54ehZ2J5kjYFmSmA12MMwyX2s92wOJrrPYRsqvOugZmx02p44
DdcXlm01YcHsUUBSLU9aViuzk8/Ctnoc9TdIHLdHZJJDkkAk2cFE4loXV8+WoSmW
ZlC1xT+gsdmDUBiX4fYS523xwYnTxRrUweqHPBbgcvXKhb00yDrR9qutWXnc6TS9
Jzs7tTe+dVbsDR3Y7nOXcCrRGBdTD9/hpTyhApQgzgxM2OmN80FMwsrYa0VosgId
lypjCbSxVb9EZr4AOLdIDHGcLEkwYe7AOBTSY4RauQBegP0TZzukqQWgCLlAi+dr
SGPkojdSunLmpXyHqG3juna9I0Sh6M4Uhscs4hU8CYdwIouHC1ZPLcM+MdW3bymQ
se2IFgvf+lqXqSrlYGy9Am3HMo481RtorrX4P+qeOhbYU7mNgsD7RUaV0ZiU42TE
dJinXZ+wIeHaAUsRH71g6zmeBleXRGtRPgygW7BF12NOMGGFDczV4p2wlqLcXTf4
cfGAfWwwIfNDD4F64j8UwJ6YRUUohdqIdw+X38/6kkvWPNS5cQOLLq+WYszCSazJ
wkZnuWuoAH5vU3GUU2Q7NLWuFSUqC6SW959frL/cmXbEg4OJ1vFcB76yH1fJxgJZ
P3dWHhw+J0KNRk/EbxfFn3IHtVn4SYLOvPLOu/Mjws9L0ys9cgmwJHelEhlpoBxd
LljXen2pjkMXWiwIl5XzZpi7oADqzPQkc4Mgo6GqrIPyYFzsKGXTxPRLrcUhbrx+
21nztkPSPAQ/OhUhU6AJ1eELsjWvW3CQeV2/PrgsZ6kRVOI27CRD9RyKckCVCDBJ
7IH9+Ro1WYD2FiSGS/GmUsVSqXxT8jG7EqaakRDy8syorl185ApDMA0BVqPcZyHX
UNSQq+doFqvWoTROTzj9By63dOeQiP1N+/YRArUIk7lmXRH9b0hnf5xIa53eSyQ6
ZNEYqHbpQq7gGKDWWr6MvzbF1S9Vho+sENuy8wV4ghKj/obcdsxVuD3zSzllWwmO
yEY+vILs3jjH0JTt+5RE9KRCn+Lsxef6+qhc8z1wAfbtn0GaPZHmhEayPDDW0Et/
dOX74oCAc9A/I+lxT4ct9jXemS8Nq55PVm9kS+RIsunyh/TcKelPd/c9g03Bf9HJ
Vl1dApw7WC5Y6TveeK+gmZqfN6+SAf3OwNXDM7O0j4ZVdQgbKKF8qTrWYjjrY7G9
0Mbn9y6WjbGiqAzNueC2FgshU29LCsoJpDSUrmPp0vDstJmdY6He1FuOWJlv69LY
BWIb1IaNYWZNF7SvrZ9fH6Ii2GYYP0WZMKjPKXiS+YmCANx+2Hh9C26me02pAN2j
3WlDTHKfbbRAgqYYCuZ67kivLJsDQU3/3yNh2u7hIkIzc3GSW5hgtsfkonhqpwgR
YmHc3qEfAn56Us5eQ3XOoNaYB6Yc+WBNJxjuVvVf1SrWe7UCiDK3iboRPgHzvSig
EwWqvdgIUb+gUdtOp+mb1F3Hyi5jaR30jaQaFMfVcrRZd1zho4owdNfjSzpMBiKJ
/IGVKkynKoMlUqg2BNwf92MnqetqVrwYcO+d0lhu76PnYNCGb/Y672ZTce12ruDf
2ehM7ChKbHDTu8paIphdbSENOT8xUlJu2jmEjZPE7tLk5g3FVzRUBvJooEOOSV3e
ltQNWmLmHVCaOY+q6Waj1e24U30lIDxPfkdg86AJ6wDw4S6Ck92jUi5QcXgyhsUo
5jBpke2Q/NjKzDqKI0Q6MX7QnjuqHNSbhpWEYpXWcylzvHUk9psjwI+Du0ManE3Q
t/nCbF9PnJBY548OAHU3Wu1m1K7cTD75FE+6G4O6u1WEVz0Biz/CYs4+3aeJ//DQ
zZ9wt0Squ/Gig2nNrkGRKFWd7NVAYhr4UPuKCMAaBzEk5uANcTwh/mO4zXC52m7p
W+0GPLURke9ypptgE6DR9pRqrXrhG+hyzinAqEXOwEd3DPVffNLD0woV/onBjrdk
DPAeqnzxllrP6IFsijtqzRY4deOvrmeWqusDkBPUTwUJHTxD41m6ZCy9B7eVidwJ
bE3Pq7/7i3u1sFFIgP4U1Szd/EcwhtJoVsb/XM/fBvMDq/VFWq2QTVoTnZn1GnQJ
nBUa783XxuJmrjWhHSiAKsBEA/I47jTyVkyOvE1B+mb5bzhKMVY4HZlxoA7hnWU/
F4LxAUZog4yW5ZxWxcEc7El8QQnZwC69SvYiSWDbIwDX8HRpfSq5+miPhmCPPTe6
3QT25hEBuTDiMgoW+l8Fm0G6VcvTmbxQewCNjS66JWocpZZ7rlqtxp4W62K3xYyH
h/LtBSahiAdcauqDcENQAy/6uokoiO1jmTV2MgsZX8LfIszmY8VgVrfsIzLtkX2Q
pSPgSDYZncunerdhPCdiE8YPEEvyYFD3qXkDzmwXvZ7TJwYpWGS01HjmP7EQcXGc
gnFk8cj+C+K0l3WuJKfA1+EcoVHZQXtmWoUp6hqdg7Zt5pTQrqAtGa+PU2NNWPa/
V9CWc8qqvuBkYS6333V9KD8nWyoscd8f93/XvRZumii8TRI4YdWJKU67qI7luyh7
5D1zAPoNspNGv8dLJXFm3fvhojTU3ujelBisIGhK2t/VKyG7sRsmxwB0WfmGX02M
x1ki3hKJPmlKyJiKZs3NstVkzgmeIJjqUhEkwM0GFV5lBErcuJdIgNb472w123II
onYnlu/rXOquUrjlk6Z5RGMDE0XDbqjbU7XXxT6h6BYfhq1axk4uX5F2UT+z7DEV
Pwu1Su94C2Venc6tS+ngKAzt85l2lHRdL0fkqCww9iGSydJ9mObJauRbgx8+tHYQ
M0tL2dxKZ18P/fhdN4V0Ikuhd/i3jdACOpVV+p9hH9QE9kXkNZH3rIkIpQLRMd5w
tA4vp85NyZ7bN/u9rgbAqz+8jmHHI52D8mWM/1QiO8vSCchd1RVccqRpgFn8RRrl
MGxVHDX1wUDJn6XNn/+QaHPoHOYS0AkZsQVkIZiUG8HbwgwZyV2Rrz4nv6TQUZ6j
/NTijWTs2lqY/qzgpHvSqjmY6YDEAah02PAQ+DDUOWYQCCFvlapN8HkTcUxr4jtr
7rYPxHUx5p2Nvqt26G/e+Qntp6pwb4ovDLuOfAdN4jQuFA6srXwycBo9xE3n7ey0
1zZZar6OnMd0fThA3SuTtEgxzP+U85xyA0eF8nMcQIg7YFRskvreiHPEGR/fgaQN
0spzGD5kRP6J/Rr5zNg41ueOektetKeuNsXxNx0/zUTG9fkbY5EBw8hBkHnHcCKQ
agJD9434mmf3tPTNzGQkxZB1blbLsz5IA+Ib/cEgg9A44FUogLT5ukPvMGJlGie7
mLOK6dKYTf16magyfyf46blPxLGGxBFHwerRG49eGscxYAdoeCgcOoBBE3uAxENi
W+eIq6AynEKxg0Y0Zhyl36lGGs1a2FF/wfpCqjZ9YQsDg6qiBgsZwL9rH/0mM/fg
SOdsNMaAhj+eg7wpNottNmcAUZkFKxPzi6nRG5JYV+P6Q6HJWqARAseryeqUNiDv
2SwPHUoJwCO2FqMA0ZyFYc/5FpoMrkAtL+L+omLe/DFTfEL9PRFkoxJkORw18Elc
Hez6HZFCt5S+oT4XB5JtnGU2jbfZFFw5h5XEBNjZ5cxbrzgPTdtkllnsvvtxMkgi
VY+Xk5f5/pkRNgN4dd3IpOmzes1OfcL4CEu73s1KGraSTCAXc+x3Mvi1mx7+y1+6
zel4cLr760NkU+BiY+NWS//bArACqcFxD/3unZeCTTjkgceU2Bs7fFolyisfnCKB
Bm5PkwvXhRir2+cgzmOIHo3iKN5rQefip9g+XhITfSgnZKyAzeLoTwCDGRxDsGSS
/nZTGVayuXH7yFIu4SCzv/JITL2z2HnrOk/hnIwWQd9GPn6cfNztgwqbGAWvO694
TEP3c/tRom1Gp8piAh4DKfTAOvOzNEaVWBSOQNBG1k5J/CIF8J0Lq8pru0xEKh22
GjSzfzefzj/fAXnxHqWa5niEu/vM4W/hdhvRpc02iaKipRunAjFFPQgTYWXCVkgo
0g5q/iLgqB2tJv/l/3sKwaBSSOVVL04U9M2l+GB/ODro148hwD+TCD4cxD9xdMZp
qkNZnMElBq2k+goR5yrC4dKgcFP1yQbUnvjMT3fYXWR+Dip+d0vIeYlG2OBVOAvF
jSEZ1XlyisspQJZgdM6FjQvLgUXan/PQRWcUPA+A1Fk3xIEdcDAhRLrC48nkxBY3
ZlTSLgBIE6JJ8HS1r5zs1VfdNBbQ34aZ1i26e9/EEQajkyKOVIy8Wm44v6fB6fXF
REr5GIUiIZvvzBhRB0znzxNJQp9O/ZfcWvQU8UGqLtZAgU3BGAUDpBv6Ggbkwa5h
et7I4fZo03L7RvzK2cWY6lbPXM1wx0eu+mQ9a2R6Qmx6C/zTSJ/wEt2qhAQ8nIDH
UIgruWEtooeidz2NTKzsVs+0y2hzAM1sM60KwLQJpDnzwXPoWEk4fL9cXB6WDOFZ
FVkgKBTilydLSgbrkbpkm7L5Z1Xyv6TZp8220JI0viF3VULXd7VkyE6eCCCUMLdB
dpsOpXz04xvSEqTxi+lrDqMHhiNsK9zm9BrocOZIsMqi8ytI+tpBoeAe5IV9+Kct
C8gWVk7j4DkR0gCWfIlPmTtc7RLe6JRZslbNvwTm+pb2QbL9Jf9l5sX+evqCNL2f
6IJ0+1LfPsWutW93bf1nFZahPo2sQtl4oM372W/1hSKnsK28AXXpgorCImiXTGRR
B+tssdoayi+Xvd9qhHx9IhnImLcUsT9cJfFprV040vaPpXAwUGC1rxoR+SLkfehq
WmXF79b6YxPtxRjxDl0oDTm4G9FTu9nzX2EUrtSX4N6ca1U3P1s0wefk2va2PX/Y
KDhLp+u8tSeN8wV+8/4NdKpssP70tmHKStoNawkzVxoUnV4U9R9p3fgVS4ssn+KX
U+9xaK8PgzA3h9VBphdFnJopyzf9CxD4DGwu5rtXauuvSuwnmNX7XSkxntsJO37F
iORH7Ph+jozgKdW4ohIy47XgZt4D/sOgMXfCWQrBxuBu5hoHFqF80CtfryXGVLyg
owFK4xd4nxcxXHq+hUbOKMYNdkDu12BeMOmn+pwHz/RcT5M6W1sqH6xAF5oIE8+v
sKOwj9X8H6G+ehC4RtpSKuV94vRGYqnjs+MUvDVXR3bcTBohV0ZRCCYy2QCjFqXU
mYyA6sJ0O74kmWXohFi3a4i3s7/2xJf6IFpAe5uV0Ufaf+MyDbdYPo2Y27VC1Zlh
vJP5xuDPKn5wT4g23zGi3Xb/cLdnb5JdWgsGdiQOFhbenJfsf54x2oywGosQLG+m
Bu0yhUmaZI8+oe09FLB+kUAsZqKHt7tj9SyB7ORPwLNR6XBZwiQpJC+VxJtDtYa1
WgQn5Yye/NSj/wzEkn/zFu+689+2dR9L2Adn1Uwt2+UFDnU2bak7LkeXERf9cky+
4Jq1OGnIHJYqo33psmP26417Qc2jAAu8IErjlJU3XlVDci9yCv6Suiaiff2cT2dk
bw93MfW2bQrBHgAmztb/I3PEDvWLC4UNS+Fdoskaupg+rJgXkL3ElxoNwC0O41x/
NP6QDPiPzqzQTjCmfUq5c+boxAgYOhtag14tXaB1u0PgPg54GILdQEQOJd5T9C4w
hjUnAAeIbZZm3SSfqOpQ+ddoAhXGQgJgdy6L6xyEvcvDJs+B/YBbVt9YRN/HFibY
/lsR8gGR11hksNjQY7GZ1bA9YQfZNG3htMgT22afZYgsvr69vmhC5gUi+5IsKe4F
uWERqwfY8mkLtxbM3KhNCR0/1X1fQgOgFiHUyTdraEUyR/LLlpDObwP831WFFaOr
wqdzDknecP0xQR8RAH/GJPfQMVo37N9PeQXJ8bKk107lfCxTvcxhjTr1xzL21zlF
jycfjyHkeRu2MooghR1Bg46oEEgf4opF17fn5tjEUXErY7MyMPCGDcsBXe8H2zL9
joD0JCPIDl6JwYF23A94m/PlAvbYcLndN8Mz2gcdPUMCBJo1sl2UW9lumbiBh4cS
j8Qs6eT7HsmTJFmyjbBeghW2fo1JnRJ1pGS39IbMg27XufpqucD5e/YRYtRB2C1B
iG0FoquDmmIOXcJ3iHem+9TuNjHi29b1xOkNaiiNdt607m17zQrJEFeluMWG24p3
woppqllPGBSw7zuTZD5QEMK8w8xGQMcrzA67E6yCtfZHsvGDWDs+oKnKKEOq5haq
NfTQXOLX2IfmAbnWDOoHAkXXBGTHj6yN3z4N9aza6EsakgwhZUs8oUfBTg0JyZfk
wHX6qJNJ98McgAS0H51+eR1TmyIImORHvN6odD531Iwz/ix52fAudCN+q6LcxB1k
TWYmITVlUkD+Pmq3MfnfEHX3Yki8YHCSjkGAO0f/ps+OKt5kYHgpE4Z3pDbkwlnW
aovmbu11K6DdW4LoaYBvYFC+0F0rHzme2KoXlbZf3Vvs/5oG+p5A4w1NNH5/l5h7
TbKccVoXSovgN4ZzWut/RzM+7xoGVu2rq6Q4U0l8mCwVJM1R7x4XINA0FBXaZLgm
w6PVGoEbWb0dsQdTfqueycDyUeXFCNRIGP2ISIs6w5fB7Q91B/m8/26GTI+/D+uK
5NhVMn0EYGcvTsv68wRgkAe9GDLqQepXR7bEzXm1N7Bf29R4c1cnXcV69t/0RYfH
kHaNeA5e6kX9J9rvM37DYy3MAsUxg0YM0FxKI3CuLksSDbRbvEXvJ0Akamp14fLs
e3bKqegdDWkVFnHpwme3jDGyd7E840O0PFa7p6isCn0aywYeeNvI0id/YR1Ot2VH
k9MA+12zaGN9QQoLCiaLcKhH/4bXFHrakVqZeePXWY+TBFRHSoLVagEFn0DPf1KA
A18MXz3Rt4fZfllF64SKe4ffnBokARK8OCa+GS5mXg/sEAjly3XtRRNlljaDPU1Y
n+ioFP974P+yB9YYzVTH3UFxkglCOmjydPReWa9sIt7JYayUcGXhyAGciOE9BorK
IMCQcjwg7fGIvXmZaVbfpZsf0pVqZMV8/Iqo+OC8NKD4OxVTQnt/vn1AdTNjgY/x
rJDo3i8WVa5Xufea4ntcgCVSNoy0yL+bQqPXXu5E9pK5PJVlg7q2dIeEH5A/XpIL
RHlzM6oDbf96lYAcIhK/ONRWkhCxbhEhXe0THDmRobrLqDjKw879bU+LdzIStSjc
J62LQuooka43Sglj7QIua6LAFn4dlPAK13CSGF6ehp0EubI7nB+kC5EeWQisBQMJ
/dmRIX9tx+A3JQb3GyoYLJu8pfo7NoaCrERHLeHvmLZwjdE44CH+ZB+qdHfya7UW
gGxH8TnIOziiMwV6Op/DrM6to+vlDmeaYmUgG/Nkcj10gNlXiWKbv2yU7jJrX7+F
fjiPh8I+zPtCe98AfYCqguM38UlNDDcyZbATup9uUULSRc37orEzP6Nrcw0hYI44
iHpH7B0vwA9TwHc/K8cl1w3fI+xriyuD9fByJ9MOkH8nDZSkn8QsTqQAo0Oev3qc
TsVo3TiELIgJ5Gkl6gTGRTYkn8I6fNk6hwAmxE05E0l7YG7S0YLQAs94E1s2eu1k
ggFM8EYt6/VYcdw0JqpC6RMPaFD+KH4nvAHe3tiKg2LM3fRZEmosI+MNoAh8Xj9x
7tfJMBBIVmmGBXog4anALb8kwiUDk4J/hl1FgolXUgXxqnwG6eBMnSZYXQ2/PbMm
pL+C4edNy+V1lJXUdNZLRsueakUib+tmKs5kP5zQf+p14d53eRqOR50PaqtUKpCq
ozt8mVpSOw5mYLjJYfLJYmJZlS1D6aqX9AOJ7csI8GsNOY4FFVTZSDN8sBnc9Wur
+CJe9SH1HHZUWR8Mw6DHqZ5QGD2AtL6a/jJkXuhYW1zEUNb03Y/xURw/vV3mf1ss
1KhcRaJgt+E9F0uw8i1woIqB4ujULbw6uUiv5WvrxBtN3K0dCJzk8TvXeDrF1Znp
o5FsH6O6gKXUH632BT70umJlrhdkcLXXu5inEB9c0I91O5o1hFRN1dB7/vhasj+9
LqjLHYg1fL49vVZNLNLpIjnMt+M26jrjN0JwrBFZLkuF3Dh6FxS819Ai+i4WaiMs
1cw+xBu2EegWrsmCgbJGW9n1Zd6y7fhbFNZ+qP7WaCs773rKDLH7gvHl9cnHHc8+
toU4t7Ina84WZUidLJIEdRTWEpGTXxLWlkr1Fu75kMUVa4tK1cj2Crfz6QPF32Pz
0CFFkwf8hGSlrEJbF47/U1hwj8Dz6TIbe7zpfcJVjCyhR1cGyADzM6z/NTCljKMO
29um2V0mXm357smUJA9h4bu25rfY1OgNQBQvAnzyOGSPbn1G9TNktWycWIOmRJv2
DP+oN53OrXILMCwEdC6DYzZZ0RoAePTJfkAEhlndW+DABEgQU4fUQL2W2b9rag9t
JO7eHvUvNHvkhtULWHw0R6GNHzFl85FDmdq3V6uLO3zUIPgd10fx/ezvMZeYLSfF
8wkirpKt5MZqRFOHE4d8cyc5Im8h5aqK7lG6RBgQIGh5ETb+nLD0Dc4I05rcVvE8
r1/S8DAkT5KtvqIyrfmyLdIW6J8RU8sixQV9779gq1NdsNWH9QaWD0lKMF7dGxHe
XWk8StB0k4TggQ1q8ihhodd67AR7euCFXF2yeq0iFjUpCAbtl7fc+ChtFfFzAekM
bUtPEGdpgk3lReAPCGNsyFJnw1rRUrbXnj6hyUmEgZDeljEru2bhYb2N2vQXvgJX
zQOMJjx4a152Oti7GzvtWX4KVlAMmxzfKEjzEeXWLKditN3qZTI368TMhxF6Cawd
V5bseUs9pXCJbrQxyqrvl4KiwYqhb+FLTTjXVqkpg07ZtpysYP68uPAfUXoFQzMu
8H0VHScQg+nexOvhqZzhcggWSxwtlawNxoWYTHdy9fny2Q2dXeiQipSc28IHBlP2
DHOymQEmwIt4jalAmXa/P/1XE9ifOZyvo6S6dTZBHaQylZziGm10Y76GVz5y3Uf+
2u7Os3e4wy5+cmPtB5cn7W/mPba6lrgbEYP1c/pAnvPvOTT4FC1sz48P9aaCjJet
RyJVATaJalKFeWOVr1xIt5TQRV6F+cYFTeKS0YTygUGs9VrHYZdTRvhRqsefGFDd
yo1eGLnCxvrWzIBbisQRZanJECAj7F/yU+5gEMJTnbekGxwcwSKDtaV8xbLc5L4K
RN1CNYDYjxYwCdG7Ue+18kaSGz4wnHx2KxR420rHpbLI5lVjydHW0l677OenOPi6
nvi+tQ8qWCmTTxUteHE120WDYNrgbBkLk8ZCAUwPLEjh1ue53SeKj8CyzRlvBGZ6
PNzByBaW3dgGMdpR2fPZdrfqVv5eG5pYY5F9lh356sBP4n28tAdS9912YXu0DzKV
UqkwIbcHvFl2+Orth4I4pUDS0/hjK/8lt9Cl1AjvDnGc0axHuYFEwRT4vhTrBFTG
l5CA5J9Myi3rEpE5kIg5vLnqewnlewM1rl46AJcO+UrjeZGiiuGC46BsKhGZeV1b
+WrsBjTEsmFwgNnmRgO7NoJQuM82FYu17XS9gFt54IgkIfuDmEEXrC6kt2RNdly0
PkQ3nLtkrKpuvaXs1nnvd80dPnLCb/iLj57J7bZsByk4G5Z34JfyHnuyGFbZuyKe
0JbAkM+FJ92SX6Dzi2PKLd17/780yC5Os8BtTy5pNFN+Ma+Dl9U4r2FBXLrFXxj9
lXjnpWuXVV9u89ZTTKUI48wa6+TCyytcTWwG98yLQrp6KXgDhxp8OT7Hx8a7iobw
fFxqMKtA6x5c9KSnndLSiGPu5uULNrkZ3kt4uq14L8f2RUZh4vNx0RjtSlnVelNy
7wen7V48zTVijV29xKlt/lFxLr3rqFYmNAEAo1IlWBXrXj+9ZhwpVzeaS2JiliDv
4oWpKUxNkR8kH9npZxLaeJ6aQbSEy9W4L+SP18FbqG3w73PCo9wgQcHtLg5Mjj2V
MGLZGvt9tXGYPwMIpgYYIeIr/goudr76I/pgw5Nimgs69EWnwj4HGS44VaGDA6zY
7PtlDsjZhXAwlgL6o9QqAkg7Q5I+wtrrTQ4YOCaQrFe3VUbv0vqfZZR5hrnVaEvL
rfdDIZ9X4ihvW9gCwKIaxV70pQF3szORqyf1uD2oK8DGDy4NN/i12HMSAtoJ4jy7
8pRH/g5/iVxeiyLIP/5swDvD/ow/bOEptd26paUWdY+RyrKmTdfICX1/HtnyvwYQ
MagE6XTgl9wiJMrcrKHjMRCMP/Rh5edgqT0+IXcx5ZsyE25OXTRve+eAcRhcEjqE
OKp+AFgh6mrFdyQ4yWgQNU6L/2LUlggrsm2A9g/4z1s2e+MJ+ooBI6Lkh50wX+2Z
NYAegCeABu1f6CKmwm2aRpCxSLqi4iaNpN8ywqNexyBm/EvvJKRzKEnQm3KPNxLQ
iH9CTpv9DpgsBXVAUkrNCM/tsBkh+omSdmZ5UMP6EY5C6DaietCCV6+b1F3h9PuK
/dNRrRu6AI/VMz81T+RirCoEeAzlevvEludkbYwfFa1qm7QU0D60V0R/IiPA9JE2
BwVJlgv1Pt0eOPFwUgouo/MIs+UkoqPkBPMOUkoSpEVFMdasIR6F4r8v15iw2EYX
/mS1xEVKl42o1V4ue8MTolhpxZJ1hv9dlYG6UUDrift144DQe01Kuvur/7hEqXsy
7b3LYounv85LX2eAjxzNj07Wb78CYhEVL5T4loViOraf0M7X+t6PvfILP039ug+7
ir6HFKJEHQr11iAP97NQEhz5MW8c+EP6H1D6WiM2ID/6B8gMD+zpfgdtRyv7mo/Y
3ZUsVxO6hmgnrJ4g7ksy6IcolRcPhBmffFKGRM3MX8siIU8xRJznDVWt6ohuQpzq
NtNL3DmmDFaLBcjCN6CEdQVY7OudySJLlzhctbzYakjBxleDIiNRVA8QLem/ZzRj
ElRb1xZxebpEIy0RU+VKfWc/DcwihrBwSf/mXiL7Ow1TQeNQK5ga1YB15Q1Iz9MI
xfOHiM0DhAMEyO//4DpNfvSAMcojtDUtoHnFLKBJveTNTICWe6zNfor+JAdrwZYi
wAdWZrrCrmyiMoC38nqcU3AvlYyaHtLl2ZdhwtpOrAMDc+8l9gJZqsKSRsMUUnz4
bHJW1xkfVyN6olMRLvmTe1owMXUBVONVyuq86SWDPV3sjRCHKC24UHiY7OvgqXHU
4QvzrKPx12bpsgkc/oXaGs1irBGdekc4dC+w20F7rAPhX/g1gStET8idvdthAfi5
3HRQFKKdZGytP1Hp+VYkIYjil8jehRanH3jRCBzc3MmV33JA/A1MVN23Aq6HcLLD
yTkBPK6fqE/0BOJ64r97Nr4cy+qVz5Ym9aSEFAEkfrzVuxd9Z2nyUkrskUnX0p/H
iWiKa6fLT8FOcl6D0fLULtD+6tgDRUZZj1p2BYfd9NZsQ2IYpLP6OD3M0h8E/xEQ
uZzE452HCBuj+o4VxzTZXvkE/26YUKpDrvqHzPG28SbdUxgUp1FLpANVIDTxFuvV
2EFWwV8NLt2zXtPSn8vMBMiYptvvcRkiP0PTTMXmRBl24c+pzyObJlFbDwMEhReQ
Ap3vS2E/rsYu/zdEkE7yfvpJJ5TCuYenZ6CBilHr5i6Vp+GAVX4+vFZI8nhuuOms
KJ3rJASAKdd1KUZiWwVTwAwrH5UYQB7Itur93KQxhqXvESrOQzF818E/H/DY5jL+
ohC6+pIDezsIw2lJCyv0RdT99gUAlHBtRqfFzfkmQtTMd2YTx9D6reNAwkMCP5EO
F8mtFrco4M0vuSWN6gB2DD2vSZxNCu01cX+6MuIhWQ1WqT5S/mtQSaK5mYuSkh7H
1o4661gm8w3F55UTyDEVCM1OtrZEa0k+8wkeXczm5JHNDmgS7RwrDs7o8l2qSeHj
wGXFc3KDAh1H6m/Sm1nV7CfUrdH5q+ZFeuL8kmHQgPH3VVQOBoRivRJyOSRwJA87
diliogH+GQnliiOaR7MwZc2IanNoOkM34QEWrxUd7yrUJE3Tk8UUjyfa/GI84mL7
Nrhyfnkp2DxkUgkiOEH3DLqPxRlb6AE1dQtleKJSCUMU0Q5f83neQ0JUV0H1PS+s
FWJnnGbx5ztpZbp3eiGGb7x2TV5QuWE5brJx04c2ttaATzLOzNQpjcBirn3RD/LR
G2ZQvTCYt0BITSZHtIfociP+ONh5/KiYh/YTK2TccWpsf2z1C8KBoPrJKCzg/z9o
Y6lGU/WidNiWoJhZzX5GJMdE9RW47S3vETLC8um0kKAlNmm7VOsNkC+G8lcMHBMV
pKOp2bJpRZa6n5jZOsj+T+Yd7ovhGU/LiWs+4hrjJF2F1CDsMCSSTonWwoNB3enC
ZleSh99AWbf5L4xF0sVFtWNaROX8JZUwJklSTuMC9xJU7P8bmbA5WCFls8b2Qi+9
E0eI819/1Yym7WK/C5wgZowrPqbi5p9nTH/mR1QPt32g5v1n36MYFwReToQdfC7l
3CsFU8HJhbU4QKp6Dj/5oWMr5Npj3E6xRq+z9NqykhkU1A2PtV0h27/Eas3PwKl6
EPMsBww6KYMon+ikR3qXfd9I2RCdh4rZWc2YenYyly0thOBvh+Rp/qNxlnCcchRQ
lFzRmu5NUyFBTt/+10P8uROEa+5z/DP1ICGKsX9hh8b+bpdGsJkyYhUH4E0ufr5n
TBIkamj5sGLWSU3WXyUHEW1ZjYEd2oG3mz/P+HIHppQzh5sAZjIf0bhtgS//Rw8C
Q0xYoTjO3v55N1AHMBkP610jbe1UaoRjT7W7EgM9ANYikWNu6m02clp5wnv+o9oG
mdPI74Epxyx3JZ7C7JDI2AOyK6xs71hpJIIGWeyE0GwPogeIqBa9mJafXDwgvEsO
ODa+cArtaYX1qN4gVJ1oQs7Tkr19lT1qWMY/emFCR1hWz1BrfrYaAg9qUsuwQFwf
/p9zHtyQyUUNOSXR+KHcVyk1SHG8MH/XeiGW7qbUG+KOR77lC9TFvQcbR5HzNvWa
FYn52YXCffztZuQn2m8aRDmBa4vayXNUDyrgclWJx6GdeD2Mg0GCza4WD3izZtuK
07ppPZ8EdMUwN9jTllbXySbyNUYJ0tCMvD8hutBcivw/XXSu20UFl5kCGXpvEKeW
sjKDs3nZnomVmoLnzNCVTx+7CkS7sMMenbOI0Ll6WcmFeMzeyc9/PQgT9NT8zEGZ
YoRHNs8oV5egJKBmCij/4UWM5aYBRTm3VSkWJmIfZcss7xNpYYgxK4tbFZ3++doT
2JhfHYtSxG7aEGkFW8D9Ajb74KXw+Q+PvGirrXNDiJ3UhBeXzcQeP8vWqcmxulO6
UnrPB2/m0ebPjL8qQKGbrSPTzZzWUITNX72nPzzPf0//b4qXPiSu5vD73YAa/coX
W0sIkArrLULCioEq+Q1NNPDDexluzaAWSNsw9zsgftseV3osrENCv2DzpAyknrRL
kSkSOz0yaGqHfM3NsqlyukDxDjiZwBiU+QKEYCSh29hGAH/gWE440ZOGfQzKVT23
Py/H/DxwoFikD+DaQ0aUmq0+mP8XuC39zNXYheZZJoVUVp9KF61wY7ky+9FrpZY/
wflh2IeVepVIHNq7uEX29GOe5sT1Dt4XD/NyC62Q9OW4acqYtom/R+DxCXK8auvK
0nCo87IxE1LG446R1OHAT+MWlAF/g0ItnF3SN4BUN7b+wtobQP/tF5CP2Ml94SeE
/GcQ2B1+/QDRkmKXivs2hnvrd8Lm0xcEiQA8Fmdo9U1a2D6RDp1ifuDwuRttQbmz
+Obs7+Mb0g32yvO57syBKL+HqhrOAh0uTA+D0DvlQOxjnyG5Y1C91BSAlHdtObhB
ya4wB0kwXrupfcOkGNByMvvoUUC+NUJziaykbD69BhGLHc4o7CTwqEFsZoqN8o7U
goKyivFCq7JJ7Ctp0b5JOhJJOSMQ1diycLKxwVc5u0Jz3VfunaV92j475tUbtr6i
cw4YM/9k+8dhaTiyXOcrxo7i2oB/5E5JRmeUVi2s1ksKsfJw+zb+A1BidPtA6Bf3
u/tqTURws/knrZK9Uf0BpKOZMY0/dows3737bq5wY/N6McMaRPRIt4rKZtcsVGCI
5dPt4Xdt3b3c0/i9mwzR4i6AMhx1EUi6JiX+kCI1SZSqCuBgxDwvd3jzxYHSL0Wd
Gherx8d9iawOo2cLCBles0mxB8nrny93vn2FN+YSprVCCLAfLobUXrtXliZWk8Wc
DV3Rcnudvi8XtqDNOA+d7nBmZbjV+kd/z7c6tnv5RHvTPsTdGPV7v974RfqadFpJ
E2PhzxvDlQ8CUv5TBv0UUcl/lL2hWna7R7d/MWAyrdbo1g9tRBolTjyN5xOh5h+p
LJ/M9HyngchIcog3IjY/WZ7cl+CnZcXONEaU8j+np6kDEslni6etZGBrG9fo0Jl2
0GPIWxqDHUl+QnG+YcDoMAOJcu3YMEYzwZi5PUlHBcUXBC/5GTs7IxEGVtbi6IR7
7NP5sQlw5k2EjG/yfSKnRtPUG6lnh4nxPnusvXTYfpmChI9soxU6XoclApXFDHpQ
QoeXPWqNViW9DIBrSd5cqojKZdgeXYdof/bV0SIaaPkH/DR+ZmuBko5bpXkPjcRN
FFNzxoHYJS6da9mqM9a0NZPNc1SExTxCWy4nqvr0sS8fg9goMBI57mrlQAJjliBd
jihPlrbjQxnczUEzInrzzoXrYzIL6Opv7xqCRbYxEPUOz12lGs4or0Wk7aaWav4W
ibgBJs4KrniLm79q8ebKApRDj91QzmmfRDF7qM9E9V5QxCRapKufCLQluMXMPXau
8rMR7rP1A+AEA0LpVkNm1sqZRnQow7Y9HUU7ME7J3E8YyaDcmC13IOU7eE/sx/BQ
fsKkH+hEMBz8yRhr9EEV70r24SyYupJtXprqXJCQ5imNf2yvTdkRb3Ul5F6vZXEL
TCndJtowHieYkJjPSYW+4xlcuiafqe404l7mzMBhLNmX6T95agp1r+iSw11MGRo/
y+IHrNkVTybt+aj4BpbWX6nnmLgNVUg+/Yi4CfmednqE4JVfqmUHzX8CKGt5AJz4
oxEsWn52VDjHWW7OGMDyfvoAnFR/rw/o+t7AKrfWKgfhcSBLJW0k6ec7Vil5+RuH
b4vJJr3bJ2HY+/r2riBH5d5UoXii9eXc5EYuJJeH2XYzp3jO98NwRjC849bdbtE5
ryasQbH7/a8u1bbmEXB+iXeI9lbDlGTrxE3W7vHP5NMWDiiXDtzj/tGhak3Bq/yj
5Yp7eLW+IXse+QfEgWO8R+xzVI0BG0byVPEJ6hIbXIXEYnd2C3jKY3EHptvOvdbT
afoTpNkpFiqGrxCqqFBcosC+EuF0U8wpwjZPQ16FRYJQCh+gkf3vlmfQmCh22jrz
EzzMsdwVkdjlUU4z7ln25zeDci8J+9/wxr00WgUOo6cC6Wdao+OQ5ET9gLQjSnlE
YVYauSEgjHTcI3BeIkcxJ1Zvg1Fi0z6bJJMG5smd6SVOiJ3pfl8YRFrTMI2VnFcc
XqnZbtExdYz3Klfge3NDkvHOBPpXj51ZFiJB2eIaSsY1sheECwvrIiyx6TIKzyUG
8QqJPQlmIOUSAvKvOYCHpNhjI9cRQyeCGwfs5SP1sL0TpqVwgyoFCFbXEbkhcrfO
36loxF1nB5BkpkKM42Bp5aNLOa38A6OU1GhQ4gSjgXePJUhLKgSnQgBfOPmE/dTH
FW8K0NiWdeESTDHDO0P/X/XfX6ZwOPWO6VKpXASL0RT/5vbDtTgn0Ptxgmj782rC
vLR1ysgvrdthQeL3UjvNqtORSaFHqxlWH1EaL12ltplAEnZfI5fsWwSXiBmKthJF
5XE6vmIf2Sd/BNiAZkTmt0YeS5srkBt1jmG4oj9NYz59CqykC2KYHyWwILMPNz0+
QD8doBLiGy+rKi/or5n0sxO1bHMGgUtIgJlEbszXct4480o32tMwKJ6su0aA/rmE
/048fKxQ7KAwZK38O/IYcqVkC3jp87xZCQZUzDdkZXqRmxhQjcqoOqPhOxsN0ln6
fTD34weWIMDvRxwkyuSbVas1w3wkNPjU+D5DnRgXR35Xt9I8Co+mZ+vjgKDL4ELU
yBs7MsCQxlK6cMzerAhsUvdclapKFJ7mFOHxBrFwbKAH5Q/F65NjO8dN237BmW8+
cLOp+RUB3N2jmt/7aPpCWvNOGvUqOL8sJ9c0+uCZZKyKSngxxjXPPBITRIzG1JuH
lapwtHQvCWd///hVEvxUtWR5X7v2WL4+shg/pl8VblMXdlUqBnGqHttNGx7SCv34
smR3ravpDmfdGinRlx046ujswJ88UTsBlAKEfXd7eSKDTjw9LbFANhA5zpODpxRn
4OEpOUyuuowISZrms3oCB1QrRMVJjUnyFjlgIiJoBcoARomOM6oYIXMgo6XfOaYL
OfUgLIm7HdLcP9cydItGY7a2l0s8GvhbcP5ECr0Ki3ZTlK9rc2WhGfaGe0+eVmps
f5hfnIK//DenkrA1Hse0KCSlcxvctompC1k9+h1AGcOYJPX8wRZ3WRmsfudz4+h/
3A8xmuo2h4rI4Z+IjNU23gWNixFWoMhkId7PMyxoGxE0U3ZfcseUIbzx/skUxU4V
P/j/1ALG4cr5KeMZnp0HrDuLrdTimD2MSPcx7dtiV18O2+ohcY6qALBt6zZkRkX0
HEuVZXF7YuttSAmfcubY7CjmEwoxXiElThlYYl0YWPLWhp7V0ivHJXJyTD2+4dZO
n+an7QwcXQM1kbAEgiCwPPxkRBIYoVXYHaEYrHg3Bq1/RGVzRtGU4HO3AHdpdDxK
9FDIIkxHjQBb7CoW2H2QvpFl2r2IVFs+g3qGbE36Dmo2V6is8KFLJPXkejxyY4jm
F2wYKRAgx77LTF64hUbLH+osFTo2l5Ur92NaB7+e5Y0ku8ABDqh+HEEUXxTI+Yt4
i2zdkVFNiohX2umPvx7c0fSn+wO6ZK9GYbANigp5U6DtXMX+XijNgwkMVD4jPDRj
li6XPFg4gnLJuxJESBFWatuMnJkZvGWMsDnkcrtCuFAlY4dlgS6qk7YtgbfDT2o4
CLxWWVfdn99eZ+cIDwZjARB+DB/nqJEbGtRgeQHx60OFwVatMgPCbmpRIRv8ys/Q
GuofeJG0dnQ4qBy4wSxyWaRJMqnM0M/VexPB6nG4KK0IIb4BDmuvvo1y4f0ymZpE
o0dJMX4vOLsqDOKAKZpT77zCECtpeJiSv/eeAwNnsVXKIpWX+Z8e5yVig2N4A1QI
vu2QBy6wOe3Il60r5aE7dRoAdvSFJxV+D/0bg0aSObisoWEEwUv1EYorGdJLW7wd
oV5Y8w4A+GvVb3wtOFWxToq+KnVHllrFQSxTXWzsHf2k2y+CbwCcrixQ2POIGp+8
rJwuh9r0J95dU3I0NVRvTYJIYEU1jyX5TPlr3noGnyPkOWJWBILrm2/f+Sl+aYAY
d/XQe5MjsO8omrraZB9bevA3zhoRI4JZ5f28Qk/ppS1/ER03F5X8VgeU5t2GcaCG
8XijrBgr78FjAbiIGRt22YN7RFxQEELMRXrcJGB9J2mG9eakLGRaX2KGm3WhZznV
Q051PbRp3thRmXUrVktU2gsGpMsq8VIr5sKQchouYKIa90M4LkAJlFLCLQkkxrML
DIN1ytw3SHE8jAcYL3QROsUHe3FLDfm+6VFuDYwoScG/OH1GM1NQfFX3/eAPxO+2
GcSzlUDbVDUZAdyOR+oKaDZ5zcylUG7xd8MqyubjIqqYrH0Sj4T41e0AodvQ47Ce
MR8hOzUA9TN9TOV9/ueEFSgD0Cjboi+XZFnASRIiVveYiD5R6zbC5KXXoxhR4QDX
1XBs17twtf9pxuEtKTsEafVC5KJNxln07o4U5eE2LQWcNyljiANaCeozxx0JgmVN
a7uS6mmfGmChs2/W1V9m8OzwlP1h5/Y8lJnE1Zmd8JqQjDp3uKZiTBGPMnnt/A6S
0s94hTaNugcpbo6ymQJbqrmOQSERRaXYgEpskZpm9Heoj3zuyQK6PPhhGWfj3xDy
e4xKaAkku5sNR0vLCgBbTIZ6cCFYI2hx5ogfZ48mdnfJ8f1Cbx2HJSKJZD9KFx+z
cRgDbpQ9dq92NOxMEZvYCPSKF1HezrvxGg4/NgQgFebx3xVt5Is8Eq5LmY59npqk
52/0ZF836aY3D8TMNoMOpPsU3rI6q37dVtb5m9GaA3jY5FPCd5KzES+Q6/ycCvo/
uQCN6elp98HRCX3MWU869WtLpTtMK3n23p2U0VqlaSK2Z+lycowpvWdxGzL3QEvn
zD+saifq+3i0cmA29jPYLXgTDLMgj9lLfaNFbcdDxPV7q6Ctr1x3oVQomK4QNIfE
aeCKHOab9hreNFiUD7/6MMhfQDuGoONKLsIKRSv80pt4Hte+uKkkcvOnv0ml65Aq
EKVxRH3quKVKoenzrgxN+PPSC/7Umwe8+wKqZjj48LG1Ex7pfJTZ+sonIQfR/gsI
RBRXew2+Wnx4H3leaVxHtZGYrZ8R0Pb9Ph6otL9IIe7ijJtM+wxpBHLHBpsjuqsn
ntvul25jOd8YSj0qV+bzLjH3L/EAnouNGjOlwc+pspjrM7n6uzrrYLljbv4qKhDx
+p7tkwbn9pu9URjzi9KSVAbaioGLiwVc8hDvx/WublZZW0b2AEBDrEGdOLD7yNEx
LSBZiC0cflzE1VZ7hvlVcF+XOiU44zTIe4GUmCm7+YhcMSwU4xG7foo21Lrthq59
RP6VK+vfVDuLWDaLmCppIe/TGTIZZvDOGy3iDBuNt6hBor6zFGuqRfGjQqhEcoU8
CJuxKOelODPcVcx77EH7jsgsmUt90lYnIu1ZEZ6KVgZmt947uAjLfLFg5p/1SWjP
hPbxozHbU9oF18gol1m7ElER3vatT8n5Efr9Vz/TQWW4ateIZ9MP43wPmNcVAYF5
JMXKbK0rqNFUSqMYT4rNtUL0t30r5XygH1qZ6SQ9qZECocbn5dej58iPsk56e8g3
Im71UvW5beQhg6BFWLGOgRP/P5kegDCxEHXdNQktIQYO4ks60UBXbbkw4CgkYycR
FalZVJnrqhBv9uYXaYcENBZQdcNXtS8K7tjBpTCjNOseyU7dM6Td7Pm7FpFv+ocC
qY2Q9TAbFQ09CSD76EH0knYLcZZ26zO/1KPxp3viYe+ayPPy5GU5lH1BXLeUqMVe
aUCmz4uPofBVJtRf2KzTEuiMddhVkNSBWn1ubNwFhCbUZ1/QRzdBL9uAV31D5AEv
VOz2ZB8+SdIQca82b3pOYgqmDLUkZb86QIezTEmQe9nsAgRnAXXwbqa+goK3JuIU
pKW38aA89wRrO4etbBVfruDqB92wzvegY8oT4UU/XLlDhBxot1r2lJV01AU9/0uw
0FREzFZRe2I36laVwXAXNMZ0TYW4O68d6pkl1nSFdZdFVUgSAgR3G6nomvckngYp
eumozADFEtZOf2Ww3UMEbGukj+6XWm2yAHiYrk1zB49RQXW/5NC2wPJtdtiQ/Aeb
xog5npIffeTDU2kOeZIMYG7/t/mM7B/OpTSNvzE/zREpFaA3ZJxGD/e3uCTB8OeQ
UfaZ/Pc4fVVYNt9LJq2GFpZ66an8qLFjkKNsbQ1PWkxaxZS97JZGaAEKFKaJCzGU
bSwucsTvllKc9QZOvswF6AK4jiRUdScFEdgzHtYJOAFW6aIpQdeBuyc2itxxIwMP
uvDxneyHQqC405eizP9tCPSaLqHWtsvj++cz4Hd348NcPWemCMHJZzPELPFAsVDe
32AOJ1GYCaQOD/tUgXD2Rdf34sAHddKWNradqxwvKT7zgIt6wWtLLBk25Ig96rkB
f0etqmIUJaaIdO7GzoZIAH2qPCX1vrUuy30Efkg5QaAl/WG+gs/pd030y/ALk5Sz
/vEHiWTXd0X2Pu9wYpPJgMPtczI9Q8AsSZamz3gKAaWBAgI65TH/a5FhW/+K/QRD
sfk4N0O1hjhSVFWNEnMDP2pMkPPfK+sWN9EtEv5pAahiQ/xiF18R1yWrwo4pqOSb
CnF4Lnb7sOabseSdvrs9mF7CWppY7aN7rd4JqSVrT4KrVpcKv5YFEcDRtWFbOAc3
vYGSTOQBfBeXtNs7t0brbxAUd1T3cM4uIUIq3a2ZCLvdkrV0QsfsRP80WMCIT+Uk
kGqaPp0ClHIAKAuCLV0jzpSNIvUmJyud7zyqM03m8AsVwYmOSJfAJMx2ywlJbtoA
tNBbNTwd/iBzh6L5JCzDIORRa1Y1fG0OBgH9RXAsXHWwnYw1/iicarkjLl0FRTcy
9bF9aDE+QESzubGyN1x3ahPg68NWGAhGeiFEkC2wvYxWi/WbNUwWmrdzf1rO+JNo
ihM0Jwv68xKyn4h5HngCLhdjlgRUAF6VcQEiTTwVvHDTwe3HxKAoaDDTRicnSmTh
OePaF0n/huYWjo58iMqi+FeLsMKTI2RRr6Hr30K9AXA46LKrXE9L0BJb3KZXdxm2
3TQz4bqMAEaScZAbuiX7c1E6VrX9aPAr4/wqGwjBio4bEApXLgbQzsbIszLjBSRb
M9YXuHaH38FztMalbVaNnJO+z6lDJL/mAsZGS3nsFqMP6xqcVdzHgRfpu+94KVHW
eW+TxZH+hI2TVHYRPVGHwfdm+Xuow1ykAUr5aGv3JOtqqgaLS9zWEIYIUzYRKr98
4vn0bsNgCqA8Rgc1/ihb/GmE2g9vmaOUDcDYk9chpV10nBT1ofmsNIKrYg3HOTsP
GhdR8M61gAMefa7wi7IPE0EFLlJ3eDKTNtWgM+tYwJrVD7on1yRyz6+TaL9KHsCb
o0UMh8GNG34NNGjZNhtF6kSravKnGWIvIIWXKuqwD0scUYEJSUBmuty3GeapLegR
gbfLUBcF+EuciFn5zS1X7iT0xJ22LQAdcNrHixmFEKumW6ySo8hG4z1WACttpTFd
1I4iQ0gkXHCW8bdFSrxSkAhHBBmE4++fXYoHMFimtTuqB6/qiH9sgdKprIjKj7n5
oAYDFzUh4RRk3WekZYEa4RKqR+vXXrOy8hzxAsifuY1yxSdJ6ywWGo9jyrOkRw5w
fVzMXPI6xDtYuiCA4B+8EN3cujRsNolKeMatVDP+Kw4e4C5F3dKIr+EdHMEucYuw
RzGYM9NgJDw4QAfSjzAyZuT7COhj8T6J5QEu4B6Sotmu0CKHo/odPtqWsmZycID3
LN3Mas4ji/QLiOn3Y2z2x4N59FThb/+Ny7r/ngWVsZOPYZtdzh/kIwY9jilx1P78
F3megOupo7aU7FBX0AnRGxEP0kLURIRxM2LM9L5TnvP/o6/USHjZkqDrVsiy+OOH
/tdhn00MqBE3bM7Eh2MKkHsXWb9SsCCpK69+CbMCrxYpypi2U+UkGzb357b1qzCQ
K61ktmrX9LaanQQJgjNWbeLMnNTi+yjHZ38zDvc6pSdX+2VLXBBc7aS2+xrIHp/+
LRcv+pWtDFc9Si83uBkijHqsLA+JiN7ydqR05L6Q4Kw1XIBAwhpEpsPRfIJ7JDXM
gHda0sDh6QdwL7NUNxeaIOnvJTw8SDZX9f83tWFzXQOD4k4mPcRvYT+fZo6+cYPT
kP0SlhpOIVNDjg696C/CLAgfIYJkwPlqo0bgGAVLBDXhGvn4ngApch1gNcfaPWCD
IR6pM4eaBPnHJInPr+EXrMF/sOP1hMbnI0OqA+h5YAvMD5teyK+4GWMAl0KMyi0O
rhXl9f4vDQqN2AvdS+s9aFKUXZGZr5HKvgRFsDcg3uHJ18VvOPabIRdlOCmuaKHs
nscX0YA9bc583e7SzyQ5aRlbGBUTz3OTIgremsagZnvEHjn0KPNC3bHdfAGIGaCM
eiL/hkeyvD7P6yxqHkCMKYSnsmiNUZsDqxkPzRrnwkHicTlDy5V/Lr09qdPLx7qH
F/eSh2P/itcZ+bJX70wBCjjk4ENPpfOKkbRWlMWwI1/PUzZ5OpiPh8HDu4eQouDF
VOIg4LvrLlrTsU9U8hr2/C+eUxLEEbEeF78+ZJsTvHYv4ldsOHoNh+hLYt737ljs
tFKp+Eg+8u5AKKVwCNL14C8khYX9wGUJ7IpFEmhFa4jnlMcYiLUiECy3XB71JfPz
00sEamyoNLdSyaqNxMk6RMzDIJo/2jcByNG6R4V+G58MwI/SCh0lsf7KLuzrWaaI
zll+sHwbz3MJ1DvLuMqzaeBENlGa86FDlNBKZbQTSDa5ywkhomvSePXxheDGzH4h
/lCHEmiTf++AEn5c5PmMORaR4jhRsxZyxV2tSv10UTdrkw1aO7yvTn9GLwBV56A1
ZzZZaRiNOg+Tie7R6f9MrzmJHpV2TWdXzYHMpjpFujNfufRMXWhT3+RG1girO94w
Y/jG8a8lkg0hbQnb76WfAbsjGr1M2YrlyomhifhRbxu7YYP8SbRnwMbvlzjtz1k/
512tGTpnnp574jVOwJuuBv9Y/04UszPw4DEbYHaBGiqM2AhuEVGaRA04KgWHSWQE
GbkWJT2FSmB8foENXuqgqNNMqTDEqiePdXUuo+8a8jiVSBvquY6zKKRUKZes2TMe
5kiV69yRRm3VctyymkuHD9Yg92qu09Vr6067gLuxkWwnn67Qjazvkj0JoAnZBy5K
xk8WzlFY3TAqtaneCn1Xeb/WdgW8rGaqZjTKiIpGM/57rQQjX0xi5CoNetSmqau0
G6HnT8cFpqSXsuyKRZzgJuahBZD0PUm6IlRMOjMlGOIZA1oKPB0zgjsacPTYeXKS
VWRLT9F8nH4gRbEoOarfaE/JNdKrlRXXlBjwfXn1X29kZqo5jOvGKSxkNwqLDdGa
OAVJnxMPFqi5q8hO7qLvICQZdwFh7kyMLVuuqrraV10uNu5uUt2zyP2cW+wSuMzi
EH4bRk93lyUUGITWso5nBH+vAYiwWaiqCK7gxoW4gNr4NDh7WGV6ZCIjjDySF8bT
+wxzaq2lpxzpFhi2Ff/VsTlf+7fRPEBfbBwbOug2qKr/9rZuSmLdtMbUPODKT66a
iJZQ0HscI+uQiLJOTlt4u/gq0Ge5EhP2N4M7nVpB/mQS0kvTRgxXFAAqE+UV3muL
jOVcZ8P2Z0Q31BLfh8ePiYlXG0X5h10dCoWj348Tj12DEkkpxl/IGrTZ+QhcRqli
sJ56wFSveMV259Pet0UjPyL5vVqxZUmcWuE68Ahb8Ud9+C42+qvfw5Tb/uLEywQU
u4Jgbsfw4Zv+yDVS+w9nTXRvgIYmw/l1qQYo8VKtwR4phsT3elnZBeTGHV/8tmIY
eWfp0fFtSh36lYN+y2sDSapLe9tZAIwQ/VrlQGEJHuisiTKMTiLgSXWC79TXQorC
PibHR95AsYpwwDobAdTeEIcxbfWQYFLePAFsGIKkcfjCVwNTHYm+gnJ+nFVky3Ku
Z2U1CBKRtCsF69pTv2ldBnnjdIl+08AGIta+rulpmC/bPrNCGnaFEzKBDn7PcX8g
5B1gSrOzoI+zBL1tJmwSEmZodGOOAuWQSqDAyEpzASt+RXn8n98euY3x5ohJfV2j
9yum90BWHGj2qM9PJhjdabLX7gARq/epESRnnUE2ynqMT8sKpzUxLMcnJ+SLx3wH
jNXLon9+bn0rUaajAaJc5aLcCIkuwpyWihV1F84tmb/Kijg1uvW7ylA2Dtmh5r4P
XEPWtFdF1TX5QXTXHuA074d7Gg3cEUZWC26vmUHHdFYwwJcuw5LMSL+InlBQkuyx
cYtnXYBGPY9r1a+RN2RevpjazX6z3D1lNGBXFb7EjR+yg4AaKBlV32jV2/VZm9Pq
P3dnKZo4i2Mb2rTK0t5FfCBkzeETPCTJ9zf5edTMFZM5pelRu2UIkKUr5HtkR3RY
kzuJmT7OY/wdExEQO2fGrkGD7oVjVUsUful1WNeVJRIHzpQmd7xY3Hn7rceabK6k
/I49JMMHWzJxfSZiu1JS4RPuMvHRkqYWpRek5cUGHDBdT+FRkf+Hrai1LMlIGSy6
Hg9T9+iMKGEWMR3l2CwHmeo+vUQNnrQ1oacs9L2z+ffv2ZG4xMDBYv13/CpVHYC4
y8iDemrk4KA4CKPJoutucNW4NNxSrw1DLymP02nWhoPwwbNVdKNiQ5Zjv8snjrwe
AGZD6Y604hUaBx0iue/p23rQ8HcJUoWj89lgrPWaSXOsSnPFflxuaQraEbzJnBjx
N5NGap81CZYZZ2hx/1JD5xGx/0SUQEeI7+icTfDPvcC8FCxydNnfswQai+4zWPlD
aQruTRljUPpHLuGs7N3Jp64eIs+r9XyWAnZhLxe+NaCe9GJ22p2vYX5ivIK4nmLV
rI949tgwCUuflTBsy3SXKLcn+FfVOEApUkgE3WqrwV1TC4O+3VRRV5sxeJquALGM
ShEXxUzHfpRlnH+kZAF8zhAQWAzbLaJtZoivdbJbHaQTlLn7Me9UQe8iU/ZmxBCn
RTMm4rZ92pxjQp9AvEpnZZj+y6uidFIuTw5x+jXKechpcyCCjTeO2k1he5HrO8NK
O+nZWPyH5o6Oh0c/eRFDqaqB7yjahSywgO7odJo08srax125j29/wJbh/Y/+nEEY
lWOZoBzXUHc/loQVIOtHL5KPX5bFMWL+K+7COsbt8gIsLCMd4wnGM7zMZga9PUqG
8O/1MN8DCHKsusYrXatBqtWaJe3i8/2dQ9G2W27EC2i7mZRQ7Rd5sVg/dStnJVdP
59HwHagmIf18piqehEWPw/ug5lQzmAc2RhF0pIE4NiY+adunpIWsjBnUi36zDMIz
4V563FMRO3yETOqBflTdlMY7mzFFF/B0etgU7GSZGY5D2YG5RJo/y8FjPHqv6M84
4fi+hQwsJhKflRqoJiZX9mLk4AMQ3Ra13Rabd/hliHdLOFxP5xOn/0NVCAG18qA/
EA2LLnCbdc7lmF5338OYHHkSOay/tvmA43Z3UUUFXqBzr5+m3RIOo4hQLRRwFCuY
+u6LfqyAin+hX9OfkIFeihJfkHMjzD2BVBOJXFd+52VIvItAy5Q56dtmPnKTEtIZ
dG7UqUDxIuoyOujqWGqrclfOFMfvhqu7KeDBVhyNMDNxLonbFdTyfTN1RSj1fOg9
U10VwKmY83cxYb6OOdlsy3EPZBfpR/BCAHIaO6beMyHV2ha9EaUlpvWI5eceICXd
Tc90n+2nZuUfh2YP4j62GP3EZmkbaZBMXOziZj+8xvCJGDBdHJoje/LPuqlUAx7G
9XFj7U3qifO/cROjhYHFkKLP77sL7gP5U/9Tc9ePxmXvlnvs6aG87KewxZzaESw5
1NS8B3hvrG6ztApXDm1qqgoFordE1g8XC9Z8J9U33L04AZHAqB9+H/QFmCUJKXtA
pUa1qDLGbrcvjBXTpAm6a8JCw0iPVRViysWzIC92CNI13WjefD6kZScClaUM/gSn
vdyZ7po0OrC8KkKrc1pUVaq5lTYIhfWbll7e2jB2Wt667SI0/2yAAIMe0k9p062d
0u1tgnsAwF1Mba/kArjztkFFmy7GkECgxa2RspDDaAY4gSn7rLs1X/K+DY7Ztg9a
JL/yiq48Os+5l0PIlPBwVRIi1XfMJHpcF8dWxkwAEjEwdIJNp5A768MjWrJ3cdU2
trdKwZfmjaqYVUzivnac17GgxexJ28CJiJmGX9+6wGAJi24miA+Vww3wFeF2mAvo
J72qmWYMx3/5V3nS+sTTUerlZIq69yHDz0c6ke8ApscMEPdR3EBkSU12ZzePefLg
i1GdgprcAJa+4dFQAHQblIDPlryZYNlH8fzfACrokqvDPat+U4bPg4OywUjuGYig
TNaHnAyS6RQ9szLjdJpzGRPQS+DtSX1+UlVRJsA3k6olFvWU3aA/J+GXtbWaWf+r
IUNqKaAAZF1iCxbwu+j/LzLUoVAiH/Q3AHndF1bhM2sQP5kRHMIcZ9E51XhtVvQg
9NG3ypCBDup/LRChCNWFTIkG749VtPtwrMnnqioLwNr8dShRFoVVgg02JrgQPfC1
whDxfldZWN0zVoPEV+gwWRQTIalOpx0D0shV39b/duT9RPB/6G/sMgo5XBBcijRc
pOUE2HbwF+QFFLVq758jUzhEjVGTtohamAPL6B/71QyFoy644n04ud5AsD4JMW3Z
KU/QZn/9+zwAMFwUbkx5boUgtSSQon44VIRMK4tDBIlJrlJGlcCU0PtJFZlyDzdG
QIsl/i8ZSHuB4usr+xRHmO+qC/sjXP8YMDRnbI1J9FqJ54T00P5JUnUzt7wQiYWB
69kLg3G0neLDPhfY5vr+v39MsA3KXaDezffzOJ1p2YB98jx6s0kOXihT2l4914Vl
95Pc7xQeRcJDn3PZsm5Jllg0LHbmFN0ZHtc3kTs6/mYLdTZfUf1qgSxSVkKQx/oR
6lWpjnSRSCwVe9GX/Ict27cN/RjIh3fChTzUq2IO3ileMY2zECzCfiqBX4w+IhPs
coTA9a5PWuYJpHW3N33DHOHlVm4jaLulMnKjvSBdBI57mWDwsPvDowDWkbZjnwW/
CPvHDHNWHMf8O0la62bSw+s4KPK+lR6x1Zx3+OS7+xXdoiY9u685clyh/M1rUH2c
7i48v3x2P/VI6BYU1vp8irHfcw80KvwaTGRjGIAEpB/0KDu5HvclkEy0ajWjcL5V
v67WP2/vF562DZ+kWcWrEnvRgzoUVhiGBeq2+D1kO7oHBToRvQEoOHUjffbQ+4TD
RynR77y4R7qsX/58RbANhHue1AeVNpd8k/ZgZrXQlA6sTKOnpbqjNmZFJXcvDFNe
/HLvl1wUPgCIWK1C0AE+aF6a9PSehRfyi9hPVzQ2PkmGYbGSYn0JE9KszdQEGmLw
bGfB3fxi3MTFdFSDIZBUzokNSfdSqWB7Q8BoA1mn+ABpxizo1SPT5n07VUoSTh6P
QRWBRIlWVe2XoqPrBOThoUAej0HeVRzW21al4UGN/96hgQNIltlg9Gw3/eNyOIPi
7dvRmND8XlbLpa54jx+CpR2eVX/NtOWDZUuCqyQbSohZ2yDm6mjAXUE9lYC8N/Os
SbrfdTnh+pa6/pc1Kwi1RY5pJRJHKdgEWoAFfpu/PUBBRgpZAZouzS1ywB4NRNT9
cJnMqJrT1tSWHhYOVuYYtbG9ziQcXnd7a9D3grVM75B+/FgG9QGKIxbVeeWnABx0
5ixGX/DnErekKSIRUbLwJTwHVtfOoLx5ng3n0ODmBpHclNNtIv+9cm41uNPWBFUU
poRenmsRojYPY8az+0kHENyic122VcfMWPQAAQXHBOMRZ/GazpokMvIbddZ1B/yB
EbiBOt/8n+5gkF2AGFYD06kK9AfYQUdFl1PH6xOwqCgNpNkGlRL1Nx2hH30VUX/w
Lw7y6lyjCk3K3FuqbW6vk/ZfTbTdmjqeDVkSefxZojMsN9iFVTVPUS1rcfNClXA8
RXFtY+jesZOZmWJqFYsyYbzXyWvgqm7CMXIzBbc8zkKDSflLyl5GbSgWyEuQWTqv
VWOzq5/yzE2qL8GSY38fbxQ7BAWtTkLLsZGAKqwEDk97dPdAaxxOEc1q1jWuIyHp
N1+NzZ/JtzpW8W2hLLD4Z6aE99ZTnSqYj7klyZgh27hmmhW/BSN177IYvnW3JbEj
luOBbBJD1BRdTpuwkdwPaYLnWLHbRP/FT6yPXx+pUIC+a62mOM6jQoEskgxXY7aN
vnat9ItYHYenblb6x9uKqW4fl6DvKzBNBtKDOaPDds3HC6FUlrxve/j25qXBZ4Iq
sMJa85XGCfksCGOCl7nghVwmE1BZc0MBnr1AKXJhGTIshBk5nzGilauKYV2c+X/n
IV233VpmkP2jL3Bxhp4AIz9AZbivUdea4J1KNV4D42x1HfNscIK7Zwf1Z/DNknkk
L4rD/jlwmZvH8WKYOtnwNPx5P3kcm+CA5KGWGqmmAPYGFfoGNexzf4RDmXmkgoNc
3vSKWLBwvW+/O1GRa26UhaEjl0DM7Ipw9MFkAbae00mNdzQmRFkstE64elPdQl1D
8vTkov+oLyPpJYlLQrFrPgAOROjGmbK2f1d8VUe+uQocIQci+7gIMBJbjCKwJbLm
zQlJ7QPpGqV74+sMg+yLE2xPMKrM9iklWsFsgeaSCUkGhVH0KO/Z1CSxuczSoWqj
1jzMorlTY5/6KJuMVz4efstkqvKE6ACq2mxI0O6BBiWaAPw9TOoBeb1Rg0GP+19b
ilAtsbk7yTWgICNJiVnLQQq5HwYzNVQ4BY9TCUFd3dw1fIcrfzo0zVmSKR+dnR7j
F3BcyoyAsL0ogR4Q2t+upNXg/VUcTtNAc9FRuKBj13KWXBqspJZiB3SopHQUNKF8
ER+XaZYw2xBnYnxbzuR8UaaoRRo8aohNevDZILhgesMUn9e5OeH5zJuY0AyQfUd+
bySkvI7Xs0F2x2Z05LS76CFy6aG5Aw94qZs9g90MXE/UhkGFnkbNHOo0q/EXCVZe
2RUT6cB7w3F/gFvu4tGUGjmQlIe0pq3aBcXwLDITKOQsRFKGv9FKT8Lap6jwpPW2
sfn1ZWpkQuVkifLkFqiMKEKpRcAgiQpa/pJm6E2Ru4Ab5e2GPCcsF7T/W92/QSEM
vpndtEYsanD0ZijeKHh4UwWceLEALm7ntyjlsIAEJDBXTrYUzdeRZt+W52EOtJD6
4Ce5I5HAUmsRQKIlND4waNBe+61hLQrkm3gmQlCGXGpBXpLQ+cPC6bKGjU7b8ZEj
eUQQBabOsYcKpvEQOW+FBxavMoHwNBImRhb4cci/WwPBTDgMG3L9RDUMQqYmv72b
7ixavV8c+kVlQk9ECmPNEuIbQBfLrrJqOLDYeyFYtvgzCEuh2L6Yj4IpT6EWiWqg
eqeq9NsNtyZt649fZTtdy7MsnvZmEJ1o2DeduttLyaKU0fBeHyiYVn2RxQdp4lbT
qM1+MrQM6ADaS504BAlltF745JrD5uDg7gDDC1KlhkOeyYsQYUKmWyiBBArcfZ1F
JZ/mqaChCOWcwhQwYtbHBJyw+IvTn7CL9eHtzD5gjpR679w2OLk7EUBjSp98qbFc
E2z1YBQn2CXnXKe1d1XwAuZNFXq7uHtc7YNPOiYbm9PZQ5U2jQm+zwyHzdqN6t6Y
pFV2CTZHuBUDV/KeFRKdqFqtM0RNxRdtQNepjBbMK5BG516S0lKso2/FWmXgCAKY
8jPCxmA6jkSnQ9UnEuvupCMeYP7m5uOq17NmnqznQMAhE5LsiSm8BYmAs+m4evyd
mg+lpx5vKmkhn5FJH8dVfVOT7oUN9sqIfEAnqLwpSJUbtuG4GhnetYDbFUuxzFdP
42IIB6GNkL9iuFcrLWz57xFR+5Xc60FzKofu7GxWRv2wOS88qW87MQ3v7OEzHt0m
VITpbRJjq9ihmtCzlORJ0aXIBRhlTfZh7C4wlvk5mIEGA1y0U8jndYP0UDtUBgVx
gAaMaKV7jarg8T6Ho+Kf3Vf7uPxpITTrhq7xNUolTfz50HeCcEIpTuoMW8KChu+W
Rg2R1MVa4FgY3T/XiHdiMhi+DpB5IiZsVuah5TJWR2zYjfjkHWYFu/gkyu1IfBuU
yKMfGxLYXBVD/UnxtMxehmzdVKGsT5Jm+FiA6XunhmuRUoBuYnSLYQtVw21V4IH+
dyfOSVnIkTcA+7FnD3Ub8M0wiKS8H5LJmpdgNaRb5BR8hGDGfWaDZe5PYZT+tgSN
qJe0Rq1N+Nk35mMBnOEqgNbWLJtHFLeMrsE0EF2dTG5YRSmu9C0TCrIfzK2lZPLf
fqHotlCh9KU6M0NscR3MB4aFp6PCOZhknu212HWojh+0J8kw4dstBk/zsze84kxI
HrubUHz8hd/+SgPGCujYhraOW63aF9PgBHoUJXCQWhOGas172F8EJehHcDYianHR
4wHqGnWkQqYf+nzfkrRLOFA7khyUxhb7xxOgWxZh0Hm2fcRm35/Pr4rdNX8OYqRU
ZDDxRTAsEx6j9UxiOrXBc1QkhMoi/hm8mog1wvs0Dg4GJMFYlk4OFIpWcuOoQIi5
rJ7H/ZzmCOdJnCA4OWLs6PiA4oPIbBI+qFU5FyjfP5oibRkmXqn19noE7O8cwffh
XMzQ0TmP3N314Bvhv7nZO6ysUUeHBNoBxZUXioDQOf8CeJdg/opjWGFuW4cmAEjx
/z6LWb1maXP6jJMPu4oxCBFA5TuBU3QrH4wxS11QaSYuHTdxI+IVW+E4hAjvlZRU
TLNhkvg/GRJ0dTbfw8TNISlLFNvkGkdegz6aEW5YxBGsrCKp0KShDXZKk5OeopKu
MJU+M032ZNYIXn7UVgsboaKxrOKnNwyqYhO+S3l6ZROY9DsoGxvbDr/ksDCGO4rX
jTpVnu8YfI7wmF6cYEEell9c6i1j21y8PFAOuTsZWgK2nupMih1d2jsy5Nw0jjQ4
r4Znjokqjf8T84u8Bt3NdK9wpCFvdD22lb9Lu05mxyBm1JIyPuu5t+2sbRyTSDxj
lK1D0qS4lV20/yLYu7SgOKFm5Wo4uTRvePt/KDoPHbmsS3YdY+bxkyOGyy/SxeuC
hDADC8o84P662yRkwD7+nYi0uVCoyCkiogo0Nz49/UxQiaKE7ZZ2Fa01sOeRI0cl
ZtKJao5UbiIMaFa8W8R90Lk+rJu+GdrtN/KhhTK4Jx45/zCjuHxKz13iAjdYC3oG
b1GkbVSAWObQmRtaqUHVlwg2KmadON652Sz4nse/mZsLAM//2ZGKWAO/gJqZBSHw
9B7UEbBBUsXwkSKQ0qyvr3krw6nXQxUG/j30tS/ZCfAcf9T6YnXtS0SlmQybRjFV
SlkFzX0KG591bbP74w4EJl8XmPSqSrb5nmT/MIck34oO8chIv6M0VNFsonx4XtKb
Zn0Hu+WfKXAcSRpCM0krlBhRiB3ppws4pM8vIDU//FnujU+n5tL3NU4FbV48sxnu
M3FTvB+ZD1SL3vifI4XBmMZgh+/gOllzBeZ+KI7by86ljqnoNhmzZig+3GIv0+EB
U7XtFORZFZmYSOypS87f9Dhh1a3ySxi7fdGXf1/g35czlxpKDgVk1rzQuIIg7s1s
ZmCCSYcvVuq00RmPPJbUSFc/Wtnfjt+VvGfd+FCSqzowiKgyS0odFF5Np7vbN+Xl
lL527WCGf0URAMq8PgrcZbgbaP/ufgQwTa9mWTPMxRELI1op3HyxGgtwkCGkjRN1
R1tFO1D5DXED3EpwDIwwIvLtW0iCBuncl0ztdUlqS/dEmY958YGf1z6wVAw8yTp9
+9jdCRqvDJzZ87p/tIXIBef8DaTsBuJ3PQ1UQhb6aLFDt9mxhzq2MxDfc1N/Ex+3
rbEDRHYwmQAW2Jz2sxcIMZQ55LNu8P8GUjebVTwlDoQi4mEFmZimoULSYiraAiGc
wt6ZEXUxm01/QC4uq6LDRJ+vXcEIBfmMoTy18XaOBc381cdI9CuNIdKqEQeLBtXv
HKxNWv7/HVsA8wLUYtlH7t+2mQGeQ4r/11oGcbyWamsr5vvjFNPrtxeEdAdn+Lms
18aU6Fele+vvXCakPUP9BI7UZWTmDLkLeHetl6YT3kclh+JaH2/ffh0Bxvsv8/3w
ob1cov+LeHaxRcWP0uiKPHg1g6TSPnACQbbN3G/1siGaV2nTiv9S8DcGGUPZKpTc
hEt8Veb1ui0bKsgC45Yy+5a/OM+7mcckrAOZukARSFHPbP13ywcBqjLLMEwvrdao
FDP/nKBhmjFDirpf8NKADjaznmKF1igbhnnXu7EvcKEa9uQJ8KSowCJebVQTwh5S
z7IM/QTNMNBWmMRN8/eo2eXeURIRQA0536aYauOWteac/OTuurtn7hQvexp7QoEr
Lk1teviCars9ZGJkzEBBxlHEUPcFfVQIBGt3atcIo+wcoihXGThc5a5FIcoBaXVP
827btPZXF8DnkmELpTgURasnBX1JuFTHNzibxgvS95yx1MmqK88Jmsdw/jZtfs03
uQH+ARm//gw1ntjkkbVKfWdqfjAh7M1PsnwTqQzY2rEgj8E7pVu/S/cvLsXJREu7
jI2AsHq1pGHDbJox4DGq5pen0FJMwg5G6mZYo8b7lOEt1uCFWd1KJhP31PF3zRDM
eMrmFNeS5fmT1T9+V4HV9MxzZVJFW9poycpb+UA4z1QyUq0lf4cGFIGkXA3kRS2F
4WU382yQ0eUU1o/rL7minmtG70ZseF2oaQVzohjmsVMKYUEuKfY+soSHzQ5et6gJ
2iOA6IR7dHmcsqa6tHGctUQkD34ZlbUb7IVPILmJeLKKgvh6w2EyhXUt4K5GHZH4
xIoLn/leYN13aePhGdKRykX5j3+sA3B2t4yn7iF37JTfjhKDAG7QLjBVJPZGlv/3
5vjCJ4cG+UPkhebj/2kQBdQUi1asGi6gBo6/DUG538JJ64j4/Nj6Y/DVAdlUTNem
ttsFH98+uRsMcQ0eKIdfT9zqkRLDADilNUQcrupdbB5Rkv9EJV4tJu4eIjvR4exT
TjU4wJSMD3HSteQ8FAuDhFo5/t3aitSFG5ccsuVAiGIcQxkmsuxqIYbXfP63KdwU
/hxHMKnxpZN/bLN0N5gQ4GHdVk6U6BuC9RbC4a6HqMVAnzQFT4wO15GSWhbAzpl1
Kb4LmRjF26xfR99soy6tQfS8sJsXjqeWKAAAMh7FHzRsmDFier+ripBIFHpmR2FR
NNR/FNiCQ0N6yaAEwodCQ+vxF9mftcPKkTeNKx1nENwprwda5TlJFb7Ler+wXCMf
TS/1ql+4Do2DtLwaeZF252AwQZ7dw2hd5Gnh0t28Nyum4t5VtC3q/ZtvXneFdwei
a/I/OO7nOEQn1YAOTXoqEMUd+hXM/1u7up8CDdFMNP1PaEAhHJ8fz4EXh0cMb5QM
xOWW5ttPl7lf7k812wG3jk3i+RQ7E8Z+/wBOQ7aeh2PLhytBWeADEDUPs5ILkRbB
Dp2Pjv2mW57wbNqEwj2uac/irYiVWwAYI0+UTG1cXwCfBhEFtlOJSLtj50N+2VEL
Y61ZBJN2Vaof5MlyaNRFpvZ0OvesRByWjd+ZjdOViZbp5JLflV06bMLFg9RBkk6n
TGWp5yms2KYq33qB4P27/uWcjKuiF+ovcob+X1X8D0fLxkGKNaR8ySm2CauZzexc
NeC/wUlnKjRWglWRGq+7dAMpyZb0ljIgEuyr8w9c5s2bpp6Uoifnc9ilkTJ472YS
9DjZR+7ALaz63Da4WcTm14uZDmgNBIoW2zuVsNcUzE3UJGa6WejEkrrqxvlyeYfV
pklonzVyGYLAhLdI1nPLudAwNegrVzrJw33bcbB8mCfTBdUHcLJgMNgkVTa+AHez
4V6iS2EqK5aLa/TR7Sh+ZU183DSw3A0cxFSC2t7+nrsyC6PQQbKjXxdINL9Jse/r
P/7AVodYh0atEZqasbEfcOKNwelS75c6Ky9la3uLsgjzDhLSwRTs7sFNldZYsyyP
qICvsYIq4tvIoZjaB946BX/iPidd9mqbEoV+mZHoJQf14sYvGWKDuepi7WRI39RC
Z3xQv1TuSxq41vtB/iuys5y4LeB8P7n5OFRk8XhwllyUlGm1uXfQevFlYWFBP3kz
WTkUchwHFDZFm6NewwCokTHfKpCpEhpHiZj/a2Q3O7M0YzTxmJRZJmkbkHX0di3x
AKkZvV/BIbrY0fAFCMx7+V4VxcPcd0WiLNbRz2LPXH7JjGnqd/nhyeK4DAjy5qs1
4bpLPyvGAW5w//IcStXtiKTYZG+d4BffzPo5JvSj94N3jMOQQZM06C61bDX0wPCE
+2saA5j0OHcXSEQpQJUoiP09F/gWV02StL60Yd0i6K+EBKlPa8JWt/8piwtCDCam
35dpAhL3MJz5JB5RzolZWpn7PJyllgiNM7yItbD/3TIvRC9665owKykKtvEuWwZ0
EJ2u7khwHOVIkvVbEMEpRlonYJ2k1xIm8mXEBPQ/pVddIVg9bxPzSocBC+kcHnSD
pwG4MaTiWGnZiq5C14VCnCGz8v8PQG8a22JldJ58YZmiX1wxRabXcs+DADWgZo2Z
8eE2HC1HFN71eZaeLjxkDHP2F+lfThkSygc/AxpCCDs+HUU6Wpq6ZHSn/IpnBNwc
CQMGgVCcaLPxLfHEbtaP0oaz0U4Qdikwu1bU/zDMynqMsu/MdjBEcnP30SQxwpQE
849q/yZnQEPZtS6E/SW+7ZsbAztmhL/t8TRJDVu1lfi4OI2iImVV92Xcz5HxkLG9
i2M5oVuA81S6oJFQTmZA87dR4akrtf3KMn6jNXlJ8yKzhF2lppr/p4787LEIQOx0
yeh1mC/SDuTzoXsiSuwN02z9ivYxUa4T17ipTxNmVGEPzIpFrzoFYCVTN/S9CGcD
eog0P4oR4HQp4+hU12NESjvIXnAYLHskL0d2AqiR7VvfIc0+5YTbyeIAGFaLYPIR
kKWRYWny+30ByBBwkHt8DNDTIYodeFD/noGSEMcF4FMTmG4VDu5msnyUvYt+Avno
2S7kUCuYPWMXOxIHS8u1ROQWE55Kcgedj6pNO5YmhoTF/uBH5S9R0m2wyYL6rUZq
BQksDsjTMrOlj5oSYbbRu533sIZXcngNgWra4EyGAt+hMqRKKaY/QmMcf2le3pLU
s3t/uRcs3RJ+rfGf6jAHtSn7gQP5VNB5Ejb4NPy6VhYtiZsq6pNm4lCa9adqGAbn
E989EZ0BescTFhEBwiWxXEKoWrsWEe2AEgN8ah+exGxqb8Od82WWs547YIHsCenx
RJ3eImQUbezcPOIOOfQ3YoCw17LaqQqRjD+Cg3J748IgF/Yy4YrWYnKF8Ge0PWst
P92Kv+c5upP0oJZ1oLw3RKS24xGuCELq9O8tTdJzmwy8T7f2J32X0JIMm8cywUL1
Ws/BNbJLGeu7GEDVefJOX8/CramvBYGy4Z7eIw+5uPx8OvuFMmDZKQyBRcodKFk4
ABvLxT9TBv7B/Di7zKguZj7F5eMHfnS4eHTyaXxFBObY92hrjnZqZzbwIqUOQGng
LeRUJBRnFoJSf6ggKRWUhsVZEOw6H1NXdDyPIcr9n+BKewbRegF62uCQc1lrjjkb
FO7+/zzDQDef9VZNBfD1fbU+zWVIQyJEaqT8gARz0kyPjLmISt+pPBAC40AUAfGp
UsJTpgWRWURx2l1c91s0cIrW9JBR7jb42EUdk0VkY7hI8Um8EsZKSwr4sNqAJc4X
rrt8rS25JouY9sDrx9wW3B+r5gn1QA3NjOmjk9OhyPCFhcwgZBTFgriCZsiDRq1j
yHM0Kg43IibHSxP4IPs3NxQTX+bbWCqcHKYUa6BJjX6nephBR6M2B3MVgtGGzH1e
WWBcqDMuEpzlhXxjl0ZIXz/WLDqTG6a3dc4GH8lFChhDgZGlH16fIMNptHvp4kVG
Sk276Qs+id5Ok+6dqD7pv1exUhVq5TPltKnt7v80E+Lnb4WtY1JIbIi+sWvCT/Y1
UOv04tJn2WKjmrVG3wcSexSZWP939PT9VQ8dK9LxdLEA8gkKXgOqSJMI2bKlrPqJ
VzrqybfPAx178mZsN4GQgZ86MYja+dbK5hTP4tsi/MMTnawAeACT07bBbS379c4t
EidhTGUThjd5JvIXUkRxVVxsrr4X5EvHNO+pHg5DTzBPGibUex1g4S9mQC4gWIGe
THsaQdoTD9HtuFwAXbI0kEX5q3E2S9o6zUfesPeGCg7CBHb8pE6GwLfT2QTCHPdG
DBb7I6ovJ8ymfxUyHINcqQI4c5fybXB+h/rAfNz/nnaMuoUD6b+k0qwan5Lrb+I5
GN+u1QJ2fK2askCqhZLCBsmujaF99i9sboVGgLYkdPfRoJPAt5Vtchs62D+2Sed0
va8s4qld4sTcL4/IdZe2Fv0Rvh4+ma78nBdjw0h1PufKzxqiNy9tYkTPRaC58VzV
Ogxhr7R9vTtR96xPMwBhemIR25LBOiTGvDGSj7BBsM6SkXr9xJ0nYXnXqg7PXvP+
l1Q/6rYBph/rodZu/9p2+jBWVymjMfe/YGt02tXak9bK7772aTbL1Dns539MONex
WeaDGdBpeKqgLMN+VuC8uaorr0hD026OMx/3EW8cFH2YtJRVgdiBPDI0W5fsmDcn
M0/HfxJ2zYCBo74puwAPXeP3ho+tNK+MNWNqxYHy4JKSFAr1Bvt5/unLtJjJfUr/
0lDayON3Q0nWENbK7rKC/tQqs5MLSRWoMx+4NqZ/oNbAhZ0+IO1pCwms7fuLuHcv
o8gxESSN67drwfhANCq5JvSjpY8UPas57l1Ap5409q3aiVMLUMsELldxCQJ0//Ha
Kcd/74DkhJ8wT3FYxYK4Ppdbl5CIAXdjUPlJz4TEcCWX7+pITAlMdz3JVnHNg8pM
V7higknLUbiQOgT9Qn0ewNNfWRbBwHxmDlJn5F8JPICSvGbGZlPHEX4vDaUh4xD4
2iB2MCG6qgzI7pk2ZtdnzXvvnKyetu2UhPCzmeAvT1LBPtDU9ulK3yXv+n2lgLgu
ieHlqGTy201pZlkYILRUXKUGuLgD9ZuMrDXulVm7P4OFbQxVQNPeTvE/OioaGZMk
5p0ri1L3aq3+X6+4tdZ1QNJkFkCo7EELg0vSpBT37RRGFJdeb0jz9LeAPk2GfJNQ
8QEcfZHFknG4hNmDenJuDbyUxDMWmiLe9kqAwqbasTvX9B+xKJGLZQc4bnbFFotT
+peAcQk19+7ai4daXNC3meIRzHSPYWZ5AOxXGbfRmYb9UuE6JDgW0czvgvja8kIH
1b91q57lEa/TDL+q0Nu7T6Z+x5eukwy6/C/wQYikcZ3p74CrRSdzEBEDxfarngOv
dUDUkqRvKcGWV/H37jB+kAD5NNzL97M8JC3kQjCA4qrP//YGWI/GK4iPxU0jabVG
wSB5YuSg1h5ky+ADFgQwQN+DX/Jo6KqWQRXadQwmZ6yXtU3gPbImGTHXA/je43bn
cZ6MEaWpDgdzoZSk2TktIPT7hW0f7IQtZeGY7zLmyOhWyMd2u96rI1322WIKAIuI
ETUOjiE2SwdCjoFHPRkji10Pcts2zOYWs2IVPPAeZueWzUuXxUc2oBf/pVrn2gHS
G3oGTH+SlWSCVtr5fjeMcmzprX94lfHf8chQs7PWGws08kFg72YbOF7of2IrSu29
3y1+pMh9oSP2wES6SEnS1LQGLJz9ZCaeyCLqqotTfTZ2tsxQ12vpEMWROvwox7kf
Y8PnIAcbt4sjZKyOrJ3iQk7wc+eeYMhkoYxNeTEBAwbP838Br9FcpBkFXaj4zgTS
Hs62t72Bhec9jfH6adrEFlIb7RnTio58eVJe4f1RffH7Dmvai99SptktjAmyJwCq
7LGj9hvInFuL6kYHs7x8M6dYkmiTKTq5gvV2QpDXXGcVuhTGxh6IrZl6h2UpCy/k
z7WnUj9pBfCljqLGfqgfM8k3dQaQHtqE/3kJIwgT5I9isPG4c/jz0zdpu8hxscBe
hhNhn15UW8nBPkVvrKIOw7Rhbjys5FLiha0xHou1TBMOwWkY8cZvhKdUxFUBEoCr
lWQrrzuGkZnGMqCY5IyJWBlRvHK0Qj8HNbAN92cZY9SRdlybpHw2xb2e/pJhWy0O
GFbIMY2I+tSKafXks2+mkhjOeLNm3SZfEJlL++YUBg3DHNlzuXIAudAf8gKQRgew
RdHEP5vqb5TG6vh0xhqdvNLOA1XEnQxr8S8ufreDHOdVrGe2HXl+87AmPPvI8T7c
KES43371PFL3PpUf4lmDbBjjj/L2hXfNtYn8Yioh4JKUHCFDBkPTd+7q8i9dQJ5O
42jAnHmwtcRPDtlv/3W2rIkOxnm8ZnvMUDez9igqo605oFhohVkFfPogzKEln9b4
NU4vcCvBP+CkBt5y2G5R1n3xjiEOz0gZVBKVjUAWQqNy9gkThTC0QPztW+xQl+22
b549aYj9sKpSloD4C0gRtLwOzcLiLQBK8e0TrgsZb7WLzBq+FSafyDfWAZU6wr57
hatBtaI63I3JQFzpbD5fV9SAONiF8Pz440Kiwrd/MOtDUC+cvHc8vVUE11YGYr7Q
+iHLcdwDBUWDtoXxrn2GLd61DDK6zcuy0yQvrLJYMZlnuyVy6H/p3AVXlln0DQ2k
YQvxrisX7XOkU/NmViDIHTLat4zan/e2ggoX8A4bJWB5pA39BTRzfPYP/1DUHlkU
B4oMoW0owrk+6t49ZJzsZghYMNqbfPGz+xpmTZUU+ojlTSf/zqCA4BZ4k3dn0ANa
rvWob+RvFOb5jC4114m1SlJHV9yD9D7dCRyleAkojBI7CqChrrsdx5OKFgddXahC
f9sxZ6mpZNiH76Wr9wzaRwPe165ok4sg10+QIRzMrMrpE1nC/MiWvm+6kMOvnxUE
Pialds/Jj8EPkx0ZEhJ2FEsks48Pc6xcNzKGo+q9TWA1Oz8uW+zDoZZ/EX3fWhWr
VSoxQmZcw1umBHtUUvq+SIEW7g96arcm11y1qSokzLYOdWSYg91KdAwM8dCjQcNa
KxckXztXDp/ogFaEPFS3jmMZ2t2NY+CRov7HnF/v9lecKkf2zD3kX3ez7i1gkpA2
bYzJYuI0cbB4gfxLt5yhP1dgDs1vNIQG8asqsEjnpitN1dksw3OBd4NIkMD4tGVp
`pragma protect end_protected
