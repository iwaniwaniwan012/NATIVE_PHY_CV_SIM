`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aAwzsGc9agVCEPfKReFp32DjM29qstMg0+9b8Clqgr2gg46fMH2FtfYr2r+M5Xwy
wqI0+1XQ+2zft9B6LB9LJ0HEWMvtCJeaUhf4D7g8Pjmy0EWOCnvSlBoiKEotuOO/
hrXFmNe4C2exZm0DylZhEagEbt8pEJaqFmXY0Hq5EcE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25424)
Y+/hHerrrPXA7W93BtDeiaZZPum2Pl6yg6WvWUAUuUliN/Jk8UQZPpxq4DXDdFQz
vQr3Ypg2jMxoafnWZ1sHPyq29nqa/WKsnlnnjD9Uwzg2ewOGvNQfJZKS3dHVEsj6
3qnfmDGy9s3L/86K0/wWg0NmQWkmZm2xeZtJHOqEC+1WabSTRfvpV6cBdjFyUOgD
lVGIhirrg11I9dhyqW65SErCBxBisMtQOcV4rA/8OuEsNOfvmBTxZ65dV5k0Eh0k
ATYmXMTC/5gjimO5owCAfTUzxI9Ml+bumey7qzZ8AosVCBTiBRwWCn/a/m2hOEf4
91JdmZUFf8h6X9QOrfmLl7fgBq4o6f6youGzEsQFGwutJG10tmf1Pu01m4/NQ1ap
bYH/oCL6AiCCHu8lzzKOt/e6vYgFPTTbBpASqp6xLxZYFwRn1pqvOA0vGlno6b1J
Nhsr20dTzVkjCFSsGMvBhICOxGMd43yZVEmd8sCay5toND7DR9vstXNOSxr85uxK
3SrkVfcpsjKJjI93iCgnFL01Eqm++M7pXnf1LKL3qwimFKHdzKGPcgozdp9kX90s
T5ku6NbAPYhBOPrR6n+ul6BrjoLeYH04AwgozwG4/wIEyPzQ9MYje1S+4Ubv7K7x
0aBu7QYmZpjrhBdYHcHhrxcpGSvxC+uU+EChN4gX4/AmOskiu3XPWkyPb34DHpxU
hYJ44u6hACO89WHl+uI8B29tjMt7sVEfN2YdwXwmL3cOiuyRsog1fXdf/HlzEOJu
TDX3/QLuhmCAQPSd544CMZIHI5RzVyKkX2wL8KCXBdfehTRrvOUTzUkFSJMLhNJq
H9ZOwVGuiM/H/76Z7dt82ksLN2BRXbU1k41aFcKAgEUubQMBh/4RRV9j+JbkdUP9
xcW9g+Beg8KHVuyLrbzfQbIoShZzMnlUrdnOK5W5FPMGs3lyD3ZYesM3lcwPAkXC
sdeMd90DP1cUsGTOPBgmulGWy907ejgbAsp099n9y7e1C2RXLK1r3uRFww7gmVen
9lSnlRTmgfdeTwkavguBWNqlfkdF7K66MI0ESg2rjHH2fSkkOIPBtHImJubkGik5
mA1xiKyMUZGsnT44AS9WcOAYhCFYjA3IawMwW/CugoAcNTTANLxUdy/M9cCguPra
QdR7NF003+d5jXcjpa3QcFcu72El+zpXilrcmhHBiBSZgBw65E2haiN5+fhkk6H0
+rcJ52HgT2G4peyAX45sfcB/JJuGED0PLKrM5HWtBkLTFOY8wvtWwo2BsHRjItOp
+pU3ZEVmQrkkuL9Nv2/t+icp/DxESAFp6hAspgANoJF6v/WYHPZAg3T2TwhUYWfG
9pUdNJu/W1Wo6vn9HZ2G8w4jJWLMSzI+gT/vpNrsebKJRTlucNDxv2N0Oaz3HKTc
Jdv64DlQpSSMUNqc4uGMCKOR/9AcRMoNUhnJRoD7E99TsdAPXe4lPbuwYfpXJoJC
OwdS1RAD3Dh23qtTPsd5XCqAzTFCiH9t9sdcFWmHujr6RrteKsd7+z+wzRRNIFLm
OvT6KYU72W/3uBrTha7k73tteY6iscZK1kFhtjhlMwb0jbI4z6WEsyVy3+zhJGDb
sACVFzUwakARA5YPtNG0gKLnkCWXI8Nzo65tqibP5IMcowDOI00e43Qd/r75qvKY
JPbqpC3TW3R8fZZmcHhu3KhkhJkYUBQV2axcekAsloK9KJmBF4zJtq5zUItvj4A1
lP3PhgOoIIsNWIfmYSTdZTUc9LPaJSbi3nyZlD1YOVyGId+hgujuSQ85ntu6/d9z
L+B6sI8ih0STzsJpCw+RtI/kV/PjtqoShOa27dhbqprh+5g6DJMCxkRIjlUA9MiN
OW6ELQhdOf7Y5SIn3ueCNStaKwDa1KWamYvPrUnfP9KJ3TQgxoutcmeH3iEGbY6h
cNl3e/Jz/r2vP2QnE1fDv6r0cP44OvmdLdD5jNjm20PWoHExP0/nqG2VsCAf2zXe
cHa/THQN6u1EJGJPjztRtaIbrk8AOg3ShoNZykGmIxYTBshg30e+M34IusacXika
OxYQObSmKb3uOA4QEi8RQUkh12nK4mme1nXmxPlkkRGR012N+F9ondU6qzvfztnr
ZGDPolIIjRKQ6aI4JnrOa2C8UoWEMqy5aZvy+XYSHlsCSXC0c+CxG95RfOO5kPF1
wqjk8/XDcYs9amWo/CyPifrT6ThGjL1mff1FovccxE8VI9H9LZPYSvaL4SUQbKEJ
nDYcDh0TbXlMwVN9rRRV5pMkLMqdDZxo/FhkPm3YUAh5bsMQmPYjXBOfxKgHqUQg
1RU7Uj9ZHcVTxSFFIMoidhCGOq/zT71A4gsCg4T/9tu6T3Z+OLcRpUKGnaYKYMnX
jcsaX4ydPd7JIEEiY4fZnNnzsOnbfc5/EwXiuTBU0VTPw0u5TM7KJoftHnLtAPge
oHPoRvK/LtQ7wXebYIEYrtRrIo1+z5QiQoNbxiBfEV8JtxKPPzzEHW0Q1wACvqSZ
CfX38xuEE+8SNBVLZDzEJXF79ui5R4ZSFZ/goItdcZRaSMTl4oUkb7BcStL1Y3EB
F/oQ1w3xcyCVzFNjgQIBPZ3c/0LSjlYPyzPOWnOpnW6Tjs4Td8WLxSJgWDAqE8ib
o3asWuEi+ZlP8RuvM4cc3Z7MeM9r5LmKccvRNqDhzCgowLsB0WCg7AB1t8+g+z2b
0W682RfDcJ4EuWjrASXKAhlzb6M3GPir1eFOQ+TcuffwIqtirGCyIab2ZNFa1xFL
1SugSV3gKlB+QPpLEX/CRuP6VGW2XuD+tkFL/J5ZpkPgtHdz1kZmfv/CmEZavXKv
Fxyk3t4tTKXUMiFXzm1uutkpcU64UwglZtQmELh4YQI5gfQ5JBDMk4tWuudltaHN
jcVGWAoJvcWJiFABp/66y1S5AJpBKdSGI0JteRW4ksWysMzGmM1STRU3hAp7Z9Dp
H7dHuWmcgZ7ec9pleMlL6vc0zhpGLLqmJVIHhErIL77wl81qWoWnXi8LPkSxQt3G
yrhkI2aVihFM+Zc5Hr3nry7xPnwF1LTyByPtTLkDL+OCNKkbV+Vl0hXcUtiZ6p4G
Beg279thkWurVW2ZHXoD8tG2k/wkgGwR8BrlfLL6lspIz4wA2F/UCGUUQviEBpgJ
xuzlYFgonbnWi/bf+fiCGkP9RDYWj8RNK9ej4UTWUgYAW5pzZh5USzA4WIYTVTtj
NvtHTJgFgGxzkxBEvqt82CcBDDI7b4XWm9QnrG06bZkAGwEbngRpHmdpiTIOjjHH
oqS323lcNjlS1POs9UeLPeiJrmbIJr4bLg8jEzAWUhQXw6qXI4m1nTCxUlRkfgZ+
zUXvOM53I0W5XlHKvOnA4w2i/06M0xGJGl2aj8h8pSNmnTwrljQy2Nsw4ddQs+xT
cZWXOsSh0udNw9an03OSHrHaNZmP7g5OkaFMgsoTkmSqDfmyM7jwHGX57JWwGZIL
Ma/6DNf62BeIr/PfMnanfMIM6KXZCnQAhEWeBQ+5YhTBvrtfPeyp/s/WJ0yRJSw4
58UshlaKmsLAfb+DbWzfmIIN+MbazuRNuqRNO1xkU1ckjPq/+1E/bh8dHzGX4zpC
clb1BmEa+HdwjR2Kvjglk4JoM6TCFbB6EoGJgmN6FTb4fsFW1srIjv2go5y3uAko
qzPihCA5D8o5WpNxVD4jLCRVhw3Fr3HVx27Zi3r+IKQEvFYpbW91ewBCxkWxkuQ5
+4iINa0R3Di5cIa9bVYKmX/zfTHux6HXFgAmIyzb8QkDF5RmkE/XM6m2iPXAEGwM
UuBCpSPdX3kTR9CwOK3XxlUCIEqb26ZN/GMzkut5a/Nt+vDLJN8rCy8Ep+1PvxMK
kDt3zSSyXQEoGvO61ma3OBz5YolKhC/0RtnPFPfuvNbtjhBne+73gUHVJMGPJhV5
3yy8HYfKzebGNUWEIQfPwSEB8oqidewLam+FL7+IH6Gx4+fBljF/wGbzlE0dCXKi
w+jdQIunfhfkJQmCJvOwUmYj8xHm+ToMeuc19JrsEPNcFJEtiVZ4A/uRpyme16J4
4tcmVrSZj/iaT/1xQYKSImmyB3LWZqA0y+6+53qfqv7kGdVINuOFG7aET627zd9N
H+LROyyDlG+1LcyfBLpRROdnej0PUYhFyDwfeWqiwiv5FFewNuMxD/MVw8gdCthO
gimcAW9tTSIuYhUvCpiAdluQA6WFjrDesHFujVm0y0SjSDMHWdo/ihtlU1B+gg92
eZsdsgpKLx8656y1448+U1ypK8IRWUfZnAWQ10ccLgMsXRjg3Tf12aaXG6s+Mtq6
rK682159KIZnoKnFWD3gUhULNvJwlsiLulpabnw29NYb4vY5yOGMgAcOW8dz+gHZ
uvAaer7gcSAsYNAOok46dNeppBedVhugA1f2G8g/vimRcOPdkrRqGntI/MBYW2Yr
hFYGTC9NXyP9+nI5o7gDOHa/OjUgZvGNo7AlKCEKWQHgT5sPmPHzX3j6lOSa3IG0
ZXTRPwR5k3Xyg3ERKkKTorfdUkZAmoxDJYm0RZbdVnbbg4uowlQFW6WU1vQtOO7M
UonLPlg8VVxRzVg6FA8KvaEF88Cg7MBwgiQXo1YXtYjd7TbL63mI34u/iNiZ1NIS
QUOrXdPCWyXZcIV3PoSMbY78CtrrDo1nHgekhkmo+2c7t01xv3VbSeBq7kjBoGDN
cdKr1sXn13Z22W0RSCdj5v/cw/4NKzk35EvdN5895uTMNsAJXJOriDjrAmWoFzhC
3mwIwtOzpYbU6J6z9VYpMmr4D5gdsOAwSRxAbUItHfPZ11F/zKfF0o3ZYEUqWtQd
tBP3Lyp2/25CBJ8+6z4PcWms+SeSAezl521Ckv7BCsSUq1YqfsfZ8zVOtu+oQFc9
ZMbKZ5E1YeixbOWswy5fOAczputd3bG4cxpC4rNhvhDogEVlB2eUFWvtw9nTcav6
Wj5kRDm3IKMFWE4RHoEUnIH+9gpdG0JeRO0FRANvl7SMKmG3/7cuLfqmKzp3N4vf
OnCeQ1GnHp4TVZ8Vcs+pnJJqOUOZYXGfLdyA6bm8WTC1ZPqhlul7k5KnONadSNKD
GvO7r8qrYHyX4JhxeE4Xtd4qDy54yOuPGgSxoj8YCicYoz9BR34t2FXX66K9wYdR
t7IdaYagbQySkVGp3j8JTuR6PDwcM19u1SsfqJL+MRItqC5MDCUdzCGJVJLb5Z4O
WnX5n7e2cs/ColjUes81wFekNAScLXW302vWsJZDkpNLeeg4/bmxkvI/9EKu1FIU
Kt8lJkkcOvRL4U53LF4K5JNAL2DGXlHli7MfezTFq7OOBD4vzkZNq9zkIn5avlCA
b5E6b4FsFI1wq0O4DwGspKa/d8UnN28XgM6JvGSKJuMZs1m8mMbuXmzCDs24u3dI
AfOuIVUGnKkMoQond8sLcFTtgpcSsIluy0QxbqKFkwHYLthweX6fwPo9+m9YWUXv
nTMHaVgKA5qjVhfxATrEv/4w/3Ty9qBzNJON0QJVIahVqiLUCPIdiMWZMi6K+Me9
demigZ5aMziuwUZmIC+tvfgY+lBvnHG5eGxF0pnzOohm6VI1gQYYHTJfnuxdQMrN
P5tpvQ11PKwjt/DxJ2QsNp0lDNItxCqIsAr+FaczkiPVAGtYCXUZgkKHqnSBn4QZ
ALYrGfljDrUSP8K8vF+t3RxRsHrbkDm5kp3yY76TfzXlQXGRg5PUp6GVbhaWtZ+z
mmuT9WO0vcstPC7dATKvPP8eHnmMwUA0KY6wrnRoUT9H6nxhAd5A7jo2t1YCOD9b
q5jykDg2LtbOaqSWgasigL6gBYxOpRw9bn8etaX96m4E7gfayx/49GcM85CmYYck
x9DlJqtaMVSevPeooo83T7Q4xYwi+hJlpxvRW6He3QBka7yKFrLxzULwCA8BP/HU
qBw/no7aMXoXunzBLNNzYu4rGE6bwZ/0xbgoaPJtj746VT3GTQ9M7auftQduC6KR
tFb5VC0Yax6mNFoU9AmsVR+hSVTefICFjCMPj5ZXZ6FCM522IoT+E+MI1ezMT/VP
5tWFsiemWY2phT+LpcKAMFy+IL0AJdrStiR7yG8X+MYttJ+yK7ScWpp8zcofGneR
SkNOSljPsIH512wf7mT0tWZLLVGFuxhePJhlwig9Xkgda0JykJpowJwhsg5yAtm1
QyDa2/0+R7XzUdDAaHgaxT33slAwR4+5AWRhXrkwGBdEBkHmLErus2D5R/1RLV3Q
o3bZksRHSJZCymo4hW3WQM62VKbaSd/MAxmGcVRNzIuV9JQirrx/lZBB7Im25hIs
b1SVAukKjCP8iVdiyqROY6ZOMLtYafb86fq53SeUkvQO++T1MJ4i4Ku5XRMY+UKg
5VGTGFfu8V3x7qisnyRDA3LadjxxNDobIFhEk9vWAod9AMWrLcwcUfTWL9X8hRxR
lQ0mJEy5/rjQ8MnZ8Wg9EyOxh2bx0fHnhjKm5MN1qZI6uFZ9fh31Uc/Gil8ypU77
uquD70uzL7fpch0NRbr20kj0F/GtB11h/Sv1Zktov0erkR8bd27a5IAgZV96+daO
2EuHL6kGvszKBgN42aVPJ/AMPxREOVS4BRg0O3A6hlUbrEip2EdazhHopgtCZ0As
HsBJ/LRPuU64yiIIjwbu9hXFwZSe+p5cG3XUY9QHXs6R3aBE4IkuU0rdJUW2BBQL
WmJecXLj3v9pbOqh/8dUioOkkpX9qn+pwGZKVU0CMweIFXyw33jSRxEGCYDyJLAI
xfYVigm//axCcvUuyCjp67IQcNhy/d6qaJ9XEEmU0rV8PHVGDd/ht16zFPQTqvAS
h7/sKjhvlTSCeQKgVUMWBLDs/tp3RMoO7naMk+I1HI6+LHkB3AuFSu2REj4c4g0H
jd4xwlGMB8PJNFdMnnbEzaMR1tPyJBaxWAAymBomx35ak2leLrE6Gxt6KJSgeY6y
nyBAvmKhrKPgJZsERp/ZSmOdQJ5nHm+/FRrD3IgGVwWoo7FW93BQYSFslCtrQ8Lk
hoD0AUDZj3G6o2J8OLAc6nLVO/zOuAds1bN5gSUMjG4XWxUveUyUfEpU6CGW8OKl
yXg/UGQnvfWg67Nnzcpa4plaeGf87HLeh1UaJ5mLG1Bx1DSwhzmGf8tDa+S+iaXj
LXFU3h4ttR8Ck5q/tGTiPObPRQu2cTyQwFg6OyQnArGJUgF6Hjh68luAQ9pCI4bq
AUzz7aQKTXqr9TuBNVD55bbAgqzRk1kNfG+Y8C3Lft96F/GiobbxRjI7/vVRz2GK
JV9iwhTXq8eqzSsyQTgK5FZ4s4UFBNwLttzbIdFsKoxq8WcLmTR8OCkGmxtzfwRF
rYFv6IEk1jAsNHFRx2cdUJ54BDHC/qJrkBGJ7a2Le6oc7tzTbGgYWLe+fxMckdN/
VcUm7um7KFTmhqWCxf9KHidrT448u/mGQB/T49BNysjHZD38p/sWZMDSmG0vVwLc
YY08lw896QwRueRHZMqCLLWrpddtoJbtyiK8nBo/rKO7Q+pEBfiqt/w3eMvaGgCK
CPMeJc9YJhGG7QAHpARrLKtVzc+rI86fHYBgL7+erfAB16F+fIKy06WjWTSDlOPL
mpoPWXeyF7eRxefGST0cSlM0Kjrw+YEI+EyEp6Qmh0M6uv8hmdVXJrlAjra2YQ9s
OjDQZASGnv2EhPPcPFvuTqMQsotMiAGsbD4pBE4CmzF7x/iTnyMeKPRR24U4x2SC
X+9E6mLxf8mLBw00rRmh01eT2VoGBunw9qLITRtMm+iCYtLqh95TZ7Am5sFcRx2X
qyTudpy+esgzg38AwofOJRZHzeU9Yb6evhelbVPBIblO1sKnoLZfZBLJtziTbWli
Ghn2tyS4RhqXQF7EiJ73Qf2fWwrTuD6TXBl/0B/CG0x/1xbo0mIcbMIWgM5E1BAA
ahYmzktkiL0MGi+u4yD2RfrdEYYWibko3tJbDkAaXnZ51fEqV36iRK9RSJFs8iPb
LsGO8gf958PsBoePBVH4sayqZRXik7AAPbUe8GSwpBcW+5gHwSTpYPKjxvwLHFnL
lUQpZeBoSme7sediEDy2EeEXiMFCmSHx004pzAMbZ6NPcjTlIF0xLg2AY7zgL7uT
85EcMXvg0KaduhWkc6kQsNefk3l49F5Cg1zNZNzDc8qF3dcTgUBI4M2ZjwBctB4v
b8Ou1z9E6NLGso/Y1kfr1xyfraR6xM/epY1PIv84zXwAD+zCvDz3T2I0PRs/ZW+0
77zYS32/gBedUG1PpkUTlYdwUnHelmchdndpuKGc99Ksb7zN416C5FK/1zG16Ivu
aKjfiKtkNlpUz1OILMbQWMM/DMuqP7VISroG5CaFuU8mCZjXGogy0IDl81rx5EuV
AfmIcwOflwR3DBH5gHxBaUXZZT5AvdBuib89xzp0/23AMT8k0AGeEw5Uqmi726jh
o+LyHKv6X2OVabmuG3UN8FVw8J2S7L+vsjjqFPb+TXhVglLw3w1ikStabPnD8eza
5Hyg07x1T2nKiD6sK7RyYkEvJaVOgUuRJ0Y64GxpcuqGSVcFde62CgfAtfIakTrF
FSB+H8Bx2WjQbC8I0JzsVgdELhqJ3e5uqVTxLBMSf1kAPLiJ5Q4G7qWn6TeUyCZE
vD3UbrhlRBuuolQsaSG048pGcL9kI8+FVl72dNnsZQFo+lk2Vj9DrYfz08WnNfsY
Bf8aT2ee+es4ViE9Sjkace4p+n5c47JF0HWvopbspyjh4GyDy7fSlX2GfJ9rFgue
ugi//FlHbq0MwzzVgVN5tfR8FAGbRZwl/sT0WIXdHznOtLX39NqqN+ptCuYpasRk
o5cR3I9Sv/bOuOu+1GXzerno0zVgZCHCeRFvxt7vrU7VermyZ0jzC/lKnSu9c/GF
nWwJvy0MCfqDq8Ov3ZQ1JxT8md0ogX7mqpz/FpCzYbX2wRnHhDajTzQJv0BsTu4R
c+ewCsls+2UaBa7wEVobG40W0O43NtpOs4vBckjSxo1D/UzwQUxhv9+h6mDxgW2g
C46XdCOMJUfwZvITxsdUIq+i/5xlxSn+UdAVOl1WJ0D+ALjjaRB5PuOBhbWUT9WL
YDrIh+OH9gXITcK+a7RN8LA7HYh1MCjtbz+6+V9PbMEh1vo0zjEqkWKByCnUV6Pk
1rNDWW8wkqokdlVdHY7WQnawaoIyHhxs0gExkdH8p0HppdgjHWu44O9l/cTZ34iz
PuOxo7UgCxecfd9fqo6VXmdAPg5O45oNUyFqdzr1P8uIlULKWIcYWEZt+8pWUEZz
4O8mJFYpA8AfvVmy0uKb2U6Itv1KYnUTbyT5Fx/2y1Qty01+WBYJBrCPefuEo6z7
/VIh8IifulldB3bLCbo9y+7txOqp4zbVaXOw+f3F/weoM4bhVEJckk3cORXwCa0N
V8Cj1CnN3x+XGEEpMjH8llcn45vwi0DxYqg/jSL7kEoiBvHk7Co1vQz8bVoGwdkO
i1v1Y+JIN1xvfae4dQbgvYmo4+wWij9wZhDMeGpnaXCWW2F0VQ0WMwHAs0ATzEJ4
935/8pJ/3zi3puiMTuHD6CEKDzbFZ2N1x6HVBLf1XQxgFTZgZq6Id5yJuZQHAgNd
IaaPmA87hOWOfK+mU1sPTlqaTB1ljHb4bx+d/zYWirweMO8CE5c24+VQkGSepwSA
Jt92SH4AoZodgntPGolXIYyEMCUo1V2SnFiRZYr+w6S6VJgWIVDb0tuPCAwPONdG
JYkF02EIW//BS5TV+6FoeOVAHnLydwYiSrMnN8eRgWL3ZtEaNIHzdL1dw0l9axA/
R2I4OPNhrhu4cpysZFz7Jux1EhBFSZWVKXq4ZoTpHq1osSkEwgxY2FZo6GR2ww0c
Zv3S6tuMlsG+JVOU0o63E0YHlw9f/yb7lE2I13l6aDxtiAP7Dz3XG2fth6EDOWoz
bPsL5q0K7CPCPmbNF9F8SB063WtDVgZjuBAOfpEJtv/tKpPKGhTtEm/pIqgCI/SN
uG9Str9kpZRow5zNtdE0cOPtePbCQkZVENiS+v4mq3iea37hEZIc8Ba8c0WYzNcK
JtQhvBm4QgkunGTcrCBkZUblmrSIM8vwvwMVu/+Nd3yfpuPDVc2+h+1xkD0650uD
g2brz4PWjrqDLRSEqqS4iQO0TRr1Q5Xg3EKTmsYeSB8J2gohwld1rTybEmfIEHDC
sQ5NP0bDCeqXWQPu/gHw4C61Bc69KUc0xevRWk74XqqJwJnG6yY4Q5cR0f2/tY26
r4oDQx8emZ7F5TyZIRJvsgtjzlpwwZ6I/7hGVoM90ZDTge+Fk9mlCHqOOLozN/Kn
LmlRYjkAIK7fYrxBJtWTqiw22PWgtIlDv7cHrjNA5DWH6VMplFxVbSWAAPJlvQ03
gaeepRC/2Z7v18MTi4mUOeRLhbC9B3hS51cht/61WWY3mWHhQW+iJ87kgyLbL8pD
mR7EvyeG4mxc/V1FARFGHENn0iVGFRBGE61cZZWyfPeVAcVgnarcSI/QphRjnywJ
ZrtWaXx77pektbYPHdjOwR+0y9ECoiIuGX1QfFkyzHr845B4EVKU9GTLFqJRiT+P
1EWRrvO72mVU52S9bTn7wLoHE/HNuPpxgN5xFyyNDC9rTraANh96iXZ4biKjjTra
dxDfvdwjgW0BThPFAqxtdBD6QJML8qCG2ggISyTg1LIEkKj9UbqU4ScmZA9zZtVs
UMlHduGurjjiPTPDQjjAuAqUUwRQb4W+d9O8J/tPwZb3IrYmIV4AIf5YLmaaRlrv
kY7HKNsJ+PwestmCzl4t6h1JeTmUR2wddbkYwk41Xt75T6ljwQxuK+qCzouljl4t
Uw7onCsRvhCF7UGxkESSgiqbgZ/SCs6z6hygGdogZkZq9rRKVZAJ0wuRUjYnOsDI
sdKYgXInx+9Aipv8s5vSlhfHU9YqgMJ9gfZu8+52aNP7yF5RvjmE47SL8kucfR6v
uXa6xm4BqhLrEWagel742nWJJ0Oduy2vP+bAyEw7uNgmT/bLkmz6KFtE7DeAg1U+
//a1SMGa+wNVhjXJUmNyI6KC4nkJ5rXVXUOWJklQiGX/+LypiNM1snp5Fr7ZFC70
Xwh905pbH6qrF0/W/We5pko8LmC4Ev8IBP6/DdmD1CaaEMz4FjVZSUfpq1qEd5CH
UxgzhQW7ePl2XJf9lnuPniMm+ZDvQTcXDu3kGbG4w2Efl5Cs5zULW4f1iRRYCP9K
vImksZQSayIqpi9fXh1oKoIYR0nJBeHV2sQ5RVOj0UnBK70B99snGUeQbyiKbB2S
tOQOpMDeqJeJB8GrFwPXyc2oZdUWDV7JUlEirX+zg2WIxd+mbNdFyBCV/3Le+zsU
KBcyVE2ophZch5h7PGeQycLVqg8jTlzdABa3e6IkRTCmWP5Je9j0FM27GijRzQJB
LhofhNii2lroV2JNc2yMupBK8ryWRI8lrbuHov8ZxYkPHs1CRf8pRE0pw5wIMD+d
BtnYOaQM/Upwhsq+gPFfVOlinkwcdo1hKOywHS6xJOL/DZyw3/XH6SapchmlY8LG
HHNIl0XGuSygRTd0SqYywScrb2YiKXFzH5hsuZCGaDZQWKFkQaTeyuM+LNJVmRNO
1g8zvZnbdb44Lln+sisfOFsT59/gMBmwYUlpmOMnQGihJ2RjNori6p+3iUxDvLeY
jj8VItEAoTSjUoZSVG9Qkv3hdrCRHEsDru0ELQZq/F+xoYBnME1hDYcemlBiq30w
kXL/fEYCa8xX2Rhp1NG5QITfuqLQYY8zyZtrdMntg1hg9oEkD3Zw2XC66CfvQBKe
KdAxw23VdoTButeCr2TAcfYujjfOr1PAHnEuoI0YvYxtoZ1U6XL0zeYNdrMLvlzK
HsGGyoKkJ0t0b0bvF7+tQjtQeIAC16DBNtG4HCaCyGqa1kz3q9h1zVP4zewh2zVd
7VgQcMWr96F4fZdyHM+S4reYkHdqJWxc5gqMBatdG1Hna9LN3wHnEq7sOFWMHABR
B/fzC85Peuzdu6yDpRqs15awnQ9QMxJ06U3D1vHLmo1nqToJe73fJAk92BwsUz8D
x9c8hI8EpZ5/m/9R3NpKbODki20zjPKwk/fdvIaYIQ32ObNHkZVIVI+HMFizQZkk
BD8cKdVolwW2Nik1b/73/qZnfe3mYRpjn7nsi62Jmpi2DW+t9wMm+RfnyP4iuPhH
w/ajgFd4UAhinVBxwg0EWFJYbBo+IFhxcSkanEsHawoT2PbnKhMdUmeDWTbpqsyT
tr2g2j02XXle0iko0w6iIkZDA6syfrvR9kG/nXKOh7k34pSSE/iS2SG2AHvwgOZk
SJl7Q/ZFnjPM1JAd1GpT7DI6edcsHUXJrakHwVlataWQGTWd0wCwPaRL1vUlsFkA
rmtiHjJan2lCrqXfJpoUm4oEFXheeb66iS1nDlay6wFwOtx4KtWesCeO/3x/E0Ia
AWfxtqgC1FysAiRY7z0E8Jr65Z6NVKYVQr9ekJ9DTCD/+HvzEFJXOv5O8ZeVJiXK
hL3RVczF426d0UNQotIybX6VmeKuVuh9PW4OW4x0n+gce34tXzwSNVzvjEXkEEwo
RZlSF/WCBtCaZX7FlAT2xsHJRxZfItpBAJKxoCuKIHc9+grJSrGVqtgFypg3nreN
cYoIZOH+rzttAVxRezTPeeisjjcxgK2DzhmyX5vRu50czCLbzWsB8TbSGEgVLX3T
3mSqfJitdkRZoVwiStTuVv5K1C8TAY7G0CjBHwxU+kkbnZusY7qfYcrdddF/m8Z2
agxnx7wOGoifrAU0dBYvse6dPPbWmltnQQvaSZeHcx+und/YD1k5JT/wsHxwFM1/
AEO8Gw5qgC79ejeT5/0GYLP5Pmk3dLJ6w9iVJMm3SFLklZt2s1AyIsog9rIIWN+A
tODPtmDAwKonctYTjabXrNCQcxmy8oVHiGR3+kvmUBWtz0S3YLEwMxfyhCSSdWx6
EpRY2X3lKyI5JvRIiKZyDd3cUi96+GQIDwyq6Jkz3mLOoYJZ2kRLdiFtvoDqKhPM
cvFo+s5dQmTKPs9WsOHcu/xqXDN0as6nZhMx9Yl2Wi0/eXeZ3i83IJCUDMKtZ5U8
qkq96hqt8Z+IX92HAGJ1fDLiNrBZC6vO3H0pdYPPMY8G0NbhkAs3orqfe0Pxzp/4
HU8dlR8MYzqvMvrs6+IOm/25JL76GjFqo6OSlaYcSpEJGfecj4bg/YjFMnJOAJdA
++x4ZzwkiDekRJTXKEr0VPNy+gdB8b20YADAKkeq+05BdVtLQ/RdFZPjzk3W4+9J
QO1j9Z+wVxrjPbhLMcb1wXcVRBuPKb9AFBeuWtUleV7mKnsqikaQzRGDBiuDmcJv
wkwOBEs0wyPAV0HlblzFLNK76AWwpPy8G0TrO1gIPohusqgoMnsrrQu+zhT938e6
uWpcLASTiocUP5bQ2wzeyy6LH2sbEEWlCxxOL+aXM9EAqizv21Gf7nHnT5xvpZ0h
WMQg4D9mXmIGmsFiM5UGfsMRXGYEMjbMSz++6KVReDfGtAnpTvFI9LstnCAtw8wq
MTh1twb+97EpcH4w15DWkj68744F1H114aLmOGtw2PPKt7CzfWQWvQVH2kvgFxLN
W5dL6HVGz+XZDb4mWvmrnDIMtBZMWZH+DK1Ahox4tHghtQnwPMgJX0ZLqf8zJ7sO
siAUAuWyEvoRXa1ajuX+HC4l4TSmu25pTZzMiM/oHF+QUuI5qHy2Rvsyn3umk0On
3LOS6roISsR2wXE4c7WiNCeAv/eg75cLoRDyyeWH7zKAIZzhrgeF2A8JEU9zYXtN
Ogl6NFD8zF/dN23JZZUaXq/SSbZ5UqVQy0feTE8AMmfHf6Ud0GtieT+4XyJo88Co
gaJOM8CDm2EWBjpXVR7GTsMo6+nle7OSzsVLCPqk7okYxOCTPfHNfSvn4/GtCDs2
dPuShXiHqcVwfuDigNjQ6ixUS5oqHyoCXuYJdTyT3Qmovo2FTcWDEXEgZ8m3jXv0
2vOfY+LaATyxhbYIz/rfPSHbZnPXDSRj62Xxiz/bhedJiCN6Jr2TykZG70wmQ7We
wI5YMsvOiSITUGX0sRqjxz7Nc/CmrSL6Rdrmb1IJNcwCo1Y+L+bS130KzJs+asMo
e3E/jgZVISLuNLmJ7qSCQKJAZSjR7APNRJs7MfvfBtBDkcEqAyvRaVPRMUgAYCMN
/fm2z94No5ev1u0kwJ/GCVrgBQPJUTSfQMwOJZXhth0WHMXdLKaC5EXGKBQEzjsT
wXiluh2dM0A8htwhODmBxa9V5APFV85A+0bL6eI9XLkpe8ZpXzBDg7kBvPSZCsH0
LqLKVmSrK2Lh8oelzPc9dV6ZbUiKt7zPerREYPh2JnhDS5hFH/hFGm1VxinIt4TG
gyqAXIR2OPJux4ma6DnkDGI9lyNNzaFPqL7sBQp4wTNLDV18+O2YOqC0D0qPEs6p
JIVpwVRJawP0jNxkl452OnV9QCoPhrYyP7XDvtucKqT+/N0Srji2Bq+j+rwIeVUx
s9KneMXhBarjMfMJDnvRXMD8DGNoI0N/xvGc5mUSd8iyZxbp9Us3vZkPquTRvOnp
e1hiOBVXDur8UDhJ8NCXVFbx3FCh1eLCOWRPQmZoosfe3TJZVX5wHz/xDKqQA86G
pUhbLVn/1GIgmlsSb+Kh0RewAmYe5GGxEXSbQXXLgM2zcb1NJ61YEoAe16D5hXWt
CPyf8EX3w+iP1jgWPLhBlAw/bS2P9ZNfZhyu7LahTl/fYvfST9nDwpVR1DiCuyk1
OFLg06SEWEKcI0KY4R1NPjhcBWlrkVjFewTHBNCHu/iC42aZoQ7jmGddBgQS4R0G
uYxC2IjrvoCveUIVrrsKlFh8tr5VPaMw7NZiCSdBUcLtkB34m++y4LLFX4mdtNoZ
JIJU8it5GQbV7h7d9gH03TqAeiTR941eMQwsPyCdpVEMv/NLeUtkMI9U+oISJDcX
2m+pjsJgBBwum4azN0SxYkIXLaUwtThLaX4h1D8QlWX0C5B8iiBFLq6eDYre/stu
gfXJjOvyHHMGRn52yBUhGxBRNi397S/OaVQMC+6bhxIzRy+IooZAAo9ZXyHYtVfs
arATzX4svx36Y8sWQ5HfhPwZq5CSB+/tb/s3rfylg3hBFlsw8Cn/w5WWdkcvbogg
Gfviw0tBr55tWElQ+tNXrOkFSFtXVkNx5Lzljo84CAupoe3l9cNNVqNsbIGQiS1U
O5id4tF06uqcaqF73GZ+FiQzDjQ6g3exzMht2bygckuq0a1QAhh7ePEKlQOnEa5H
O2z+E1pc8aTlNv4+H8QTeosuwnTUptRA15oXeA9fLkhmoAJG9W4wBJf8q8yxFBAu
3bmSWiCCWYjz3kRgviG8HC471xNhq7oGOT3jCrmVVYXBbwMSXWemEDb45ItE3XmX
NpK9BR6sSGgni8/Heg6GDEtv6nSXIjKMkllR2KlFIcqO8MnbQjYfs9Cl8hXjKdl3
Iy/3wXgcNoqCqKwc8UkcsqMN9uQt7l8fUlSdi05pkRJ2M8FuIr+4VqYa8QHXBi+Z
9tjZXJ74x6laytdI/ShzTPxRHRY1T4RG2A8DvXR+no/CClEfrm9yy1V2ThuUWMUf
gYNZXPysr35q1PBWnkyvnE5QLwtj47iZnv5JAI0vSS5QENZcg4SyI+lGTVU/iihm
+JMmEIerVFQBEHyTYczB/1PvLXXmV7yG4dsPow0QvTo8TI2laCrrqXXDXIyLleKe
eXDxnxaEJS/78d2xSS15TvNcaqOcqhlwVzVo+8kpf3IhfCmjDijtYxftnENZw0uV
VNFG6eNhvvLBMUIO+KFzcRh+9D7v/CTF0mjm1FcNt49RZkmlWyM+tVRp25VHXQxT
N3W9Qj0M3tBwEQUwYMF5NsFqdVvPhtxYmfJswDyqXDKGBZnutvo9dVClr+AHin4y
T0SwE0P6NJt2tVi7jKpeKfei/zpUZ9KNa+w8V/6/bK3XmgQIxeNT+/ztA9IiLG9G
dpiSy0asPmsNKeVUh5+y2uTRYqFLbp5NuOEqKnTFr35KqgZJ2JnMPgzfQ3WsBfSW
YNSS2ExYJIAY8dwdDGw41VZoGX0TwrLJA2RQgHOmqAGpHivibAyGrhal+rkVmfDw
npgSFH7NO+ntxn0qTDSAYWbR95vGogAL9kMr968pM+khsPH6gCkOCfExogwMvqu/
Lk81OhDUP4+3oMP83GjBkA86wYr0JY5i61I8qhlZ/vAoJUUx+RqKQmB/BFSyV8Wi
bO/O4H4FRtc0VrPRlAqVTrn1aO04E67rnf7sO04hn9zT5eMtfPmqfdG8F7YFyXqE
f0AOwOSLOvunf9ppRYHKgXf/3i5n7O+tzPr4PeScs/KK/B1n9R7B5E3GBYijqSoX
Ctd5k7OMtc2XX+YYJxGZ1vnu7f/MT7dYwjIKLqtXyoMfpiK7B/CbFV2+lu9IXBiL
ce5fbVzaWUD5NHm+wb/RIh3zsRH6jD3BQceeCye/2WI9Pr08Yp1SDhAeJSopLAXK
92slaik0/IpiLHunILg5x6nXMVy2/Um2wZBoKWgykd72wOzA/Fj4DHgopms4SPYD
bn58CsFZt4BaGuBsnqxHKoqRgg6kKGdwHCIuwWz32kP8aGeKgN7rORI820ltuuxv
SR5yke9dZETMMaMN8BLuE2EmxHqtcGe53NrYoNojjb1yr8v3f9Cs2vA/YmLgdjbe
Trr5Yb+W8wv744FsBpGbjpI4pALTqyDYK3jC+NYLfqbt88RZoQW909GJgGZtnEJ0
hqN2Pa4W90bhc+kAWwoml/951OdFVjvb5lDOWH00Kbi6DpfLfwn3qML9zO4TgEWF
NIJLoJEdyr7YyFYEDxEG0Ufa26m4Wn+P9UKCbG7EOq3vOSoLYkyKLCxs+mwAUpWM
QAGFLtNPvYwrPyLQHo/GPC5BWFJP/7zJ1WzrEjvzlMNdGbxziRHYW98bi3jwV0V7
j2P+Zo14BI2j1cz6+e160zJaaTEKOD4h/sdV5ujvmlJ119W+b/NqLHscs0F2a1PG
Saa2glAiVHSzHX3zlMg/QP8i5XRTCXp9yc/J2iUPFz6Esh1JrtQpeMYAEirWut0k
qS5UaYZy+OsNbREi/6KHVY5IMjotI0S0/UFzsxY/jpZab9W9pkqnj/2CtIrvql3X
iEVmZ28RE+7Nqrc4wvrkoe5dmTUWBbL2maAD3OChDKRnxZoPnPGfG7Gv+TVCfq/W
KHutHyk+LrHKY6CJooOYnb4kkMvF0ILI1DEnIfCYnTNeoQnt9NtbfrYiwjnWsDxY
skcl+iHf4rn+hg0SLgHvdz8Ec57MWeQn8jxKYAtxTcS1WGr/R4QS8RbbFf9AbkRm
Xfy/RVN7pmqKsZqAY0Z/bKqNp0VaMBjxRwhusA3xOXzhzHcOfhbdBWIqP6P8B9kl
v4lRIjGFisuhDbc97gK7FpHtKUCvL0ON1pZXn53pjrB/qVMEF+w8qgBAlAJiZva1
EOEpPU/6l5Ix6OKNGoP2TRRtT3tZZr6YJ/aSj7GVgE+3AvuABvZWv+RyVsAy/u36
S/xi6DrTdpFsdDyWmkVZKPoy5QllWdeFiUsmnrffHrpyGDCoVZo3YM5vLLo90gyj
C3jp/vSwJMPU228eJACdoIRiT03R7BdRyOH6M0dkbEmsJeIZlOvGBgHlSmybMfr7
ts5XoT0oFuDsiZbF0lfDqNr1TauJD9X5RpZlS7NzyNX/iWa7cLuL7zs71JortjrZ
tkgHhGJFCGfeeOdTKz6NcaxTz3C/pwQHIYWQ4+r4ihkp07Pz5gTjfNvF6i5jsX9z
4AmPtTUk8APBcnrI4LODg8UwIJLGXXzbQdLoIU1jeskUeIWYf4XrLEldiqPeNLIn
TwG+QIc+xHU3DvP4Snu5K38JTec4A+QhGDsMIgWP2P18awJ+19lOhPg0rYP8S//8
BaDDI/D52HC8/ixHIsS7dXZM8qMJSzQ8lEwAnG5cU0EMNfBUJ87QaqSwXQIuvr8c
mq5gdZpnZef3jVs+7JdCKHMVS3c6Z8WX6wv6uMxl/4qJRuy6XtVjN8hbOsBJgw5Q
pbgYPzsnXoQWK6SnEBj9rTKxe0NhLah4PaoK558y2ebXQU/3/8XPRwj42Gg/gNUV
vQ4kXRt2KkHIeke/BNAX602LKc1KgzKWe5CfndhFNyG3FQ2uCQkxFafO7bSBuPoP
9RDgesnuN1NVb5/H1MdoAXJfhVWS0i6TL/suoRkmjVc2FfdYfOBNhk+V84/iLhxl
OeuV87VbBnYq5Xrde4YTQx3j7bcxpWKWpmMuOUplZZO69aJUrCffqjjo3SgQ1BVg
Ss+2pSK3JxHexe+uniJ1T2iY0gXLEfVLzSPsQN20hUhQSsmK8tdUHqKxT3yBlZK9
RVE1HBoSjvfvMTsShAEQ5yc24GKTnD6bb+t3EJ/y6fh/UWFsnlNPfGvq/AO9Lzv6
J5cvFOP995a2Eea+oTjz+RA1hrMBRK5G18/JzWksbagpLQdKQfTRsjvIf786qgwt
TpepQFqodS96WviAZJpsxMkFMoIQ/g5rzkWIEE1AySG6xOuSFQWqJZSM7kKMvI0Q
+GYuhlvK4Kx+5vWwIMa2NkmS9tHrD41ulo+rOQYDXs0Dd75QJRDT/omQ0tOkq7si
5V2Un5IO3VtsWCfNy4tDxld3duJjUGHYHNBeDYdNBDjPk9qdcphdY9k2vfpfKT5B
uWNmC6AS/J4al8LZ7GkwlH+BpgHuAQP0s70ltn1w2YZgAh1p3PZnq16gftpI8YX+
LuLpIrrfxRQCN7BgHuLI09+gvuACfmlH5JXkTT2A/ZGV/fJcU0DgjTTN1Zu+E0P1
wKzzdHEi78uUe/vqcDyfzDyN9fGQSXCP5hibNlLSqBJJzaROSMebz6SzBZJeiFUV
ktsFmWqJHQNYUr69Rr+Xb8WtAQM3+8y9Vy9brESwkfOuzyZMPBEiHHlQlSXOQGTi
St7oIpJIPciqXSUavzShYzUxfxfP5V4+4hPpC4CyXQk+D+vYUxgHxaQQECi3v3+c
qIFc1lNWHX8xVHhHT40ESfcYGU0RVzHqbtSwRSBHIZxzDZfQWIbr/W2dQ+77Tl6z
dKk8XJIRbWtyfSTGGs8rJDmUsYFVPaKPQFO9NqRgvCkH4O8IVINHYHh2i8LeTqYI
ykF8G745ccQWf+r5vJc/czHQp/oQqSJWzkRY3Imb14vq4tmDsdVvuN+4gvxKqzmU
+mZbL+NdYS2UasvJoMcO3amh4QIYzSs7xWTUCeaYpFMp7ccUTMMQmIS9mGbETNtl
+tnGNb86lZ75sDxlYTCS5TWoaYn80r3bWQgO8r3XKqPbR3xsylx71xbu7NvxiSFm
DQ9/NSnqZz59vhy9wJGenHR+XlF+54JfTaP3WiUOIOiEZEy1Cflys2ISkautnl5y
TkJU+Dnq3935iCURnfCOv0EprixNY3yD4XsON1R5iqb3JRE+bjcYSfcfs6+sf/PV
p34IMFLYjtOIPHol0H4qhVqBVoGjs299kA1yWPrBiW8Kn+u7vcTYJhZBA75NV0e8
Gs6K1FGDAXzhEes5zXoODe3CjMVB7Scpmfl+8lpBiL0TFc0YU46qTZPLWRwxb3jL
meb4WviT/Ruvz3ZrbrLgy8af/vJVOZ8GrjcOZlZ1/xAOrw9zEqS1ESyR7X2y6I2a
k6J92aNmcX8TQPWQoBpUHgWj90VYZsOv+0uBo2rTjIjO59P//y+i6+4kUHwDuen6
Cemlpdqy+Xg+cufeJ/tCk6h9pipf+zhk55D3F9b25g21YReg9WD2LeX5LxO1KZrf
RX2q79QtNFOySECqljQ6Yp/LG8rOU8f5l+EwtfPKwJG3JWm7zd+GE7uTO7gOTWBW
EHIIvMs94nljTZiZsY0SwN2pwdUnmD3KTfJDzIeci8Rubq0/9oQOBsWTvcY3B+SX
y6fZJK1Ao019/a7os2Kz9TIBgniPqbLB5mNgxYnPTxm/zkreH15tkXTUXChdIuJM
H+UDUYsQKg8AQeMIxiimDLxBTHdzB1R27+WCeyS3St1Sgn5oSemhW7z9a8wB+Iid
oVuCZ6EodgrvL8RxSg/winn+TvH4kRdhLes1jzV3SOkk1lsIF0Klgs9SSV4ritxb
22v6XdSLXFE/uDfYw2QxAGa77qZF8tjbcxvvE5EA7FYaO9v1IEoxfIIM38fJkYKK
QXPigz1U60FraNWhZB2pa16WZybGWICHPD3CnP0bs9LFJSKHNUqgj4Rde69FRZKn
mdOPD0u1iN9oHtO+FJSz0NnQNs7t+pqdYbrCDszHLm1Ig4FN8g2jMGCtyR2Aljob
hAuDwvqCuBFY9nHTjqlHFsqM13aIvUruk76Kz+OpAU1w9Z4bAhyQurQnVsjXVcaV
qb1ijcDXEZBD3trlD0EsOR4sAmA9KIJyWVfQfw88QufurlonhP0JAkY2ifnaeUXX
9ZO7xzYBGb4t0v04A3bNCVq0fgwG+zP1zH8dP+TThcsR8LKHmSxwT7rP6r/jeiJi
hCoIgNkmXoq12lJFEtM3Ky/Gux9GCwZ2IItRXoigHhM6z9w/yIyZf22p/Gw2ITxz
ZM/WtFQa9PfPzFQ91AvL7hPJybL9CRzKuOFc7MGz520Hk/w9EaTtoKIXchDsdIID
6HiWbC6bRaxEVM7G0if0Qdt1EHtb2xl/ClzXIL3uokXPLEuSxxwlChM2Bo5K1fNl
6MgvVSaiCykbJgYop1wTpi/7LTIGYHL7Uh0EhbL4EFxS2SJ94arp6rwHTGlMT/un
NjGNL5m+9Eo7fCMA+AC9/UfaBq1mSEGLkZNZZIpcaoJU8bh3/w/5CH8e5BjwvMMR
IsR1TwtHwdsbP/faKXtoagIQwe7trmh7aKzmOLgo7L70QQ+mkmmczhEkHE1ce81U
vc5awi0gz5uYNHOPg/9AiPynLDelouFKGk2k3ydQBx8KMRI3gTFdgRteBhWB9Wv3
NX+GqyvwC8UIkQ/lfJm8JJtiVoCQTW0JYjmVX0MfqIWZepMhcQqsqLBQcWSNyvEZ
0UgGKakGnoFZ4OA71+gnQEgkty8RfKn7AYi/YmSjf/1lA+Y08a0S+qy4HK+e/4rY
qEwJeaW594MtdH2Cg/wdpFQ+gXBoIEDRaPJIfyEerfvbM9kRocdEz/9EEM2mLLIg
jJeGKsO3Prchk7bDmQ/69KdHvTZHDrc1V693ZdllQigBM2OqfSGVGZtnsStW1vLj
W4JODmTIV6sCRAcroAX8X87GQx3pUtjk3nx53JKL1+U4Y2GHZiafRE43Qw/MDWEc
5SnpXwXw7rkqO9xYuyx9TOl0frZsejw6GX8U9U8qFMPVZxVyzHJqYF+PHZtOGzqg
SwBFTg9JlQXfsifkdUXs648PuGphxgMP1hW7ZNtD1jHlUYWCtCx6XQeqr/9HUDrX
jVVapLMdb4zeJDJrqk2rxWsk7ftHXcW0o0Ov9qnj4P05/ptLG8UH0nsJuuGN1fXc
fumLOhEKALA6vDw8yB+yz00Qc43KT1zkzpdGU9p0QsuPG95fcfenfHVAjCv09JeQ
VPZHdnhNLdHtOetNMfG7WEbObj139dkfkgPWgA/Ya70XINyYVgKMHNqu6M2+nSHy
X7L8OLlXeRgas2kOWudXHnTfn7HKPGlXPW8YuAoL4waXhrpVCpGOieqIfdbM+aji
gnhr3TRMZUzsgiSReSF1Tebdk3/Aoh2cfWdlXHW5INE9S7prDe4oM9CPyK/eF1KL
BETeH/8cWMSgWe81q7/MHFaCizbH/mJNFP6rGPkMk+ndh4zCSjB9DbNnBxKWPPzD
ceNxVg9dXJLoEIakRV+NrJNs/NFk01YU9sUcakEF5w0rRzLpX//8phWaLyx5wUmb
xLB0UdV8Idc+thrlboBA8oIW43vj3behwqxQTaU8WW2ZR8zSntYVwCF8b02Jua0t
ypDRD1KGFKtsv91u180vyMbKfVfilXxDApdDUwd8FH3bWSVvyEorN+W9RDySnhKh
b4j2eB1HeEBtkNNRlvUyywRXGKOiLT7zCrWyP3MJcXBb2WYIKK4n/nMHr1w5sUFI
/cGcZJVlIo7WfLasIPEuz9NCdoCUWF4ezekqmMJvqcUDrF8ED+2xW++rGcRCczm7
0RHwDU/nw94Rl8oTJVZtxhABBWsUIiiSCjkeSs4WHn9ZIG3uAvaEq1s7jYL/XFa8
njL4RdfXnhz8XQf52c65RQO/QyQoNRuQgWLWKEVqp/vDJJ/IP5/c9fIV7onIlD/L
FocxskV1YgHk3rlJ3OLeQ4Mit9L73DIBWjf3ff+MQg1fdoiiREBRRWw4cYDyCvqj
SL5hvxH98UA2twzT7xDArYEMcTY2ORonV6d7jbCxlL2OT5mnayqF9bdi50pBfG4c
E2UhhYqbomTXfm/bz0qhGu5ybhIeEM1Vr6yFy8fNFxTwh+rFOHfPzKM+KkOpYb99
NUKb5/iEd3y9/C87YhVZkM8tmyfmTLJA+3FUIRAp37Vs9kEJdYzKI2OwcCqvxb4k
ZDGUE88PWfoNo4TEzcAO21rDe8+U70izBI6tb+wEwdpkNjk4OdWXbqBQNV+U0KL4
+GWR5TKZSnCJE1uE+aAmopctkVFBkx+Kh6xvICmXXy9DZxELAMNvB0XR867gU6h6
Jg3apsgtcMDRL1z56rv2CWs0SkKcM4Eyh+Zl7xH4WRL88/r1l1Fsd7P0v/nSIsch
4q+T/sflo3pAzSPl4W8XyNOcmOvb7q8dgXPL6q16VSUmCqR8TvjhEqLdY6O93pGO
mmnwY8c9gIDB6serLzt0RrLCsEGq2Y2l2JircNd0+6lpdAK+2QvM9JQxBhvh8yXv
JBJ+RzlcxH511OtTnl+pWfnvvx83ekYdte+uqw3ulDbpcM3rJAHX0sgso5r8Vf92
CnwndlyalJ/hXMvVGPlqQzxlieDSQOFU0xlS4tqxXb5Njsw5mv/6vZMRZ5Y/jBXx
vam16ps1DFP4fnb0Terk5avawssiH87FcFK8crmpvMBft7liSR0IPnQO581H6BMf
BKP4i0Bqz9Bla6/CVRBv8lGE2Z3tVUiCHcPQ28J5KPO63FBJaYXgx0lznwC7GjFf
7YTcTb1XgwGZjV59suA0nkOHkOBXAqm90sviM7rtKeEvpY+5V7ntiYZ85CTXBJJ/
5wT6wOw38jHDXXig7f1Ny996d4ZcWk+uwumuuI24GpLNQZOp+DDSOgYi5CRvFqO1
OYpxVpysdVUDyRPkEi+OwWreSQ+77iofjfzLo99Lg/eo0epcaBOYULKPV/YREp8F
Z4ANjxinqGUNTu9XzftpdWVmS7JhyHjkUEZpTDtrycpJ+v0Me5FfKVmzBbLSoNMG
x0wuLLt4ES8endDm0SGxSjk1nxumo3BtdWR4WEExZ/hkBAYhG/LRq+DB+pLRaS89
eOX63bEcrr/KHNTIH8F70YINkQ4QbKlzLp/6F76tm2as9CWalMFNBUqd0+99W6up
uZNRFAgk8R8xJMn2ZP4ovemUjjhpj1qJkktLZFAxriTNvot9v/Sn1irX2GJIoV7K
cyZSvJ0igHENsKPdvK2Kmc1IFFwQrHCiPIk4gUF03Jl38sqhYsjMYe+drjt6rhE4
UyW/ebmqFCS8NmlLm/FtwQc50F0EgsaCY3CxInFho5oNuNvstNwZKBdAn64Jq2JN
r4cD6ag0uo1WNtzxdHD79SMNh+YlDFvs4UZpjmNJWgHIzr5cZQQgBlVPX3GTosPX
L7376D97fM42NtRtQ8j0OggWCzCz+XYh493fC9Nqhr4x6etPSNhzR/r33JYnYeCJ
M7+PY5aojy4xNTZfHVJuY70uSCIInxMEjSBTShhcENi+S82Q+GND9u0X/ZpS7NAZ
s8RPoPz5GMWtRNabFw5rHuXL+AF/7/5qOnC4tkoAdo2udLFrmrH06wG9bZggk1et
5VctxR3FNgVsHD2mPZlvb0Q1hKLQPkdjdOZhtF1V9Bscft4nxIkkQyggrCgh6rdL
lNziZpPkJOxCHM680w30gCIj1NTARk3kqxRNJNPr8/NlGpIzugRG7xyDNzNMU2hU
hvym0aU1Uimcox99Z6EG6Xodzx+DlC8bAmaRhRcyliuacvDWLtTV1Vrt2Zw4CaU6
MisDvHxtFtS8x2SElPWXyAvqZLvNTaHk/vPi26/2sw3XTkoa/T6bxA8+ZZ8a+zgB
2nd5km2z2reNebeFkI6ydKUyUZlYsTxSZVJuZ463273xsiE/W3OW+ZOkA/XR6KD3
MrHWMYBhVvM4xnhu3v0hN3FuMhHlIwpEeOf8u/dr8BviqMZEXEPKuOm1lb5l4uI1
iMvALit3W0+rcIDNw9Ywg5KVYQKx+mS1kzTiSL23Yn7sUt+UQaXf9x2ZhoQ5E+S7
9evZK4Op7ftR7CU05XvSjvbR2j9xvCleEAw8KK8Ceh/h5Z5fOwvwbe17PaSUTeSp
9SP2JxDT2I7V4Wl/H+IA5B13/siLOeuS4GTJD4rrs5NPvrD3/gm0YnD1OSuMslng
wwnzoZXUKBwKdguQyxTCH79BL/RvS4FAzj+FO8a52RRoHIhROdp/+j4TiBusYUZs
luU1Df3ZtWBOllEY/VeX07tqrDxL58IosIgRtt9MycrZV+hH9c+4NOYPs5cPjNIv
Ldlc/NlP/iR3DHvcYtbjfzuDttsfCxfgtd+aaEFazPkXCNxqJko3a3i/YsCq2GYO
TzntMRPAkt7jnqaf6QiTBRptP4FyB+uC/XP7X/qRLHqAO5FG8TuW5+axFxWpjPqF
l2fUqGMm9DhpLDG2OSiyHnWyW0G1Qli5u1flTg5q4p16EWsCWMcfOLiAck8WRvtn
jC9QXWzN2Sav7ZROoLih+yLvTq2vW/89ks8Y1JU1qUD6TP7Ibu/Bz7WMHmSbUoVV
jffKV8o0wFok7ZGJiOj+eVRgm2p8egju2UL6rbl7jiKeo9RKg7pdH9lBOeQXVwvL
tlk+DAnIBkNwXuVZP2emXXKJQAeRrEakroCAKRMVgjcQ6OTk3P5YvhfLO6IJpb/E
HSoqvPLpEgnkv7z/gJxOiAg9OQoZw04hDJSrCpMvDpZDQTEu3T2NBgM7u+RYtoK4
9ksdayCPgJL7wiqU+3F0c30L7ah+UfcigSSXBpDyaogA80l16hRagd9qJrhsJ237
n0C0WFF1T7vmA34jsTS2yh+oOJ2fb8Vsf5Kzx3HeB6uUgL8tkRXjI0nfgLUtezXr
03/JwegMG9pyztMwSAp4RRV9oqK3n0aAKYNi7puyAP0qm4+3ZAIUSZ6ojRp1Vg8k
o8f/NAiMtXkGs4/r3rivgXcfOAobk2Zifs0zvgyIvuZiZkYSu8Ej4+XvIr7FLi3m
GcF54xSs93fkUN5wYoHsP2bd+5gd0YtRO3YXmZnakfYO9DSM+uoEqB08h6mUwrGx
xUC8nK8Bx9vAjsokKyJfxWWbLj76kE9x5UHmx/TVl+r6xMnERPvrak38K57HZau6
5bFr9aJr0pOTxFr9y3DQz73iMzvseCaVkgsFTvvvrEV1UG3p5i7xkb9otQJCLTPg
CiTqE9Aufn1nSiAqeRTUQLnTJ4D1q2u1ryB76GJTeAvHQ2SOWy/0jf4K+N5pGle0
Hp0cCQYhNwSuoyeRz6xABicb8QJIAuTFAbAedb2uBhd7orYR+HXDIScenuP9RpvD
rTzUdzZPVXcn2j00Uk0IJ8HmQV1xH5jWnC20RdZwB6UIwM9gg81N/d0LlACUvSAX
lWC1VpdNNw5CHsqd4IOETxv4A6YVyApCz23Nxx9YyWsTFGOr09+oWuRnc29B2e6i
aFkySYS3Bi7loYpIQiH0/s3QNi6bzES8u4gnxHvn34HGESz21nFODEJruPv5zinc
CSnAtF0wAi7h9wEgKfpYeDjaaL0txIH5nkS2RC82xRykYBofkISXqxA0nAJyWzSD
tioti0yizjE2pzMkcn2l5uS+BppN8Vu6R4QGaYA3R6ZoJj29/dfL9506/eDHTVBK
3wsxrU0WCV56ICpnOS9J2qWjKFT7e4ydthKbe8HAB8tD1QR0DfLBwF0LoHNEToD+
3oUrd+Ep9G55ziE9plGnoF78hWBRqn0QJ+M2c/aI/wbnmsQEXeW8mEAkLo4x7GE1
upFLA1ugQNA+pzsZLvFYNoYx8S3z/FTpuANPfGLIJ+Ds+tvJLDTUAINgGyK0COaQ
OPx2cWx2bUwGFBPk2iZ78si3A5+A3vDDy+t7kjBX8oTdu0cAdLA6YV70uwWWEwta
MrXut3NBIO1F2xo2c8+7b840gfe59yDn2bzVs3paszIUtfRQvZ9uW7wgiY9Dz7yM
kH0Lglk4a0MKU/X7e77MgKv/juubqEwcutPoye8Ut7JIGi4YmCCjX9bc4CLLkZHf
CloktVmwXdLJ8Xfvq3/KO4fkd/+oRzWU8VW/23apPEcJaWdM2uHFaWUR7cpd2wkG
iFiXGwKrjAnlZtB4sVPcn1XKKF7Y+fuBwuulg4gttwE2BRVycRafMtV7y0MDVQ1r
XkbH/J0JNFccjh5VDMPY6/wi8coKGRPv6BE4664+rgQiX8qvHI48G33dMI1xawAX
zgnDSjFEOVukFbVZrjX7gyNMATgxUpcBy9cRpiXOwpqyKoBrkDpGd7kT9i/cjBkY
72tkXK3YwUf1vzMww461YKaLSOHxp+uGJoakdvM8okdrEKnMhNbWbfxP6B1wb1v0
RLtvgC1TYnH+TnMQaP8lno391NYAxEkJznGRsn+uGXORU7gYq8TdVVEg6sfnp9oo
I+ygOmy3MXG2Br0XaS/ZVYaLsTxCaZy86fEEq5okZ02+J3Oe0R9bzmdM3ObNSdhb
eCK3t+3MDz94cpGZSC6XhyKKq4O4EehJUgZuMgF9akSk4hAHJoz3ywP/8fBwUs57
EUjJqdltgYQiz6Rx0YYwvdweDNT17pNrP6G554firRWDDpzedgqURGnbVZDvAx6H
a11fYs4h7wYrYf+2XDDAGvzuyY7Cc5f7Pu/VicfuSfFPli26Ni9NllTC70JxsyDY
9BlB99JewFf1B492amWbXubaL9+D8Pt30N4lGObJapc+q2dbWA9AR/cQMcoL1PHn
N3WfXmhr+FagS+RG0X8br+LI59FOmkPZzMZ9SE/4OQJdvWbNOq1DilTdGPlpnc++
pv1YncS98DU7Ehjr/06+YQDrhcvM6M5lH8N/Z/T9YFCFx8QbvB7Dy8yfh1NDCXZy
edB2LvbehjANNzY2cwJ3tidfB8ZLJ1IO1mRH+nx0/2aAYlrouc95sQwys1Y0YL/T
wR2IJt7jyCS8T8zT+h4isjamb/d/XpvOqA05ThWXvwIB3rkrJOwZjv61KtBIeJrV
T2k+0+gi0dNrfLUiIG1+Xabw24+NDEJPiEmwp6iWRlHDfY3Kfo1KmSjOXBlCQXk+
xpR2wLvk5xNSCVv577DQcrhbYgzbA1SHRY67PDdu4u7JLxJ0WLVp6C614AmKRdSk
biWvja634/CUGpx802U5BH+sG9Z9oas+ZDPSuFqDvQ8ArJtv6jpQx65MKexelfvz
WQyT9+Ongbh0/Oe8vQtfgMke88yfmSxEhb6aKA/3wJD+F2umDV3i3K3UzRQVx8w0
xT54yCXJgU1lfk1zeNkgGCkY4vAZn/W1KtJa6WaxQ7zq5ulxdg6d3KP2RcHy55p/
k6GdTB6+gBkQpOG4xDrooZ4l8bff8/CTyIiYDAnKnO+e4Bgg7oRWCTmoR/a9u1Va
/l00ry8qmSlNlpuFe5NNTa42wJZNPmyW/ctJRUEbLxqkD6cLX+63Y5Zy+wkbm2dT
S6yBxQfLsi98P5ILgpTQpg5wrwhnl65Hh+6opq6U/xS6mtFjVRJ5l3LBiYIGWep2
Yl2gxt2Ud4dHWpUm7eMtq4Hk2pHOXFElfCKySWVfJJqufcriJXZjEseKqBFIS3XQ
WRHqyg3kjazuGxt7A/apgYCu3WbPIOlj4USxJme9j0uyWUkuFQG8W1l3+TCXBu+G
oNGp3s3oRr8MC+jhuFSOfEASKFF+tiGsGT+YVem2NGsjmp4aQg7dXBA5Mbu5ho6K
0QejVGeg56XBWSU16HFn6CE5BnB8RRyn6myvJx1h3zR+gtiZ6MDnqpDvt9brlnB/
HsUFX5Gxa/06Tlo6JYgpPahVE/p/4qFlGg84Clf4imk+SnrNg+NcBDnIlZmhRV41
kAkKOIaLCbrv++aklEX20k4VnyGvgjxFexUUxWx5iWTnU1zMdCsIJbuxHb3LpzGT
jUKtGJgaP3r/QJW7/nNlbYgJK6uUnYF7vVRSBEcZc4n3jtaILLydAXRwHHJikziZ
Sy2i3PBSYBongQcOVJVmBJGGS9siSimhf+nRpJcH/DmSZeK9kU9zp7gR+cMZnI7I
AdtiHU99s/Nsi2AuGBFXAtzSf8iupV4SP1LdlVYjgBhnGCYOb8MleUCy9h67ht7x
p6ZF+kYY0YHhe/7KttUgPs/+glYNGA9u+s2rKUy8L+XeES4j9LpisZiN7Fv9uuj0
BVmC8+97VO7tc0GJG5ldFlMkye1ARAF7Il9XrPSdJVsdBZSr3ZMvvKNiIsMw2rmh
JhdbxXDDyUVarOY6DMzFBKevTeHJYDFPlG8TK5BxbbhzQ3CMciZjwWftLKhPtEVU
WeClwUCNtMxu+hRmms1HZOQPTw/0wiq/qIssuA1YSazRz9ZzCkSNB9ThW3PbS1Ip
s0vNhMfmo1ZxUZ9KiuT2nU8C9kLZcWGZQU43GiCHaD0JrURSg7qY7tObEorCqaVm
OirE6S9uqPwxUwqRrODzYfDk1jkX+vUYTnbaHjrDFzhb0KlCxlpNgx7ycsB+oUUi
0S5Zdj0aB9yN/J9zceJ8l9IdD1d3QYs8fCl++M0tCCTurJTU7pnFaqhwBor7rBWZ
rtMn3XsM0S6OG+7DUv2HQDm0wwg0BsDxq77HAAyWvzrAm4ySZaJzcM7fjFzzfXvz
s1s7FU5z8H1uZXvicODEj0gyfG7rB0m7Olk4IwxKpklDKG8y4O5t6okx6E7pKZSB
vgR7pGzuk2LFW6kK5Kze4fGAaWVeNf+95EdMfzU1gs73k/ZW+yZ5tD1wyYYu7JVN
vuaV9Z3y8/MUV9jeaHSGT9946Q8rWkaZJzfKSAMDYcS+JSyoX68RJbfGS8DofSkp
Q8JYaeNNxWGQF6SMStg1R6a53s9LFqkRUEElEbcRTM7BKbT/hQQCt56P8LPYn2CO
clH290Qa8LdCl51Kcd9vhWP6p+IiEmejcltJUg9UQIjB6lo8+EKyd2cuxmegYxtI
uz4db1ByirRz0B//Wjamcfgr7KbVzhBuy+uWM2dHbPoOv2J5saxchihif3pwGB0a
Uio+WNDW3cXexBeqrokWTF5jg1vlGGYh8mhONU21QgK0u97IgQY8i/GXfO3A6uUb
Jsrbg9lMyvWES19IfYE21V3D6O0bW7CHy9chkDbjy5UsxVAngOcKWhp8+/zFRrWK
hNrFKvF9641F3+SV5D4Bsl17j+aHLm5CYcw9ilq4xhQ7Wa9ayjobGGeFR/RzAp0L
LZ+vg5cz6tQP6HvlVvNLztEy8UYcv5j66t1KWvLkwnZrAuOAN1SuQPdI+e1SlNHm
d02/kDhB/2/Ro6n/E9begqBirGDwIHSzPN9NpNYn0fmgmB6b+EPatSJJa/NsLUdl
MiFCqV/sH4QxA1jcmDfzEkJQUoAKBfEy0gLHLleRc6gC2IAjceoPt++/W1DCZkI8
0/lXfLupei3agLboZfF3LT3wmx6C6UV/jmi+e0zD3RWa/vCPdYkLMWr4npsNhjGT
Ywd7C8NxnN6aw4J43nEktyXpUyxfk9sR3fwIq7gntObJmhkvX4VVa2UZtFmDXsdl
ECLMzirHpRNGuyxFPSU+cJIIayD9ANh5ndvW1tmir98rYI1r0tDzFkNdH10QOniR
Bg07xUKOQcRwFbJs7YCAl3jKEoke89CWTgfl5Kk3nV9ngmtWglXlwe8qt+1mKtgt
sXU1qjcDuso1NteajNx9GRfzRt5ORmdIE4PMaj21HlURmKZ1B+8AiSWXvk07T+z2
O+Hf1YjpFRtgIcxyAPolm26yRAU64vngXMP8xlluby8Nq3/EYxYV4yLwE84potSO
pGAMFQvN0v3PW4hw9DM6pPZn99mPy7EArsDFstGNpS8A/rWnL26Eu92nOvxVpu4E
dAp9lWKw3EMwDBE4Nt34NYS6DZC+Y8wgmk5CzAXYF5SCeyQqcTumseY+pxGfKZD3
yga+BNUyRZWUf6fewrNU0pYVuSY1/7n/Wcr4Hy/81vY9ARcYbqw5C4KMd7HI4ws4
g9DuLHwOWi1Lse9v5byw7qH1DiDVTKs2bnoqSJiDX+Vu1HbNUlRn/hR2YxXQA1N0
I9C1Go5cgX6qU4PLaakQ3VpqdIwAZcGdWK/Pnk4SplpBFgdCIILx6YdQtZQDT9hq
c7LlqGCeQ73gHAkziIrIgUqZzY6G8I94tseu84oLq3M6lJglKWlik4yP8mLhY78+
p1GtF7LG4E0SFecOANDz8Nd3HNGum9xCqcugLhWr7M4LOVxwWu+2lUnIwtduFOp6
AedJzV1GuQTpx9OGz0x5fG73plwcvE5hOfGnS7buSnSzYAK7LSgUljRdgapsGA/B
ssbabyG88NRkRvEPc2NoMBp87kQtNoQXoKymJ/ABzyokbki9C1qsEJHswJbqP/hM
X4PMOYA/7oacPUYE1JsieZ/G/WrJ0/JHmrBvsxl6da7vQVE1tJCLoqhdBsrJpy07
D6pNa63C/yCvA0Uq9YteuXFZ0E0tKIeY6b5xW9+6aRMOqMLP2MlSnmWhExJ+K8Mu
Y3aJ5mjYgKgwJOPYcbdWgZm/jOJ+KJ1rFPalq5Lb5oTVg+anE0Lfx3zK01Mm0uMP
5q95zzaf2Kfe3G9S1aYxJBYUtMcE2XA6nAlf/jmG0I6KweFcIceJDCd33NR49KyM
XCtPxmcgw4p/4r2PyYcGR2Y5LFWbUb4xGI5XPWciMU2plqKlgi5EcESkVGmAPNOC
13T9snpVNY7wgVWpkcGvm2KNG4zbc4PngvLBIdVsVjqRM0pP5I8f07Tl2YkqeCVh
ZxD4oU9gQtjf5OGHGfRrb09x3DiUT4lGYZa7lJkAv3Hd4g5+ZuYqfdGLkAfUhgll
5XBIgHE018nsq4Olrcc0YOvEQfZO2Av0HKBiuqJHPSHjoSaB77RM8NVGBcpdZQAe
8XmvE+LBTNdeDMTs1ECfiAz6lTqK6egKw7BZq4u06ZADe0vk8WyqPkODo3bTJc8f
fJ1glRPZPWBD+oYKl85EMRMSSmX66jbBNXyEva3On3urj8MlGNiXHD7IPGd4Dzbt
wmic3LNmbm4SsGpM/B7hAI4zMeCCHDDh2MpRE5awUcvZkflehUcGZul2xPgnwH0V
oqwNAGfjzUX4gV+/sVagR9W+AD80qSQkXO9MK3C2La1fzD+eWjbvYr8zYhURRXuk
UC08lD0E2RFp562NfyIzBAeVDUJnAbLeRUmYAWHxAxZBAZ3LVDDZOO/VDV1Ed80D
XImZObPA8KJi2C7+IuAl5kmMmFE+dOMtRnWdToVVzZv8WY/fTLS1x51jOd1vzpKL
VhhjYCtPq30DIoN8KWrReIwuVquAk2gePhibSyoEi82H5+6koLf8+Gifr+XQPQJu
Nr9TFffCkCr06JvpqlsXwJ7Ke3vmjYGAuYRm/U5S/Q1aeP+MKA6EYJMTD8bHSSyw
YCdqO1LjVWiXXqlvoMniys/2rgtQyvmb+dKW9kfI5iBAQDyChKFkEFIofAUA89lh
YoLBW1mNaiuPYDyVu4xYuEWwzYnLAjx3cFcwXIOQyw1FKK8ipUlo7y0SfNApszL/
0GSDsSNQ/vCEJhA8ZvecOqYUJfHCaIathkZIv1LJyJCvRZ6Rv3u7/unSm7Nz4pC3
dfZEWSO7uFc5DDZ/6HjrN1+Ir+RTZBYLwcKnRR0Rw8O8CvHHCypreZ2PvZeQXmyi
gEpnBVf8WG8v+sDTFuJCOsJYjvTvui+NCFWuENeM3Y2dxqqGyX8aJ9kKsAONSDmw
fetoGWK8wsUBjHU/NZARPkrUkNU71L4/l4F6ffA9yjRHm5YBQisGFVBX5vDHri6g
cFcxY292+WAkhuatmz3SwPWuZG08kU+4o+7yNJNX9fPPpf1iSDIKDu0n+q48XrIk
HdXx6Y9zvZN7V8t+4oniBDX2VQCnRDSCnfd/OSgT13e+ICKIZOij7BDunelWaYuv
bNFl09N2N8DU8XPQN+9pmPCcHxlUrTHWdmWlI9PMi+EXgr4eb7daKsmQSUltwkiW
6HrcmutIEx3enT5yL2bfZb0E3StpCCE63ovOUjdlDcEdYLdA77B5Hx43Z+BUgYBh
TO+j8Iywu5uO9tiXTQ2/1YNhWwYI6ocqsn53gmQ9Q6r60v17JmONIv9WaTZT0IO2
MMqItBBL3MT+HjdQxng2diY0trkrrn7GXEDLsVIrV/Z/18UPj4GBfmp7Lx9cBNjy
oxwtOGcr+u3KqMGPlwG68CiA7ynIdLdQXayBGofYh6/OmFxEfhylpZ0iMPvXcFhm
yVwGKENLqo/g1uLESV97aXS9uRkNs8S3+YFkGFD8TZvflsC2YvPKxuLLwulOG43A
/Cqqm+mR1tMoaZAFDxtO3Si0t3PTB0+I8gF5E2JlqJeUvGBZRGgMSCCA+tvvub5r
dxABVHUTD3NnJenxeuomJ7lm26bN9sJH+GTg5JJfG4MDciUKggK1Z4wQkaxBBbS+
d9MKqXOKRFRkHUTTI+2xYsv1tvXlSopk01X4tp5C55iDCiXoZ1ERexdK8IfzjpVh
edx/+B9FVZAoZhD6dW6O58Oxn3bO0yLapyzYdi34UF/pKHLQ7Dkmeh9NA66EG007
taNrVx0JkPJs1Y6SNSJI9MEUs0+Vgtaf0imSAnDl7czdkWOksZEm1hV9yVJ5DwJC
g+cMsvJPRY8QbCwK+40AUQuX0FC8F/0RPgUOM4APbO5kMslVEV2fqOr0T7MMcpES
/abLqnCLVDFUPKMW+5gWguu54ieLVSIksJ7hBfeTsgdH2o3s7cYoCdvJK0LvGN7s
lpEICK/BBVIUJ0a+JB3mwtPLe4DxQTS5FMEn/Dr7sZ3yeS+90RNXz0B+XsV1Iou+
dcWGpRljftbU0sq/kOMiBsQF48V2GsYnivqVW/I6+T2tX95iLmanWwFMLI05p6ot
b6To86ZuqkOAdcYNJHJHMIbSb2sP+SvYT5oCQy1cB6WzP3WM0/XOsww7webPWJw+
jvc7UbxH0hwQWtcifuRWX+CITZohWMrgUMY+7OF1a1T/akBceP8k/+wZuUrqaxaq
DjwOh8ztgrVoyGdpr7Ww/BfrWmxl1KkrYAxB/9N4LkPCEJW1uX619wFaW/OD4JGJ
cpqzYZNcyI+ygZAPvw6cpOZGsjkYDhyk/Sv7hNK2KzA1IAdEvGBGar7qvXaayDhC
teq5GuH4aZa9JhDjrCPrc6RT+BPjp08ynATnrc3tFr2KFWjyg/9wIUDw0BSPfzEU
8HIV7P8c1haqCci/VKbrY9n+j9hzzxR8OFeBoIn6BJZIe5ELb31cziT9OacHpjKg
dKWYV6IS5FxDJU7E4nCFs5vys7LMgE+O7ZKYxaEa2H9K54rHY6GgH2RMpmRFKl1F
DyrSB5eg4MTcIzCYxMyS5K1W0ldBmPhqA1RyZClmkBUjDfrpPFi+oVHZHuhfNiCK
VfWEd+X18DG0hzm9Th7+xCfSvlx6884gDk8KbCiWMRGWvh5MbpEScl63XA3ulFPO
LKJviL0TKdx83JEkJuWtV6Pzbfw4UI27OqiodEhhpN2HvP1OAuLl98iUp7kre0Di
KcWtX9QrxRgLq2D7OEjZ91pIkmCWLzIRBCnqFpjv7gJ3A9P7U4novOzuzGpG9vdC
Rx+Uwxf11TXzos5XQ8ICQlVveBHgVmlnF9IwPL+R8bnHX4+xyLbjmtnDWh0B7X0y
+WNqirM309Ake8jFEPQKkcvAhIZv21fECUTKThGYFNmnu9PuHhN3VpbDZFF6xoBp
tSn5qSnNloUOTjXGTAeBne0AgCs/VrBID58Hu6I3uN3qzEEqfMVUglnla/3krk95
A32l/uOQIR1Y7vvoUcsxDalQU+qFcWfFt76apAZWWh0=
`pragma protect end_protected
