`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gn24P9koJob4hvM8rP/KwDjWnb2ygEXhlQd46QeeGN+vzwGdUmATK/m6BIJsl0jr
Y7tHXTwhy1T+saZXgA4Jar7GDmi9fYCh4yEvnR40ZT+dPxZvcLjuLaTR1ooz10s4
y8MBUKIgsvHQpqj7LqXrwHq/1oR1pbPhyJ9XIlKSWhE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2176)
QwpxgF6jR2wg4VqbZRXLTOqz8jy1VyyKpRkvnGQsTbvfAr/ET3GHziVHsBMBUEfm
+Gr1WnuEmG6lCWg6VclDAAGgSw7om3WEVwUMK09/+daiBKLwMFjBQf+x2nm3J/nJ
L37jWE+Jg/NbXMKSfBvL3yLliRk6j0RQCkOxb6MLXISyrem34Rz2MZa1WovK6Tqn
wTCB6n+gC4LGAeXAku4IRzlAXG9t3Ech/0IcHe1PG8Yg7GkXuTvqBuXqaWcRzeEY
GxBo781qP9Xb+FwLwaB10V8hn2/qgzR+WMPxm2FGNFQ8WJiJeBLdSJzaun4C7CQw
dmYVt1TbeoVDXPhy68WbuNxxzv5RXocJeAAytlX7PjS37m/jOI8AFekZ5SdLA1CQ
yAzXEiLMDAbynZCblJQu2kbkOhfa0dTPS0GOZzR/7AxmwQcphQdgWF9AfdDqbs3C
9RrxEMoVAsqn0p2IebYOdyurVuBQXYq04V4Lecbsyrt/ACFOQDGiT4HyaASildUz
avpy8mq8JkOBtr8TPMdGJGp4z03CqWwstsAkCmOmB1aoiDf2syPE7wtSJUH9mGrB
VDArejEXuVIavoCvQnlbqjzoKdDZjr/zFTZ3JFCzxKl0iaKBsFlAW0h1Lnd/VmF4
hY9Vi6MvbFy5yrDTLL29UgWiNdW+ubLRmds/DBeYJ6LbWmkr5KJNt0dQVDuTounc
lNt+NPsf9bnrW0jPdFk7qI331b2nML0QxoDsloL+bGT42UqdvUaCsQtJEk6bN7Yv
59npDa50PjsrHobmFqQ3c6qYPVe5sIjSeDdt+0M+NKqg2nJZuaI0daobb7FWtsYb
kFcuxcSh99noPM3MxA31rLMAys5RypXsMj2iJOaqm5rpUffpoqLGGJHCtJXqMvcu
j2+OSVrKhZTgpo//H0NWo2RTWYDLOe9V06CWSg0h7LhGo7P9AX3y3GHKDVg4gh7V
gf2/rkoxk9ql8Z7Xvq5L3XqvAfbyijGbXdhcpvAgyBpCCg+WfLAesBWNvnHWT34k
+AqjjdVjGaKnqI0zNEbcJRHL6dWwrtdVSC7Xq1xvi6etY2h13y5h3ZBaoraXUjYZ
DwfgyeENfG6Z2PxT6sGDJdS39tNLKYxLtEwzMmBswyzmVk2RFo5/P9I0VLRxOJNC
yUpSrDVO14CzC+Agos0xtQ4lAT038FoBPAsm/JoMdSDpIlKCNZjsaugiNnmrGlxS
hBMX77/kx/M9fh0T14jdPhCPO4sOAZZPo1jefYuY97K/cYBDynCcYp6Morg0mGDY
a1jKCgli1CSMdFMVeN6SoJCy1Uv+bncpIMTqMcGARe8jUKTiTixFmWZJIYeVWSgY
9aDzdJmJ/EiBOldDelMgtuHpNMEquFuWWhmgt4G3bswEt3ev3h1oidOAph1puY/X
dc5x1U06HqGEeQZtjOJBz1vJuVmQ0pL9lKeUlNVVEMDf/VH9wu0gm/sXWviwMOzM
pkH04mrOMHookp7uZdfv+x9GMA27moiEZn2KaH8dPtVmV+j2PclK5v3dTgWj2/q7
CjQy8fLmzF3GBcdDs/pjQy/GJ/GXCp8vRoHYWraHn6wk2PA/1tyapuMTI+Teed/D
K79MhAhaMKmTs90wiDs971IvRYNYgPITzsZrw6NJndtu0y/1jnievIks+9t1jXpg
Z0SKvxEu4NebTr3I7uzRa9Nu3b1B5uLJAx2LyIBQ+Qhrq/cn6k6acCjpfJ1iAeqi
SAjMWSePeZl6j9472J4KMG6cQ2ni0clHlDx4vd/kXdoyfkI5iZ+/k6kmloktqhcN
tm5uarq3nMLWSFUx7oy1VxjxJkami6vU+yb0rRWhjZWDwnY96tqccPYp1Zo1jfy8
tCDoly+x7w35Gn50Un6qvWsBSGegeksYxeCm2xOBKW/sjsulz/XCBVwshomMEST9
KjDqBqLGxohb/1FdnvboH9SwepUO9WW9wuSRGPbJt5p1u9rbwOEcsYvsSm0FffMC
qIiOpqlhKzKmN4ljxxK7MSCqALxJ7fTbwYO8jhHuqM99X2tAL1L5w4kfh+uvTWnI
3wRxvfmRU1Rrk6k0gkhskU3nXE73Y5awegDsU51dNlDTYMH8hlzK+/knYm1JpYoj
kyw+116V5dZESe3atVUJjcscW+VnP93ZtSNKNRuFYLQszmLosOi47hg86XpMEkLw
4rUBwcaHGV9ufZcSCVlVgyryRpPMxOs4DYqlY/XGYL0DHprnsRN/MIxOw5tzrnk5
zTpgPCfrzaWSNGnM69AvUV8YXVFNBTXkewtnSPrkLG6OIiO0xUuOUMwtreyVLAEa
wZD6sy1ZBZY1WLDJYpnuhkL9sFWJRKYQkCXzwpyAm+QA3pWvH4PIVyQ2vAn+YSzX
ARmUjtPTLEGtZBZnRH04z3iWEWmJ9uDgQKfNmkcsErDBRh+bpppv7GL15QsJ2c00
juFUoLZxOXCiRSfkCBWZWfZKL3KLrVdFavDt8b/VAKmjnas/Mt0EYD9n5DsxK7uB
+TnNqppA1SUJ7FiWahVNxatk0Bl+ugu5MzPTX4tjC2ku82C0VtGsE0uRLnOFRYc4
RxYx/T3zkIyLsQpXi/pSq4Sj31Tykw78S0Zw+nTFaGurXtzdz+RsqL3viTcYkFX4
0HB7wOxEAxGGfw96PRl/wQM/PBcQTb5KLwDoIbegcz7Em/1YwKBc8+xeAs5pKgk9
IS9Jdvluft2z+4Q32bRiAgqI6dkbM+NVHTRIzfQXQr5d0IcRBVJaLK0sxO7MmODq
yG9/EM364hHz6ZYDUF5SWdql5H6tWJbopKDAmzaGtzo9eWNyKbPGFWnaRTFuyHf3
Pn8+K5NxCjzp9d1xZhiYyb8+U5uih+7L1tJ2qpy0hnP7dx9r8MvpXtwqWtjuSDXt
OEo7WroQyOa6zzotvK/dkg==
`pragma protect end_protected
