`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tsWzR3YYYTxFn/3SS5fbHN8b4d9b059o7TWO6S6tR3aP9I8U8l7GsOA7HuouAaDl
Kzl7EjYvnfft4tkATKyh8VPzUHcPwswiETnUm4zU32PRuCROtdhiGp/URGa8qT8c
E0R993d2hqPzQUhqXQU3lOu1wCj9PToX3LeV0iq6owo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 48592)
Z3cRHahIMM/HW2RY0yO8cerYzzd2BvOX+DL84UybMoEeAcWxkEt9lUKVOAImrBeQ
RZlZrmHEOPNEDfb8PRGy9QoJj4GPgYEJcuAUmgVn0tj+nvuwsyMDx0lRmHmXW2Y+
Y8e0u8LePi6tX3BJTAXZ+9S1AnS8nTwSloS4N0tZKu/vLyF3IvRwqqxfBMiNCElQ
GqcyPmFfqVGJvv50JzU1r50T3cRg1/tivWM3wPiYKIWJ2dH13Ue27apbo5ooupwK
4C/cy/IqN7Pm5t383E3aLx+y3Q+F448LQmgB1YFHC06liAPO7DNmCBIRWku7xihO
0KZfxIAOHK0Gq3fyy5VDFg6raO3mTkW1uUnZVcGiJ6xdXXmpV5680vxPvbAY0R19
/KRRvpjh+gz4TTv0JeOgbt4enMGb4H8BC/HOc/cyBkpq7QxRBEeRlchf05HlewN5
WOFu/sliLvaVLVAMLbwLIQDYoKnBhDO1XEO2v6nLQGeXmATADBTs4cCDgYpZ/GmY
tnQKoqtpAIoA4Yxo6Xazz5teL5GbP4aetDPhUUl7pXbYqQolwsMja8JCtF0Al8wG
UnMPZCJeV4Y80iH/40jfkdInnI/wBKhm2cdoGs7EYS0PIKbNQXODTKwxMphnDo/c
ckt4a5hzpmYcYuvWWz4EQO3mlmhP6IrbZmU8mnuU7t6l2qP/yIN44dyxPUmp/UuY
iCa/tDHqGAWwFdU3WdS6hh1Vis9SNL+XwmbdmlGFbBjm7bgU1Istg8JBPodJcTWa
DXrJCLVIQjIN21BBwmSfK2e6Cl+GuZcsllB/Cj/IEAcYNHSvOKwnP9AjCMWvPWf1
dZv2sZ7rlz34u+3ftyaDVuxb6P9War8pQHZOZQTKamWR5+TlSyhmlUk7tYoDWlfx
cTMJGnGYEG8oenkquEQvbDwcjagSa3k8KOZapS3tyQ6zljLhqf7Lqtw5Nc6rHpvW
sGAGmRjx4JwMUlOYcrUytS7/FnZWB0DTKusTM8QKrSrJdj9IXBFJLztqGqU3wXuj
ADQDf9GphReLUXCBpjGkGfaDZ2Kw0bVqBYPkw4qQFIpr2BjCPGoIW8af6eAyHGRC
0VFkaXGEfb3aoYKrQRmYjhi61mmaBGJQQwcEZJQio7T/5N9FBpQ70WX52vmhA9qq
CWjEiSEPeeaTrUhdgz93QKZTEk7GkBw4BHVBQwqJUFIf/t2oaWDQ3eTI3I+qT0ni
/X7yyZBNS0IivjwBtnZzJ6uM9iW71ExZK4To1wJ0T68hfOyOlKsNO/5fc3i5Cf79
NpOoqotxfkZBJt533Y2maNqeifp/j1cnrRxZMa9fKNPoUMqPG89ALEQkLu8yhUOc
U0+xV6TWqlyyDTkkU+umoDMMowDq9eI3un7PDRvI5XmePW21keN2eZ6wvJfgyGya
kploiWpaifHpx/JgIkFqj+PLjP/bwHSHEg4P0cx8T8x7Gtf+arS4ndE1nnmXojtO
eEhmjCGgw54mZT2XR3ib8paLxeeOcBb3Sp+6JJGVOaT1GczVfGqgyOx77G4rW6pt
rCx7Fj5/T3ouJjrV40ZJwWuEFSvXph2vxoNL5BYbCXg2nF3tcpigepKfNFOwkktQ
lGEp7J+1rE4UeJWsTroxqxypABR9X1KrpEmxjkFfcN1aZeq3BcXJZIRz6d1E6fhs
yOzK1HNAuG3hvpPzg7JbNYieNiu5avktmbh/xzdRzhHMyZ1jstZ65TgrogpVauw4
RUTc/Ry2IGkuOJ3BLDqzpTAfehIK89UoN70CXvmqxufypb1zGyV5QhS8kfF5MfP3
MNSGmqkgkJrvglC7BDwImpjsL2wv+BB0F6AAB/qcn3n6y6CHIwTClQcv+bJlmqO0
Ime8VxAqNyQzv7jQKeQcDZwH/4ouGu0CsYuVen1RqfOV2qWrFM851K585qZMpYhK
fKlzPItAWZiMQhYjpMYRpRBPPibke0n1XUdsnqC+zg2kHlkaThZ8u/aShEZiVFFt
jREYO5Clv41iD3yyiQ1ZMjfq+TR8GDGrMhEDgUJbx1H9IY0rWSz96XqM6KaCstpT
W+LLPQltbCjte2hACIXCD3ONw95C2+BMnG1LlZhlVepcJ85O9gKsGSGK+DCMHgjc
cHGzr9cv063ZW+ZOwEQF0T7mBUJgH9TQENJ9GEkz7sNBNwyeJX0IkF2uzogYkQhB
NVJFMr5C9vo8XBf14aW0uuYQN13prFkboTaBGnRTlOmRwFcCt8LrT/EAFmv7VEb2
V3vmHqnWOUbqdh4vJt+/ru645q0TFux83fCBI27D2a6vstrZZtjjRTL2gquFSS8J
jX3gPP2SZ7kkyInUiAF97+bFmb6jjXERJJzQsqn9HS/1Ya1bhnWAp8wBCFrPZcbg
ZSFjgkXdv1kSPpmXE/Utm5dntOaLh/RinrXn7GvllQ2UonTovPp44yKZcDyrIgEI
JT55Vn44EhprZCtjgfp2UHHnUrRoo9RcFufd/j/Dv+Kqp06L5uzsxsuGYnBmPXhO
7xcXQciMiTMbsxte03qmlI6qC8kGKa+WppGVWZurjnq1OguMrPFKKZkH5+aqdJ1C
7shTvFTX4kLJ8P7KeMqAiyfXI8U65S8C3fH4t0JmPdQXXCiFoQWrRmL+ly8LLslo
7nZLgep7tONN7CDY+xOp734moVLt8SizWkF8VHPFFgyCizdpPgrdP9mC3QIKlD2r
pp4dMqxrI9KqIo3YxhuSYEhPAyYDSmkFE9ENpCz/WHiT9LnvGpvibYmFelDV6028
1vEYj+D3X/eSeAB8WggNdnJ931CrnVqdYyR9fKjz8gCEm6K4i/kHMhGxnayct3Hz
fNcuh+76bdiAe87LVT+8Dj0sR8EyBPJpW9tQDzP6TWaqtV2EdhAvs9Oo/21hUETf
I7eEV3fSMCRLa2+XueIyZY9loQkSWTcL0bfJE3j0YhiOnytuBgCx6vCGnAjDM7A1
l7ZMo6n1WRlziwGdI89bfoxFj8dcy9g+zNf0s/5xBVPKoi23ZIuO48WO+GaZAJY1
XQlCUiRxfj2vao8DS/nHck1oMBZByo71qpU9OLSX8ffOXTbTlI0R/mAWH/GCtf++
mYXdAqTR4BhdUo+gnGXRgnTNx581FaWl2+mqj+I0mex2LVp5dPjGPKOPUc6FhYdE
0401XBk+f1Ots3ft6oPVV4oh8Yx2Dk3ZOfnyL0zD2IKMt9uneirn57PCxobKGDBG
ZV3H7STJOqTOUkgG/a1ZoDTN7g/av3k6ABmFDBiEVFNptHTP1XBKNDxxnNshKYtO
fvUeIvjtCdWTg4DoSGeIcnUadYIx11uFytthUDBPV1/KUTnP84AoBQ7hoq9B2tBl
55MPsD58dDQ2+HieKoxowyAXpPWyiNTnK9bU4I3FWOP9qgIY0GyQZoKisakQxvEm
2M1t37onPBqKMKeuUQHyd9Y4iiHdC67EahibgTucdN6JJcPENiEcAnyVJU4WW94x
aFuML9g7JngOUZ3Pu0AcQGyaBFt7v/CuRiTr1WEfj8yPZzxwePWgLYAdDMWbL82m
OBqIoLqaU9WThu/mPKCgZ22euDLGoJEchN8cta7Z68Gz+rDX3PXbr14T2xncJ1Qr
K1w+d30movL2lnMFrpyEJI/iwC18mMR9RCZ3luo1//ItE4vHuDDof0wUSMMAu8SO
Iw951FdfRg681rhHmVY7zibG/YX7Ic8KJ8wRl+uf74qlAXrWQ9cCNjezmyDtFi8H
svfy9etN2joflXhhQUKfmv8BWrUQ8RTCquhd9Lr9yeEltXDBtzdotPcuZ+/+n4Oq
3RhB0/lnNf7M9ZRQjo6aIfhLsPRUDe3fVY4pzsMgPHCfLPg8Ywy10gNShqLnxBxZ
wx6nkyK4Dt5wHmIknJgeNUDTuN6+CMJqR45Hlra/yGC9kcwvMRI3Konlf/FBZXA3
A4WFbN08jQ/EdqogJxCbgTJO7JV28Uqmva9nnWvhhFDuMx7XhAPs4EWzLzCw8vQm
dYF9AIOHVtVi1ghdz0/QT92RgqCxEDF64M9uqbVn/SRRYFFcFPZKdqVM/A3usy9n
yqaq7WPerfVIXEboEqK2y1X6DAoavCmO0x6+0b0OzjS4bcroIeHCH59qk+cFoHth
NYvDG9hX1+eqZPL7FFQ1NjKc1hawQg1Xr04v+45OwPH2R2iXFFDL08UGzwb5OUXM
/2LAYWhedOc+xxlv5869mlMSFPDCWXlwR5UKajfy4zWBZ7OR/OXYyKhRNDf5MAJq
4AKPTsdPWrQbw7atq4wR+nOerZCY6k/Zz1P/SBTBRX/18icf/KvsljyJ0yAbqh2W
VnvZMQVze6mnXW5pQZFfnDXksyH5bWdG7IK/czT6hW9wftmCAW0+3hERvbB3Vo4J
0BTn3GhJXS6i3QrH6lwhhO9qX9snodkOGlyqFXiGWo+wdpxn5LWHhZpxKMHdaCik
i/c6JEHIfeXr9ghpcXAGr65kS7sq+p89Pqs+mFwC4+yMfnFqlaMwUGifSBRjZYU8
FN+IlSrMoljCczaV5jrr7WSLdvClVODy92WuEia2xmUsG3s2XOo6wO/XXPnzYQbJ
4bkgcQ6Ur0uTjsL7ThAV1jN3+eRv170GLxq1oKTWm4cQf2Ckbp1Ggr3PcrajB8du
NzEAa1r1HSmBc6xqrjUUkq3JT+LAu+pJbZUlYx52tT7i3sQnPltAaDnmzp9SWCmY
GvIrDv5wlItJFFp4eKdsTlV3B3l8SDaEE517CSGA7qFdS3dlebd+/yBKgJLkQg/G
oSwvGlOjnEF1bBZy5iqlUCo35M2IaGz41sLQO/G7IUgwVmITAJxEERU9+nY02cte
x/+nkZZ331NwSUECsMPsHrkcheQQ0OqN4gKvfJmkeKLnSpVtRiuF+nrnf1RPoUix
dHtKQRQsPJxw6rnwPeR7ieMc0KUOduc79yDlxGmLDLhm8Htc+YIMGJUKDwsWNEr5
gG0ePcmBqokaL3JO1qly74zQjt6R6DT2btIRrlXns7ToDuiHGkEG7qPn4vs0Wfwc
NtQzQxE6XubRNRCtwUlAbCVtvgDrsR/NzWTARNBKI4jGHDl7QTeQPhoOJJklyBfE
o7Z/n/zGQSZlJJdwb1XKi/i3XKeukLXf+x304WFCerEWxEVtGM3V277fMDgZQLm5
0kjSXHAB0nG7Bp+SM8v/YlQTnnKspTFCbZGkCJfpJ2XGcGZBcpSH8VD9EJGZb59E
H4LKkbolcVihBYpgvpYN45nWhv3y0R0UPZIEIEj9s346fqtyj6lqh9kh+rXEJ/o2
KZTUjNANsXe8QcWxIa1jpK6QU36rSN86GPELxhPbo3Efph+WtwvFdthFO+wqpcvK
g8jzLOqR0ayWhr4NcdO/jgt6BgUS1cNIYvGO6USH6d7DNz6tIM6I0yfsAjGt8ZEq
gMjPKnak1Kov6mPsgWczoR+p8MFPm1TS9dPZvVM0zJ7J7q17EqNAzYKyEe0NG3xh
hxyMokJu9G9pssD81BXr1DmzlZRJUlIKq/Nzjx4xTa0/Fth7s9qEzqbYONTB6ARH
I6QZgdg741if60J6ZbgyTOyHOSMFLOgw/tncZ8iGCGmpj7Mf7Q0Ng6+DcTeG3OT0
6hhYll9GXND1A76WznZDE7zJTbkaFqrmLzz4zOqbZh1gy+SzqIQgQvdd7PSDXnIO
B5PpfeSgn1esbxyiHcTJ4dY0Bo1aH2ijip56ZVQQrbbLq4AAnHaSHsM/qN/TuSyh
24deSI3DiMpm4TmsH6XLYrlaQZXyTmsx79BVCBsEPeT2xLmudskCCbaNAnF4pJqq
6DhxDHjFxhvf0cQxBdwjIX7ekRU/HavJDCzslaz0P5HVqJYEzu/WLil2PH8+l2YG
sq4c2oZbyXi1957hPO6aFoCSQKcdfkCHHUqy7hSrCRfEPOHBtlFAV8DJOj1+9XoF
VDioJuipq1xlopvqzfPGsI3FZN7sEQ2/kLeSXXuTfWI8eucwNaTHm/29QNn9iyy1
Jv0hActj9sgbD/eAXE1HktWbyXcOJhQIJ0JNgnMOcOCV2D0ml2E45dGm+y1AkQqU
eobql94S5FhX/XB3ezVfAkc3StGg63K4XWNPJA/e/7hfUNIfhmQ8FJ9l8xWL3lgi
UhsvsFbNAl9sQEfBYZwwMEmZ4dW9aBCh6QOkBtobNJgQu/3TLBK9SyjYlefLOPL+
99CmPunAxDA2n5F+kKajYnXuaXIcUXuVTeMjqaGpeE2d+iM/cyNJS2DNvXAzZyCk
ZzFzW6Zo56CkAXOZzbRe4+tdHqDOJVsLcWjgRhWkc3zQmjMeM9czFG07qqYwrZ3n
SBw4Z0M/QcfC4+EtkbnxLr3GPMKVdTnyLPUtPvAq/rtvJ7Ooc7mJ7atvUJ3j2mWO
RWUl79/gUUbg8kk8CTKUvFpOb6yZEZ5kt9GpKBDqIRBjYWNL8enTdt6NQGPW+bpY
L/flFB1nFDZhUMroniehJ3j5jUMF8KzqoBO5u2EQcWwQiBrc/OxtmrHCDpx1uJZS
I7XUUgQw/wnHm/oQhbA5XmRoyHUIAC002AY91o6GJLzScPD09nD6z5+pPI43qRCp
JhnWQQHzWJvFgoEetBaOqLz56kq1JhaUOpl7+E814MmcFgsvWp6zsjqkK+gHVz12
BPPD4Zevpx2D0pMjTh7DAbcrIfb7h/csqmOcvr5IaoFhWPbfRre+0LIeTEum6rWX
ybIc0VU0mvmXxJjN5EkL5xyZ4tgN9wgM2uwQd0BYqPTzTifN4Gf2DOuhb1jS+t8z
NEJu6ISjNke+pvH6ZgRjznHt5evR7PTZn46/UTyeXkoKFEZUzAOSLT3KaYAxU/Q1
r4CbEgrXYJIBnpyT2YzmaaniDIU82e+oHTajEhiE5ZlLHJSvjSXg2cFSAo6o8cAO
LmsEpc54SE8je4ll9ZYZPhKaMeHQVYiWLQtdJ3aKDaFaG5dogWfET51Ecfw7It8B
NHLAhjUy0KWJtUASmLdkhUUCyJqQuh25ZJxOPgnJh2CdeIXh5f/rwKQAkdQLLhem
Aliod6/U3Ah5Tgum3mH7angq6StGLk7Xl/ff0/nFFpCu+TDj+f7zsSc8KDO7I6mI
8AoD/jFYiAjraD6nUZLD3gRX9iGItaAud6e90y/WYcqKjV+f5ZyFjtD+ZFf2aERB
/Rp2ZlqkLtOOVpuHFHI77U8HbP1Tg3Cz11Y+J4DnJlwJMmQFUuogyAogK4QGp98M
bWuSoqziikC6YNfY6qMSkKtz/LoXeyWmZDIcZZ0/DyCrE39VKWNFYrYMOgmrp9XM
lomVFi+HFcGL3axm3+bDmbgvy5+qX3ccnd7hsWqYO+6f5R92VEnAegby7HlJpnj3
+Ffa8MYGUuiLt6PDpu+Di6g7ehr2H265GpwZYz0bbSF/BXBL7HNDCapTwISPRy/E
loJJQJEEKPJNnD1Z5sre8YQuHLzy9VLl49MiagnJeoPgIugc1wSuOiDby7bAIqiB
AgZmUwZz9mUGp1cXMuk+rTiFY4e/pw35+FMfc1aJpoJi/4rY6nrN1lfvuxPHMKCm
7p0SeWUwnvSiPNFlY8trkG2MWBEy4cbb5mPEa46Ep6zRWl7YIeqeiFzxW+wxLH9c
RnbMaudgHFDmPXTUIXL3VVknQdFf1xwEO9QAfD1ht40OmOHg9BWBnJXXWN3p3nNB
PgkfvHTmTr1qCs09A4EKAtGfVzgbuzhuML8k640lbGxocr3Z4Lo1Pssv30Gzj0Pg
thADZF86OaGM6S/iqFO+bsJlDqezuwZ+C6SdsaxDK0+ZVC8m9y8m4ZQ4QaeyQxS4
t8l+UghNCm7qa+ofmuzB70qvcll/kKM+3DOc9OxT1zE16zFyLWXKrAAW+ah7Hvnz
zlHGwvU54SDMGQpgl4z+CKqmgW8VWZBX5mbPYUe6aaTXU+zw3TYtw1Gam2+8a/7T
HnlG0zsTYVHgMk3U8wbBjsWGKTh8uFmJYZcXYFI0bziozNfv9xxTLo2ZPFWN2BUF
3XKhpa7zG27jrL/zyy+Hi8xu8na9Yq5PKk2UDjOnCfhauitF+tOOVTQZS+QwOIeQ
erzTjDuuSJp5t1mULj28cOhGSfVp21WuwhXnb2acnYBSbKxwfqXk53FrCJQXMCWE
XM4oMYco1zg0noFvwCFs7Ig7gfr6vx6Hm8RMutosS9C9Wsalbn6Lne9zCRozMpnW
NZ6/QZT87m7uqlAWrHTliU9nsR2gHGp2/krKhl8CXx6Mw++YtOWT8HrPza0sCdCn
AdYA2y4MSC3Iy85tM6dUsyatZ2wbavxMURwdCzIGsrQ7J7BL4iRhnAqMLgOUmPSX
GnctG2SxAnggsQommfsGz9CIHh+EOLe4UTzTvMIJ4dH0Qgh6JcHIRroofG0qXT7o
j16ytTpBa8Ph28a2rIlvOJ/hU7vdklb1VAif2kn2hVV+PFAJl4sZx9QVjfFdCc9J
RzbItUL9iil1YGKIxMBXiiowiKw5d4vuOaq2SlzLk6rd6XIeTCvAFmk0N4ShqhYx
hXEaGfPxyLUO7kNgZI6FKiIwjeoLpw5rwNT9LhJWyzIrdljh+9lGoCrBfNQAwdIW
/ss3XZ8Y64CjgF5R0WY/BldyaEHocj/POsqXJ/lX8KBArUKzOpqwWxvEJes5IpZU
B8SzklJsEj/YtWla9jPPuLHzSwCzbEqpWT4XMuCdXl9yNKnjmt2jUTLEJ2mnRK7a
D4V6kWjY2099Km7iaLwSTFaa4J47KVqhRIGiynReN6dQFK4w7VW9ORR3w2k9Lwmx
p7Hiv3kAkgW5nReDKlv14pVdiEckPPn0JnCIpTtC52jhfmWWDt/zA3tzn9cG7Zo3
d8uvwfOIWROsPu5rq7NDu+d/A9to1b8QSKxXsL1qlKwro2T81UfcC0FbV+grkU+p
zISOlIE7mKGtY1bUsgmC/RpK91WbyYRYZeQgXFLnlFAJN0CkRYYUX/0U0LC1/Nr4
dKM9H/d7VtXjnrk+/25MolYOCq+EAm1A98UmxbWXC/c03181ERShEjE2RbQGrxfV
gikJeoVDMEGHi8v9wrfQBMSGvWLKOAal2Ki3xvH44Q5nhA+CXbYdwhTpWg1iG6nG
EP/pBamVA+fKkWKD4vimHYM4+xSZ0kH4HtK0DnzvJcU+Ez3fyaLu3aDqXC6rgC+3
v4PdLBmMkZC37PeMj1kWT7rSB7NFaZY+TfwOM1MlOJoYgM+PbmDN4oslHRIcXj4n
+1olpYxglh65B/afMTGMTUTf0V2NFTG+jW7PjrjyBo9KhXnYqcyv2U+5kMqnpjSc
4+COt3NOKvOU/qsDiiE4pbjq3VDKRK8yyxlukQ4qilESQJzlt1hV/SUlJXjkgWjf
T7DDOsBF9rDAyI7EdW27TQV3bx5chNBlZy/+pT9k46pLXnGnQQssyMm96UQWbSsZ
AN8XZL4YzsrEHvJDbBLQ7ItbteoeiSEMtc+opZMHWe/+sWNQjefuyU1pe8LMK3Po
nPYGnYnqcH5sTPzA+6mhalu9Qb+q4tK1IEmA/sUk3FkqdwG/ueCmY06adUbN8C4y
0ZSwW+/62gD1xl730uTQC0XpjUBK8hSYJ2GWwPHoHy8Aa5onvPQhxYovA0+dF35S
saAZb8rd62Bhto/aSPbiBDvDypWkOu8+Ok7q9jqVjXGtyfaqCk0y3TcRWbtuamhD
WB/hbfizrYNlSItXblsvmmCDZAbn/CXpcqyhEj5udUUhAumEe00piTpl9gGy0YMU
9JV02Ac/Ulb//R0IdKogCK9n0WdzwScC/iOExJcPkfvUSI3A32zVkJwrINNoTmvO
UOl0h0ClRa5ysHnV5hTPAqkbRDysPU+Yjx/6Y8+w6M4ZTcUja5NiS++j/d/+U3pY
uzUwkFkuWoG0Hjm1MOpbkmu7L7l5yz0Vxmfxe7sxLFCPsQU3ELtYP4EsF2H88RH3
pt09iXgE6LW2PDvSqs3YHTVTsC8+8eU+EnZvEvW3uOd1IF2ibEPHw/XY2rPDbEax
LTKz2+jYWtd0QI1+otAyvkpUIRh+xTSzGb/WYSkcV/WNZQz8BsFi9hkdF6S16uxJ
QaUbj9kU1l4hcv4cVrvkx8C218xJ7kRrKtud+xpzX0HEmzviMqSWvT1n7mSPnJ3G
81q1dijq9zOXnY62ZV4hkZTVNtr7CVtFyZmjilwSVGM77kLttf42HlA2B9ao6+0s
t9YY6GK2J2swvVidaVpi5YNsGheykYlbr8rLo5DAnfMHUbmvjWddsAdQjWpeTkGq
4Vdq3TcnqhdOAPoKSqPsl339gblCobI92QVPrfzFRRUq9s91cJ0YgBuT5Kpb66/u
EFCdI1jfPA0bOwz+aPg08pK1N15/a4gKoOAwA4aS0RflcgIoNJZZ0qIpjsR6lZem
5KbbEs1sK/4DYDS7GWa9CSq+8X3UP+0RXc4IF0Pk/NQvaDieUGFuW/2bVTQolbV8
hx1pa4FT4AsTx48846dxuj41EGfyh0890IS6t6VqjDUqVk47EYRvFb+kutyLGn8p
JQESfJrW4CVjjoZ5u/tfHqmGJ3WhBemnHXNn6/GE+JSjnU1g3J7OzStAkytQHvmS
WVXLmcpIeIGtPLZcoqJhIniXV4KcOYAuv2PXoxxmh73QV0ZxgrxYDvQd50Elulql
84DkLDRr7Lp7wJMwrp4zoenSCr8fFIA5F7lqcX7nWc6JwMYdt1mP7w0Yyc+rRMi8
r2dIyXu8sPPuVcAynqT0ITxowLGCqMcGMdS1bKFVBX7AtwtdM2dxGbzfWoSIpkJy
ioWZNRnh6jwXomAvSyggMlJv/P4wVvH/mhti/Ln4AQlQQXUHPGV7MKZ+hEmSftmh
+tRoMXukiHsdvtQjKIVi8sDI/tguPtKO+fenOv3FH9OVuI+SXeHOkM9WtcJExoYo
6+4nOwXBDmgxFywHA/Q1asFtzzYZ7ZRUDm25wCkQr30SpT+G9EUOxH7FL+FLZXoI
HRaFn92Lu42pHr3l0/rQyW0lhngD7gt4T5KfRoSVqSDIxE53MnsD6aK2+yk6pT0e
vPQmTzHS/moXn7Unj0i6ODvKxc+ITXXuot/uuCmi69Q9o1JtRCxdftnJP997lVlk
9KaigcqYRUQaqKbSP4Nmikt+4FXF1BbBTdibIiSRCxAI44SJxSv7Q22UqndZaQlp
6IzSZLlwE8yHtnWRvEG9sMoIu8A/5E9GAq33Pt8tfxTTKTbiLqOu/k4lTqb1/Q6D
LYoAFtnOzUZC6KIP5hdJAsq790gmBjT5BWYfoUfzUopbn7JjIzMgB6biyPe6h00f
ds/W6GZMHn5VVBiL5zNxIUyO7107iNYq/Ho+9R8n+ELSIs1XcoTlt3dZdKUjbuhH
12q3giCp/Hmom0vOEFO7zwjxFpx8Fqu79+KrnuSSvjer27jjCED/FLbfsFYZQU3B
4o1i4sYeakcuxITP1+wRciEI7XXUQ4S16j+LZDy4P6yJHFpPS/V7Tyz7BVncsXd5
FjbPFXOyo6aLPeVOVK0ztYiBQ/WmWlX4ppTF4d7tOQK21c5wiH/wEiaEi1t1hZm7
OpR+00/lzMA1+jAvbFMYVonLRAzWm3GLBA2+/pYGG5ERfffDsNkXYyrPmU4OCOPZ
rawJ2d8gEVQmVF4gA64CI//9q56lHjBEMGJR4UF//ZfHZaTE+0XOvfRJDiIkCGRJ
BGd7qIB1v2i0KHzNzX+5mr56djBq6rlmFzhJTAvH3VcIu0CI8ltuXeEqqZNbsBu5
/nEo1AIaWk9J+w6bDofIPDas3uFSE6cpdaG1vjloD6LqhJZLq0KJ3+amVLRdYTee
VycvL6yMdqZJSFH+GapMHdzhiiDx4KlSZEJn1UpxUFnZ4jfwXZETci5BuUSMbaxv
tO/2uc3tJjHKvK2buT86jyhd6KO5nDxVVxWfQCFeZ2f2kX10e3WWL7U5Ua/zxZ6f
Vyk+PavBIhFPeCO0y92eSmpsjPkycM8fD7YBJdb3744LvEuk72+Z5j/tvskyZrSR
qo6Fe9q2tVZyQzhEg4te49PQ166QcHWLVENTo3u4EXOz73K7/9nievRmO12cVlWE
86jNVSR/f700dwNTAAQAI4ig5gguG2kpwbx6VkI4YzPQkYyR+NTMxxDcYjw1CANP
i7x9Q8Um9faCTtFdU9QLXSoHJjw0QyIGGbQcevAZ64jW4eLK2DYE2n5j5+tN9Hip
e8BfuR6CzwwKSdXbxg0rEgAdl6AO4erCfj6C8K1toa6ch942p2Dk8j6LxppYJkxp
ulEPxq6rS9kXVI591wSRvAsjMUkVtXGKprKUpkZ+OSmwceWIfNqtUG0lrsF6h655
BD3mGkuaTMXmXmvgmGggLly5Xp8p8bab5F6q8kMQ1+FYcE51FGwADe8PtI7Zt9Yh
3v0s+KzR0ULP6TIEObs+tlhuAJlMCY1O/ovLLDfs5VfPYVgJcr0pJDTBPfA/rbGF
VlZQ5B4yTWARr7+2nvmkzGmEOvh83q/INSbTHQ7CvFyCVloPc2yXv8k7VXqyyi61
+mb9l4hqhcep7MIVccN1TMj5ge/J9OBFsoWtJM6cCRgMY2VbkjYgAX9VGogQpoWu
qaKL9ZegatnlivSgWIr3dXF+59e5/qIzoVTqyiIovp6KLcUJsBsKtNiP2s8GG2Xf
W+9KvNa3KmRHdQsImCvV7/1/Qx6KDoPPfffO8KKpxbDYlwlRS3RoFoewFOW5v+Ad
jq3/5+GRRFo1LoRyxZe8DPB9mp1ko9KRjNai3BV8HRv/sRRqvsnxfkujLXWdaIU6
cI/qtW5BLvbZNEfrDt8Yr8QqW84liRcj3ko5JfToVtHq2Ukve9SgCWR4e+Vo28h5
GqW8fWcTFR0KfqfsrkQhs43asB9Gn5TAIQjHI4no8yK6JBKoNFSScTGOWEqunYCr
GzZ5XmqXoz9poKLM78s7aK/ebvWZn+0RI74o1A9btjxk28Bvfjp4bxufYbzogjpd
s12YqoiLoW7KQba4szQ8rtNvdmbwAraudMJ7aIcfb/tuWETOsQ9j5uvqaDsU2K8j
NQriG1UcdYjV/vbZYoFQsA+8QI2+5LrP35vie2EjjvqGiR/1la2HxXWg7izQ9/I3
wALnENJue0pUc6l/uMCcD1EBviIzYVeJzgq6h9OSmXyrO3cSSjtaE38qpi37EWh+
5QCQrkH2mCwLIMwJvI9K1xFpUTdyvl7gRlRty0T1LxAe732yaBrhHIX219bO+nka
BZcPOOdR1egXRaQbW/Ajpj94bEYMTvjgUwBDAx65wbDsLJcvkkM8rqTBnC0avJDf
pS6b78jWIFzFTTvnTkoQRzo01oYlbDHsR/SOdTfX+S4gff5CqWI4X74jq0duorE2
hP6Iu08Ea1J+1VXCY1kAkRLWkB4gPx9iK6j5en5FWSE4wF+dvks+i+rq2AhZMs7N
cpTfD+TsyiXodZmi9TielbfsxQ+B+r3gRgMdaNIAA0aMPBvNR71v7xUo0U/z6v7n
di8kawzWtgUXOn3papK3P/154dZazcE9LVPPolKCzqlmW3kh9CwtUpJMhRpH/y+T
1Yl8bYYE/Tz2V1LTbtPkj76pIDvWRXB4OiycMVtWwq82BZW1dPViuso/EwMvsQDk
GTDknpkiOMlfaD/sTEG48hhKSxnLWSfa53XvkbuRCDjUL4QcNF1Y6L+fYVQwFlC7
9IcIOFjJ6KV+o+ig7q/G5CGdPBTLXtd+mOGbJJfQ4mtvfAM6TUDCc84pER2I9dn3
zBogYLbRDuVkVbYADCmhVF/TMVA7pmMIAqZVTy+NXwV8Tywv2LcS8yLxJLzTIY6D
zSKwuTKddvxF06dlsd9oeiJ0W+lGtICk+GktsTWlw96Tx5jXUhWQ5TRdqEHExMLc
0eTCxGCf9+pR5z1KdsgTzFYaUteojS6unyBSK1aqM3kFqdKjYOSzBCh0o7qvGHT6
nEVuIb4nqBVRPR11u5acyiWWwJJULr3Xl8qSeM5p5YaYCCXy6/sKqQ4+Fwd+1tjR
/5/xug/L++tocTUAWs1aO8rz1lEnIJnpIve2dQF975T/ea/4mQdJBpT7UWFHOTWL
+8/uLY5d1PJv8K9bzGqgl/iukzsh8l/mfe6GITytH6fdL7KWeCBgMOGxjT6D/c+z
qvusiUiP4RWyYfIEoguLvFa+deO57Achx6s6NkfyVjDqTkDKvEnPKZQClEOY8sDy
TCjPCoo3BJmKdQn0S8dlhiiKKwdt6a1VB3At9EbxF/KTwT2ZWMEZMkAIkXy3pXFu
mjzulf6b5ZMCxJMR00W6rXcPSF5FBGamDs3b3Odba/NxzqE+AZz/BOjRGn0Z8QT8
NSiUfUfI9eFgSKPp2z59Bt/nPVaecABLGVa64drUJmcaMy+JgOu2kbmJa0nijImz
YqeKJlnv4GnsRdFzUopaTvtRXTtggk2592FnC7LjlBkT1X+EG2RRv6Nuqatw3h6g
iXI5OqKCoT/IGLTZhBDn/PKCB9vGF9dmh7NvI4mnmuLUQ2CRTkYhi+IjGn0esQFq
7U0SvLLKQcLPE6SXBsDpbdM06t4/XJgfZ9W69OMrB0ngdDFSHlAK3X1E0nZ0QBJj
zoKXUMIRthqYZQsvFvrPu0UjKJlJ/bZUFr9kPUHN5tGJ36liNzuUEcWpieJSLFMQ
HU+oJMEfAC42I0zKm4J2VREU1WNVFoKVulVL3v7GIxVRv5cRmtHkTcMvSnCrrtG5
SwPveoU7Utc2QZL4v8z+OZxsJSYAvZF1VPbdxTKJiwqq5btYnsjnG0Q6EyHWuYUo
sbvcPgqtR+MnCUtXVtA6LwzgRH5F7eMXu2KET4Mjc5p8oEY883cEwLZITFSraahX
FKRhPPF8u5qwbvSBbGB8YQjhDAxTOi+HpoPIOcq1YRYmAKaB+rZzMWrTab+9c2xY
X96Hg/NVNYUImiVJnouFtmG/AAqJSYuNQja2KCVOpc1t797zqWMBzmMusJKv8rlU
TFm+SdrOn1QC4J4TBFOs04HApvVr86i9hoO7lObqKRKGxS8M5bd/uOcL1Omw0wjP
FP1+Hhm+c0Ldo7+SWJIjbR6P7Im2Mrea+RvbVsgS6l8qgEBtZeMHXENSRCgOs0p9
3Vygz5z5iAbkEULUocZ//DmkSACQL3WvHhSLEgMmN9e28kcl/0hSqPChUiqzxqEw
WbR6Ov7bSkdpwuIBiSPP3xA9Z/Sxjjxvd8BqguosNohuMfS+bYSRAJXoeQc38g0x
UfqPpE60zyeiQ/7sVeFJNYtqzIywgalh7KnNSyA2YJLildfZNZc2Bx3MarQmW6so
4McMQCLClTHWFwmCdW2JN612Op5GeDnTkjZeBLEmTnpQIiTcN7NdBhj9T5HsGe+4
XUM180ZF89374clu+babjirk9CpURDaH9WFfZZqbbVfBh2vtgYlpJ3fi5PZAashb
zNAdgzCOZYuUHlZ8kJgikUWGIVcWwgBR9cstO6YzMDliIMttVBhNdomoZvR7He+T
C++NbEhewhdrUDteSCVSNNuTStTH/HXpxlQnT4F4qqD9NyYUFxqRYiMSp/3ebiIg
10cb5HFPJ5G72O3mim6j7nB4rBiKDNbhYdYGLT633xfo0FN1o0akKsM+x/QwGW8A
HnWRh8DuejlI41q+JD6CEuJwASZ8E8l5bGfMgrAvW2OpiL98LYubHSAO2NQD+j+U
rpffqR0qspWHB1j5HOd+DF3pBPr9OWKY3u/WACXvCzNPYvESXoXqZFIdSgigtlXO
sEeGZqny3zEkTEAxwct6HjjA4K9wfsrAdnvz85dwk/skzLOHswwF9oAwmrNVg+tC
L0f276bJ6Q+5095gnTDRAOTAee+byE9hoKNtrMDBZacRKonKGSKd4Gc1C6pMmeql
HuLJK400HyjJ4tJMLqf7g9DvvDDuwDxnaj6qNJtsdV89qxMo2E8s9yg1dLBR5JbE
X/2ODHd2ODvcjcbAsCXCSyz7Og4YIP1kPXXs5HCpy3B2RJFoHRQdRHvg9QSo0b9q
hkYqOqGv9hi6bszBJFcF2/P2xBypoVCsAm8XjmSqfSf7bwzqdkgHVhwftUICfVLq
utmfqhA3y3C/7q6jjaaiGOyhihJ4lXfIKorIT1CfBxHJOQMC3+CSUJ6BFYYuYeub
K+iJNScxx5RyvkUeWlzxexA4Ixn5zHODpwWTN24EhLBywiZn+5Xo9taCvXbcz+uP
CWbU86CnA9tIu7IxVJaybbDZgAiB31M/avusBGi6YEpr4kfnQlPhcBZpPvwTN/pW
qwv+HXLr+FtGQdJl5/M/fvAZNQJTMiwbjD4nPE0PIK+fwLZFTeYvo/jQbcfuD4/e
mwEKZl2hQSJKntk4jIfTtYkBnhcel3Fw9/+glDjIqVw4AH7hG/bTfE3eWrqOWI0g
EjouugYvfPsCJyiplbaC05l3H5BL4Ru5O04jVSkNNfHclwxqm9JHqfz9mK0HBEW0
x8pxSeeoipjXx7EFH5ZMby+Xg2jOC+EE0mIFu11KX3YenNcxc0jIR6Uwe5MtNNyt
sGcrQszpZDtw75fWjhDdvbWIHYIWfELrw5o/f1z9N/lU0MFY0UO+QCB0QC6dnHA2
gPrFayom3QnDCRPnF5080/Y3YM9pbqltCnpSc1d1rmWk+keMuAgtrsplqP+3YCtT
H6rz3E2bWEMweffrRszOVPDOtefI9QvdqgvGrrTJugRvUh+X2q2bjgBxJvYQnD69
jBznWGM4zi/KfVc/p6u+hDZUA9b8OqqsDT+thuQfl5d3Dfgh3xuMCLQ4TTwbxcrg
MUJygf0tZSs5F4xsWSZaAPCD3/sqw1xHtNiwhCbFkJBPZjlvOfxMmv/3tgx3zmHz
sUCnuMxvRTjq1cJDebNxnlmWqppOwJAv67VQmupPqfi0gh++OgqmMc7B6UUAQCdE
sbiZ4Jda9hhZVVsdMKbsXY36BuPGCQ5FC0BTe93yDD2kXSLDmf5ReuUDLMUpojXU
MXK4vQNZAB+iKDvsVkVj1jW5yxvN3IQJb9gz2XaNgTViEJgo6AySjT8Vgr0KO1+s
aTc25sv1duf6Wg2+aPNDx37c5dp4RWMrwiP9SjnVtA/FS0aEHQcraExdn65MJPKy
LgUHcU09EYJRMvwHDYaOnOVCLTnUKXLMJ4MQiyNGG+Q7nWapVzwbxukjbY31nC1f
bbeSFK/IJmM8SupZqAqUvJ/wcaYrv1BzMOJSwGjTNOGQSC6Fp2BL3iZ5eLcS1xwA
i1CEQd7XIz8OGR7gFdjsvWeS9+79++RgGQUrx/3Wfo7+qrMv/3lOwIoEmg2HbrhG
zisHEAUZgD0AHpXH9PLNfwFN7Br7VBlyQ4mEseElzeUgbGrkHziYrXAvT5QHp0Br
ugnMe0oMR5DpeT5AISdGNwFfCPsYiQpcSVa+DhyeOcGzZYJ1tw/6tUAJo19BBuVL
k1UKLZAg1klLTDflsfoppzhV91AuNFFxHUrd2+v/vEAn0DrUILtvl8G9eErR51cp
bDDFYXswvU96AiC62FQZAR8o6fsdKSQDVsk5joWFrmnxh0TfUfjGKowA2ye3RmRt
Sr+rNFxhd9QjF2aOhugzfcED09w2bIP6xMNZFKpsvTjtcNE7sSDZ/EpQnt9vU/k0
FMlDEPy6p8qv/+Co+1trdedVm1doUnaguazx8XQlLyeBP5oa2Kcu1SQ6V+Yr+wz+
ZcpzbLI5T61kpRaCddq9Z4x6hlXiC9Ukz37rdcQZPnkyZp59nIFQEcOfhjhvvJ5X
L7AtRjcf0pR4tpA74mb72KK6Lwxc10SrDJQYQp5O3LUQT9A9XMqJSsK44vno+CC0
KTOVGxAMRcC/Crccfe3ID+BcrvfVFI+egcudP4pwhNUwLDdfZ9dx6QvQM8wcomg0
TbVr2Arv/dbt18ZyDf+fLS7xX3Js41D351F7FfMPkfTkctXaiuuA3d1XB1vDongM
W/pDElfGlUfnMjxQJGMjU0g6xu/PZT9mwZQSON/eFfUBJqMjz36QUtxpgAWD3N2q
9FnL1dOIdEAeLvyE+KRqzeeGFZlOu1Yq+FtS7pnkj3XMPjCJ6m28JJt2X4GcDG0z
/yaAYTPJa6VCVo6KmkE/X/V1qb/50PZztt4RxEZuMVscrmj2+doFox+RQ8Xpi684
WmI/ynYv7ezN3QxWpvoEPAsa+JWXEXJLgfL0U6eb/7MuvD994J10c5QdtizfdXqp
abmcvzBr5WP7eqM+o3vffW+7iJMCguYnD0x9nPMqVebVSRzZf4COmLaD5qYzzc3r
2076gZsKlHKJE5wwHVp6XSiFn2P5/jE2QG4iyl2oztgFBjpthCc6jQdcsBiDDGlh
O/BE5X6fwXQwOG8GjHHiGnPM+1ocwADB7a95zXAKmv7it4Mu3i0WT0Kp6ISOH0OE
HXvKtaD4NOK1Ryo+XComVaWGliBeAXCtAa2a0iLCwNr+1TyGekKk5kH9LBrCaEWI
VDkbwazQnebK8SC0oTTzzEopsoJtpgbA5j6Gpaa4/qzGOkD7eqzWSNvLdTjtwx0s
2Mtbv0h78740BtzkUjAt66vqEzW3QgSVGl6jSNBV6OuAhhScfniTV7lYW68uw+k1
sKqO4FPufGAjkYyJT3ZIi0vOVRZAAsLPlwK7hS+LIed3jTbDLxAecHiVPEUasX6Y
7tLxDFnUmhwXwuVHDZB8WjBxFucS7NfF6tkkwOZA3zD1WrY71x3tGePqIYWVM3vy
Kcf3sJxauDXs9z0vXjWuNgHWCOZEvcRgFZTZP0aOJlS7SI3UFGIP864nxnqiRQm3
L2W3SRkCFx1KkOsOPulI4bMDjLgOowePATOohtEe4V+ay4CqCQ6/DAw47Hmlf/f8
BPBdIcFJu3D3bqoaLR6cccRTiy4aLSK7R5YhQOZ+h20ojsezYGOmwg/AsGvlRsvO
KNYa5nbIrina7RV6ZAJfJPldMl+zp9/UIKUKPL/m6ZUBddn4QZIb77B/44UiDrg/
7hh3kkekc5mJgXXi0N+9+6+BXGZU8NG4DrN7dEFvpstB5Jodtd3KZ7OsNHEjFfjM
PIO4VuBGPNjldcyZqT9a3KSfYc8D0PTPnZH9r08g5Z9q+W1wxxgvaCIRuCfMwmui
nkMvSSURzmqkQ6M5rVP/IdynQt9ae5tfTUIeMwqn8MQZ3ZrsNNM2hLO9pAFcRj7A
3dtMXVjm7b91AC5xjRQejJuOHOQ9XH8KrfWuBnKXCJjU2R9M4k7jqkuZ15V9xzMO
d2V2Z7+seaohzj9vjI8PPk+o87kIKD4D9RAiLdA5Pjv6pSxttp9GUL95SifgDH4I
p0Gag4IZD3aWT588rkGTlz5MsgKhrUd7mDm7te4oMcrCg0YlAl8/lhWg2qMzbPNl
9aUps0+Fueb9N+hwWanqkC8vG6fzu40DwBJxZqyNxJ4TSpKeFmGS9WFHHOWPG2hi
nS9oFEk7ocFGZum+euD/Iuaiu4rZiro6GAFgjCbrcfK1goqiCNvzBcWx2NLALmGo
EjXpPsxRr1ZqKOYEnhP6/+Y8S+V9zCg+DojYTxFgZNWW12S0vbsE3VhtMzoGczl0
2x9OIUKAzEav2DBGiQK8vTpl3zMjgWkNL6zMRrQnVhJVNxf9a9V/T9mpQvHV7aSL
U5CoJRraIrHdypcKgbgOF0L4owEWmqwqMYTSZN55aM3iJ8BeMdRiYl/+HRbqhwT2
DAUMCR4T2RMqidEnPmsHnc48SEcoTo6sgKgm9Mk6GEdZk45eQuHC9hAAZGL9teNf
sltvVTlPSsrO0BuPBldcCCWAhgEzLQnPHVI+27nwsvKrQ5RGvpD+P57OKOz39egv
65VbKAwcdjyBg7DVjlKnM2OqsmIpIAVwvrVLyy1fPjpluQxjpMf7uvnK0Sua19sy
yKiZXpHhjpW75ApxTCw+8pFgaSHxndENXU9jhXmliQDliBcU6lUF2+UVE+VAEddW
ooO5BBvYJ0svI7VqrZ1iJazZSaFUIALLgB/nOB3OT/77r/V0U9kRVNyzC+OHTjhO
2vRiCtu2e0dBMn5saqCj6utt8rD0ysl2lj5D7NFCgcsJLJb9kf9iIswLt1ZKUPOO
34t8HBXAp8qIPmrT45b5ScbHzY2lrTIRVr0TXNqEsBVIaui7MgV9KCfkHdFUjX0B
Nzjza8DHjsrA8/bZSG70Li1INMG3BjcsBj51EcMhrHrm4w+q1uJGOz6lclOv8vhs
edx8VC0ol5LHvSyFCvKfRsgy1TQl90p6pfB1iVUxAwazEDm3bMzUzMh+iQwZbrqy
E6NtgnQ/sFeoxxZIHewjmnq1Nh/aNZylOMUkKMalAmRuchmfpcQ9YBSN01c/dyk0
oGl2ZHsLttTDbBo/TJW0DIL094of42a9mGZMZwdil9ecLTl1kMlw2v8wRMMqtIwv
prWdIiMiVyxQHV+zPx7vkHXU5yVByzkmZGfaN3R8W3WVhOsgV9xc3uxBvol6oeoG
gLL9Lc60tL7QGHvLZzJlMLW3GkA/ItgB2WjJDt6AAeJ/Y6Xz+48Odwwg/22KJhdX
YJ1K+gaRV7mznIabnRZ1TdkSxZ6h8i4NIi0OvYX9wYK1ZqTbcujnwKXj4Pd/HJQj
tVWkR+39coguTqyqJXBLJiNHHVrXPFuiX/W/4oTQjWCmeYBp5sBPgZj4zE+fXQYD
SXkPw9zNhkxh/4GcQPO0fgZEJHYaZKXQzcAjEDk1el0QDC52Eu484VHW4rp4r/gQ
U3F4YI/8RIGDKC8sOxa0m4N6gZuoDPcEFDmrLx5miA3y6GPHoHWbtn0HbeGvlPnp
ps9GvCK+pKrmE1aljH2BIFRJMouGl9gj7JyfWyBciJG3/yuEMr2gWpSDSOMXVFWu
UmHB/ixquxnLNptwo42/fM1iAWXXWT/T97M2nmRejDjubYxEo1QiQvbTy/4lmAoU
WjNN6c5NPlacydWkFWRuI+suQyVwbvDMSrNiaTmBqc09wjp0GZ3G0CxwiqXijfJl
sIM3srQHtfhHfCmQwzA0mKxYX60npw59HVPV3FbtA90pqotrmnHOKTtQu9D+KE7H
3XMuEI+nJZIKkOc4N3ja/eEiNuh1e0z4zalrx4TwXfcP/DCVqWZFUcMUWXLu3dLm
52GYInaywxw0hqxL5y6Lgeuw4Ty0bEsiTufRs83mCBXrlyL7m9TktYQkwrGzl5gV
kwNIDHu6sZUqFX4Dr0gEUUPkyGRt76tH04KElUIEaKkph7HQdrKJIiG5SABIChVq
qp9PEY5gu3eJDYpHujFT1AaLVZjAAtwpU7wMG6UTPVoadaWRz68M6am4aHaU0iQO
TAUvEdgxygHueWfivEe1Rg31CXQJVkyaYL8dEadTyVa2IruvcNww3/w4XYhYC3Ri
qP/tZPX8hAlb58XmIYS21JohK1LZJ50fHv7rIrKQ5LvmzmojN+eh0Q35MV+mSSvD
IM/xOB61cn/P32/OiOT3e90FpJPW3hQy2X+ExGxDbiOydwgPTNXvy28cR/dbadYs
OurZd18totLcOvzM8+jMvXrVL3on8bq9TkGMQ/mz0zCsNJFW5GhnRfuWnQ/Lk+Ja
RPuzo2lxKqPHhxWMb3bEpj+UNxHiqztmn3pReNaf4amyHIk1Gw9FVMuCny93GwRS
H5rwKsr4BIMbiQiFcHXqRUoya26Rw24FOGmGFkMiWx4DW2veddqr/GeZo9TZCZKK
gqTw/I9HepNKJjUKOiFpoQmHRsEHh/P48EDO2D1ZuY95gCgZBkgnbw28g481zg48
RYMYZVSb33A1NIJVtVpQtZDs18CdtzX7+rk2fI2esLRlCvLnku61Sxz6GN4xIuNf
/3PFEY9GDTBtdxBFVUbmqm75lwprpu4c0VgvoqFbyF0QRi8UqWCUDFpKKScKudWw
pGGFvS10ra3ugyChqjEpr0biXA14OJaUv12qewfLVurXHdwimPOJ/tEqzXhCHdhM
Ygr9IqAET21H4QKPfBPWHVSb+CySyLR5AVPfytSzzifOzwqCjcPqUJhOONVBkZ4M
INwfTNVxNz28BfR8a5+xDum87/dTx+C80cuPql0/RbzKDMjlK9VjKcI60Ph+jIZj
Z2Kp66CZGiAq7B1mWqbvS4KPUN4eTdz1Q/4nzH5t6zCxnpjoA3tPDKcbgh2D1QEf
XnSV2+S62eMgUKFZqwpTwtuaF6LqaJbd8TbggbrJotd43G2nkRkQ13tHmUGG1nY6
9XdwMGFZ6JNthQz70fjp9tUHFpEhLlLFPddetI6LDS02Lb6a1BjEoiK1eW7iMJbe
iTh/xoX+6G1Z/qW4PogkMQ1f9omMCt5pSTH3IMO64S72ORAFPvD5ytZ7s6OimLRb
hycH+xBoug2x26pani2LxNQBlEKYB/J5f/28nhZyAVpLvv+8fE/zHACi7voPC6Tu
lho0jv59SZMLljr4majHMzHcQ4odfsFN2YSBj+udHZghYCCjyxb6OumDQpmUqyBZ
TAmf8p0ACAZ+bYEmq/8Od+PcYbw84gOWDu8duJibDbDD6Lxb7edNpQED4NhGRaVb
83C1o+ANGSB74dIiLZmDFmLl5O5PRl5ocRLapbhKHyp1UHld6llPlYF13Sz1I30u
tqy4j2jC9fSkWTvjt+QgUjnoOqIboKF12AgBjEzUJsNJtj9ScUDUKKRWQE1ji3+M
OGoVHA1Nqqm8NbpCI7Bo2gABAgnD06tlcXEgbkl3gMfti/geWgzFsEMjN0BnCjMQ
aJD81G2iXU7vQh4Z1aSvGyttpvxjTIDRe6G72Xey7nr9Y+4/eqf2NBom6XJbofOL
UdS1N1FMCOXmHbhAYtUcyANb2CwG2g1MwdQOHzR79HPgCBqkJ4s1qX3sYWrnLo0O
jP4LF+rk1QFihKJ5RyY5RxiGo8VyxcXrS23iqPm8eDuP69Ss45+suRxrlc90OTKY
SyG1ZflJT15Jw4KtJXIACztxx8Elh86LZJ6ROjpL4GEfoJWy8Gj8r9P57TiLHJ4K
yuNhHhe67IuKtKwIhjn4tCFEwILDXzCPEAB4Yqr3BhWqN3tFC+eLaKIvFHMkylrB
9xR09f+d1g4kfihs9wz8rFXAEgSWcL3E5UORaBQsSmEUXcpnZIdLPfZnZUoIVjj5
G+k05TbOPcrtfmlPV3ehGlG++U1lC4X/EA0Ni9oCT2NQ/059VdAg30TdZANVeRM+
egCDpu5mxJoqvpI6384IIqn5lf7GsC8gQlYZhHguoybACIH5yvXsWLqeZCM8WwIe
LFsmzUBGn2ZpAtkRVySN2ME7vsSBfPfqUnbagzM4szAkOM7lmSK/Gmtj/5tMkUT6
1qtbl1ljsHUZ1u/e7iuiELjaMspVxD/hmzlArJWnO1iwk1P1y+4gwNBcqiXPoBJx
dYUjHDugPtj0f0FoS+X3shuRbaYHmS6hne8bo81A6To6OOfc9T6DBnbC2vI+rvoK
8QUOoaQSiTJnWxrAWhubFrBfIfFN+rAkTkCVPAZb9XTLe+m78iIDwrg4wir0yKMN
7PeCf8HyJb+YL2fMhWgJte4UsNyWMiwcuZTQEp5egYoYBACr07u17Rz85rNSH4dT
I53PraZn/B3/FMHF9qNbeYsAB8Mu2vXjMOuJxYEId0iCswH5ynhBCnveKu7rcx5e
+qzeY3M2n0jNbtDLeFCNjwH7hES5bCzuEdsVVE/hOm1iLV7Fn7bx/aL9c0WTXi9T
wHG9UnnhNLONvsAR8TGc2lp3FOGp77LedmW/XsiuwjZYLvw8lUA0GTWj/It1KnKn
JHKkuJ6NWAprWmsfvmu07yF3AOMpCu9IUMjTxDKDGDXueomPXpIwTXqI95mQB7kr
vRCgv+FbAw/MqtxqPP4H5qG78JgW1T3Lq789oPhifhLYQiM3y3VQPpuIX4WvI0+6
Kf7Tw16ZOUw/5kY/6quMNvSZ6WklDiTXlWp7qVg171KYTa+sbLefi3QDx2Ex1za7
0i2XP4FhrgDfQ5iVpvSzKGUJhZKnP8VmwGneqypKTihpLR45FPIJGxQqEL7GyW6A
6WDxzebYIF4a+uXXbxN7fBFjd4+K5Sg+4fQH7brtX+ftvME041YMBrmWD7/vn2/U
fB9EQwHxV6ogJeimOc8VNeuu/xoV47LoA3dJW0Tg4yaE6Lbq5H6oOaHwL7bkuwzQ
jPqF5gFZzAqoX075Uy9bfuTeHsW8dm4iwYdQgej+BJ/DqPTunBqg7p/wRviyL4l2
uulyP5s6JTL4HhzwTyJCBH9LVgCh3x+a+yy0ue63eTtv2IdowKyCjGD8bCTB0K49
njzqrE6B3cGlm0Whfb1jtoTGgtv7HIqOacQrLbZWR9LELifWZPudqlvnuOEbM0xl
OlWvrA1sTPa13aXjottd16blU+qRhaDvcLRObLGO0ci85xbpzVYWr1tc0xAJ2C3O
WS/E/MhesbImStrZlrGYcBWeZzu7a8Z0wP/XNjk8VGdj9jn2HZgux+RAomN0lCWd
zgrRjnXItF0tCMhRfGkqoxImMglWaFFwDZD39i/+IVgKY19ik6RlQzWrhTw36Qw9
z5EZNjfcWjzTnRWjOXBh4bU+FFrL2d+bw4oWCP19yXihh3P3t7be97wse2BwWOFp
Of9gnYcEUw62b9uJUO+xWfrmLHF/MSNIx0RgPSFru/v3iX3qOHBbOC1YCXp6lvLc
Y1jsosG75XHoMZf8J51nlxy9VSVdY68p23hCKpifWYEKYEypU1mAtitDiZZPoAAa
Iis4xWJ1/lIsZ8fFnN0pg6wHZ+Hw90fdgNTvn1tuL2sIyArdsRH+0H31tOlavNAH
WCX6hTk7Fj7Om/gnxa6eJ29HdPaclTFzmP1dKerHYcBJ0+cenZ6dG7993S28MoDt
l9foD3Gko1qSF+37ecuJk+jDgSD2H303dsGdBKmgAekEBz9xG6X34uXj5vlMs8qP
xAJEj9/7y9fZTugtSCHfNtcyN0MklIpOZLSM1Xjs7s0Vg5NRVo/PUgfHrugBcZ2W
uLsMPbAaCKsx7C2wzMlsSSHZ89+TsxOrcAl6d1zzULei89riHPQ9FQ8y5OYl4dMs
91zPig99/uWIaA+Ls1gEyLLOquOAdhIDMFXDNxH1dha7EdylYCAY351tddQSlKdS
uddO97bWF88PinM5QF2XzA6jObr5cEd3kITYjgSd9f2i7T7NWERP1i2DAwt0E4dw
W6aJjsS5ze72R9Cmt2fgKKgG27Dh7EtumJPzFFfJ/0a8hLNDBC+EE/p32WqJOuP6
w9dzKfCuvg9Su89kJjx+Bhx3ZA95/HKUFpyzHFawyO/sN5SnkoOSngnDdkNUFO+g
oyaBrc2MJGhe+NnrMZKirN4N2oRQpg5wo55faM59HHD/BjxJXqs2c2QWhlPjmX+u
b/064yc09pONzX2oKEo9Uc4Shy5pnCdJB3tVclU79ZFz+6eYc5xxyS7qt5y97KkG
RDy5ED3fBL2/Dl5px1ZMQCdCkFXYrmlQ6XUe6+I/7iau7tUCLovCtSx+TJVlFhRV
YhHP8YJZH6uMGV6DjGaS57cox2uxd6GAul6pxe59jxgtc5pN+EuYZCcyHKm4hd/n
9w3pa2br0wElOAhLJOZy1Xk2ns2S7FiKRRZKVvs0dJvhOmr7IDe8YIHKoDvohBSh
BRcuxxnRzBBIu+SqcHWMETdTwUG7poPDHO+RxPv7vzA2QXVMxHwP4lZvP+pku7dz
nlTdZYQGLkufHULqcst9qq2lOGtvR5+wNFFeZLNKJl0R0uNSO3KiJOa+BWLllgES
4ut1CBjNnunRTNgUoAG1NDlwMQz4slX3nqgKd4e3tPt1K7ICZztP3J1/xTT3ndxJ
0aw/n+Y1icXvIwAJRXVArclidqjgJ6f7gwsXkJOQhMlbrWw/kwel66Q/qhNxMQ+L
sfl8jxmPDEJt9wbUtPjlM4Vfpt0IsVyxCuFD+9/e/uay3hIq1hidhg499p7gaaVK
cLUz1dZQ56l8y6KfyRMZUdW5YKF5nmXtmJKYU0M0mUdekGPP0+92ZMIJdqf6AZno
6nfuQW1E+PWDBqpok2ZajZI4RWIRZQ5yYbzeOkl/5WlY6hU68zQZsBhMZcJOg9v6
hCq2CHbv5uVJy+t6wukUo0pOlCXPzJDWDgxxREEp55pj3pZV2DUZRnt2CKOnTXyp
tHceyqncZxs2shP8Sr4/tbkYruE1YxIVvJB4qghwUhxQnAKyyKxjzy9X1it/jVwN
u0BLYOqZg4UtAS6LDWiYQ78yPQaYUdOwfCNaIXAY1G1eBZ1YT1ycFvboEhEhmGQX
euiUYzYgUIQvUMCSQX3ZwZMt+MXCbBAkuDcIZe2ZwIKwUx5h+xky+Z2RXs0cSkD5
CtJb1jMuIVXisuruz6ht8faVn29gvJIAtOvePgZEmugNw4/1VANuQmvGNJsAN7g9
VZnIVOXpdDsN0y3P2PT8fZZr5sHTB+WmQJVAOxKq7Vc5+zkctz6AxBqe+iq86iuN
13Sx7oPdntYS0g+jm2c1HWFGQupC8kqUdaImMrWjmsmw6eWzV40zwhUq0sdW5kjY
uV4oo/bUBZk0lb+V9hZ3jlEjcGY/sLLXPRoRhVa+hELRKgie7zM+PdbQ1tMbfCIB
6SDjUMopaQP+RlnIbETXdyt3HMLztgmI2uXvynQiTq6pNJ48lOTGyV8eDfNaJp39
Yy5Bkh2Ud0/7BnPtEWPOlP60GbFhHUYQVsmOxLP8XeglCFSuyCctQHH+F08uLxzC
tuuOvEW8rPUImwkFmF5NRMCHrNIyQSMm1BGapxpLG/rBGn65vzhhIqU1k0U+6u0r
0MauNxW7NNFRQ2b06ejTeGyyYRb972FDv2hCE3yfX58THqtAVHd80AobY0J4tsKP
n4EIEVJVBmJDz0q1ZT853j6nISJmGV/RR2rwADBKfHmIRnRdMkC3jt7LgcuY7Z5s
hjjEEFe9b7Agsi1sqZi6g4HyKX3w7t12k0x3Nxroz2cGNHAc6DuQxUosGILwStl+
dgtBHdwf92gUX69sStSpc8sqzxVJNxe3/+kFcwbBQU5fOpaWfzRmCGO6VHqUEXda
BpGWZkxR2jze8fpjw2lgi08QPY9+/HFFS2MRrKbXrJQOHo/n46P54ZmIbEGitKk+
fAYk7BUfP/IMoGwo72WjtXWcjE+Gv5kXFjdce5fMqiWdUtPC6uqK3nmAppSXBewF
9egeKr41JgbUlZG8SjUsSFLwYfpojUquWHRmuWQLpXHQ34iwFTP01d0hilEot6nY
v2DeSaaj3kFXcDRZErirC/DxnpwLtGaejtY8l4Er4JPivDBzFCKcGb1ru/sjZ0q8
Qc5rIfwiQRhvfR8yqLbM/kTTF8kSB7Hrl4vd8nRceDUFmyW0rmY8/8k6ZySgzb2O
j3HQUnr64MfbdIhz3XYLGsUQoxEPmpKVRo3TAyZw0kV+j17AVj4jhiNKj0SZxfYn
E5wSO0FRuRKL/n6taRIfDCxHFSE4qiyNqmFjP0Tex5v26EpQzKW5ElVKJVR07e2y
avYBKG5DvM2fVBuOfHg4MLI5ndWOQ5XhNQ0Z0QH7tWaZXMHnaTqTZrMM3aDwua9w
3HnXQPEmO+Kx8Uk9XRwoUTsG/dMGhZWdHqzV9Z7w1yz7jIIGLswf9/UWaVdOgEtP
CHDUhjygY9nlv0KcqNB3O/dudJSu/By10JbUH4Wws2o49HC6JNk7LvGzGrRpc8fe
WX1Jvk+MMtWwPC/jDgmT8ZTnAjoR324QFMjUiKoSnOnFYtiUkHT8C8T1H7gZPTr9
2bKek8mfrrFRe/7E5HYDxNP6dAGyG37ca1/2048uXCl4n+C3wqPUtT84CgkMPz2V
cJB5JZa4MD2SK7LgnZO5YdmJQcrs91bB+ZCnF5l3U8o5QF7V2t6pu5RoIkgFbUX7
O+1O8GaX6qSNLrlUYrEdjTm2cZchB6byeHenjO9x8T+DpL0er2ZJ92YoRHtdj90f
TLUGz4eY9YbjSp7Rlf8+i/YUeVg4U+MUVfkz80uJyg0r45Jo36bOgaK61yBkitU4
s3ba1JKBTME5ZU/o5u6TCg/oXSndjKqKjuPy4sWeL4fUkepqhTYJDz/bemRa/K/P
VvkM+kqyHzDoynY9rNZkNJsxPDvLK+uvNcZOXQYI99MULfuKKju+qLW8ryPt4SUj
ObpDFKOLPOWnfEipycl3kF2yR/1QbbauvbTDoOxLN67rQsYk2RX5EjN4eyP9HHEP
Tao8D5fY1TfInk/LujylBCN9HAJsQ1d8SWTguL1GDqTUKWctXDe2SFRUFrG2JsVd
MgnOvswKle/vd06ksXYTsftNN2ZaJX3oguap3fboEiQIUVVl5qCNoYSdI+r5xTar
smm5iuRVlS+JLRkrubFcIB7AkMmbQ79XyX/B1zyfIAsA6p6JPRLS+apfbSjgCwIR
QHQasGsMnYrRWgn6cCmr4hl4hMTBI4p7m8y5K9tw9g2M1ueW3O/qfGH96Xe0t89i
3T75q7c7pMaUk9zY3IsQWoCJjyV//h0UDPgLmNnn4OpfhgsABgpFH+hDZssru+qX
gYzi1bT11KCoDForAmG0urf4GkDrwX0gjN1Jg7JgVRjGqC6mH+KJfXAOr+XhrUsT
xOzamEf20Bqdhi/3OaN7eRQt6ivFstGNav8dL/OvaPtnsqaWhcphTZuCZ6LjeXyr
EOBXkMae3M6/5ezC+J8y1OCVsWYyfAKhXo3Vyjxvk/rdhE/kyQkBHWiB/Ns2cizl
8/kOPTx0WKj3SHGdiA4OLwIbiX7O91qrQt6zAHQjmSRDPqAdl6ZttdGC2CEFWNvi
NejueqwX5tDLhZpamYgvGB1XFh3bAIyLo+FmmfRS3kbreHd5rAMhyTCrH8JWS/y8
Gzfen6Hwi9XOqcYoEuNapcxjx+VVOsU/CPvcErmoevHSSdoJcGd5rWKarW60sB2e
XnUDmdx04JDwxMJVLXlTUH1KnlcWRzywqyBHKbTO8L9Xjxe1zGrUBfZmuL6xr1IM
QiyLozUjXC4l37E6r1ckUJwVQO05gD6UNcKocfXW8Po/tGviMfKaNH2b1KwKhKya
J8/mz8nkTTFcUqXUDcXXAdRq6Vucrpw0lSnWUgc33jee2uhE9aHTSG0wkL/J/UHE
5fnosM7s620IiWUPRmcESNV3ZEGfEm8ZurY0eeKhsTx5yRRPxoM6NOwaVld2TxnN
Me6vvPFLUQUClqkVbPhnITcwg92Cn0VgYI929ayIuFPITyKU7L24ZmEnuzZJ2iu0
f71D8EIknFQyMGuQG4vr0hGoHxAmZeHkiVGrzFEo0qfMntP1/UM+LJMiiPCwvLkl
QfpsftnNOK9iymZNqy1tATZ+M74ZAG1ZvxKj++1mQlezuzjVnGcSGUhE4tX++jdS
M2vNCUR1XPxCS3yjDsSiyGuVzMs6pZLvrA9lC6aJQixdWUT2efqLoBIRAtoe4iA+
Six57UCtcQOxO2Y8RyW4LlQXjnWyaHGm5L318Wk/CTqu6bc26njXBf/noC2JyVZX
8vyML0/Pq6wj/O0nikbSiMejI+nu6lYjvPuEdi2JqZI4EHOG8n1xFmbT2+mf+ZbH
9VAP5HMrV38Dqk4INSufqptMNd8FymnqM2yeM18jxyxRHS5Z2Mal4NBsGMVPJQ8j
OuBuP8QHHOK3/EJZDWSg1VfdOniCTvtAzop07ajiWyKt4Xfobw2eTMurKmF8CV0v
F8WaVYL4QncA3y0Wvuim34BevLtsLyI1kVFBJiFuknAQory+Jpd9rZPVsnl+RB/w
rRvQ5SvmVZ+omNPL1UJSJRrODI/STF1wbwF/z3aXDuXpDzFM3worhM61TL6pFrpV
+PbT30YZGenVwcDsBCiiD8pcqIzhKS5OcVB+Vl0l9qjblKTpWcYq5bRv5PUu2Vdb
X3274hE42kshB0hziojO2FvQJZV1y/iQB+tg23QhBivuyvX9gDPz5K22ubx/6HGs
zVL7g2zGgQa1RpuJPRXgSsTgVZ2zkECU6v7PXyFTXCBvrCeIi9wImbYvXKPlSS36
/t4QDioVKX80tkIaUK1o4ASGJKN4WqdFwcZzQ8sUG/F5klborlpB1fm5lNnNlxgn
ENSGWJms3+Woi7oAj/cbsiE8Ew+oyeNhvLeRPkfSxkOW330DXVdCqYIH4nZOXT7U
ewRCqWE0VefRPPWN3qybEzpFvtpy622MuZuKarRiepuF9Ja47sMYJpNm3keJjCex
5Ikf+o/J8cF+FYGvo3UA/rEOF3Upo2kIqvDm6BZYm0nt8g0bQUqAdUuHt3HlkD1V
989MCru1igbZ6V6jJ7aFCSDYTuq8ptDmzFglEbHuNEPt0XdYJ60rRpAZ+VKQaLbR
jRzrOiIhyWFtFWEQ8ZJfXP7QV7HzUFnUKcu9X2oDSWKwgq1ktdocEKJj5rEk9Ug9
eCFarF8vefjRAyEsFfVfnVsGlPfzL/VZYlVTswg0TXY6jtEXiaGXQb1VMC8FQfxx
qhYXNWE7DocfjCznDYUq/ywlhOJ/WTpJ3DPij9wjgHpIeth9AZu2Jrj7uaPhVZGJ
vFlIBxtQRkJ5kR4Luo7qy1XKQjVUUqht/5Hue8HS7FuJcTg164o4ukyDehK/5VdN
VSRu15EtvtT1qa6+f4xJYeOQ/n8nszWsBGbsHR7GHX9Vqh0wP3wLJjAZrdiFZuYv
T2Sv+RT4XptxHMxayAjLpT+Pv/2SZXeGMUtmIK4qZkoZQFo3F6dhWspaLZNnziJf
/qN+ugn4zOv6SKp8ZGqjRzDRc/wKA6OZo+7ukIZzc5dX2e7qI4OalrrVVOQvyXR7
NhpRlWwKyhyzfqrcvlInUIremJMETYGB7nqlKLn5aN5HtPV1koLPc3xgYwHheswb
hGFAsHLJybbjSR9O7LozWcM70yn/M83ytT/uvqIGrvHaJUlvIVhCNzbU5Y80E2Ve
obg5JeEPfRYlTsYmA9HEYgUZYutk00Yy5MaLFAajkNCSjYyU5vsy2ENLpVpMA8i8
tEZ1pU+JmaHtTU+5Z0/Rv/to0T1KDbyG/HaYCCi4U3nJRXDfDOYENO71rvk0VBxF
HD9207AHr3VxzkfMxtXHLGvNWU0N2KcXPTXfdFNBvHhzpvtntDP+UykrOH6ikfUZ
nR+09EKr8mcc60N0rJL944FtJPZ0YZyKkMgDC6yqFn0ngqk6K0CycS+Rw/DfLqK8
dK0RDIpMkz5a+DH0mg4sczPBilWu/VhZxQX840ZRnAVA7KiGMoUjeLLX2fkxaP2K
rVvCu+GbEmWd8S1l5zbwVAmCkNjalZYFMHO+3Qqp6gSG4k+jnBbLZFfLGB75yjPW
2uC0Jd5GhFzgEJOXK14jTQKJac8bpukgF33o5v+e+ET4aief9IVay57nFjBIlv3/
qr1UJt44PST+Nw0jux/Ct/4nd5maL14ffEQXrLFXLPHhVeuqJ9yCwXitOrVZX7Kj
L1frvfDGra/h363uIdPy7m848ggJjkgCVHloyKbNQX8z3L/1eQEij1Uf/qXtuHEu
bBVjfKMejp1U82vNZnR3dA306TZQbaS2lugKAEu0hfaH7ZLAvBFBOTLH/PNlI9gp
9wCC0rEjz+/pZ89Ni7OeT1379dAfaHfNYsEnuFTvviGN2CEPDSFnhkeTLOoZ64gq
vww6fQ7rrk9qOfurvXeypB476fV6kCs5ulcC1eew74bzK0mFouQYFDN2Dnus60SC
8bmDQJLUKzaiqAi0FHrcJodJLsfIgD4H92gPC4P40yLg8lEsJGwGx5HcW3lomPjR
6d8F0vyT0VWAvWh1ISgtT2JT4t2k5DfZVCamFdm5fWa0KnSxraVpL0vQPgEukmwc
n0oi39xrbinLsMZi8CmxiEy1TiWKPvaj7rVP99nBvYqcfUlxYfEHG8q+1XtkjWP5
eJNpQMoJWpFwBEwFS43MtjCG9czHOgayz4/pORL1ib/+ytSFmD8P82fGoeYuntHU
/giFD2L+ZsLTAmwFWn8cqJcVXpPs6cWQwehAqU1Srz/2gPMQmu3j76tIJ3j4VgZQ
b4dyzMZPyjGAEtao4DCZYZCjYzml1TupcY50D8uBdzhQyZ4I116K4FmRjak14eOw
J8M6LWSZp/NljI9hZCwmoikzRXGx4UCtNA15M+TeCa2qTx7A/uGRnhwSLoDkBgDw
paei3grZt6JY9BuSNFgEa238u6hwUYBKhtQ8HW8/WMpmpjaSnCorJHzH2KXrkEnj
+aDJSrb23v3gvwPMW+Rgq8BIu7DVgizgHEA95aAYw6SYafpx0AHCf0GeY1MemiXz
2gkpg+/f8tywIPHB6ioaRbdCREyQ50XuS228ihDx8acezJMpjY/9hF7J9oXUJ0EL
6RFzvS/b3c+O4vQYXnbB/FhkjxweElzlRUPwOoMx69q6TDGCEpfG7OuRDfgiUmtn
y+NsoMHPwQcf4OoTznqO0CYHNZeQiGzXZToTrwNc+SZkgSfMo2CNRGE9rCWhyazn
hG1Ty4be49GKKw3m80cjaApGmGznxPiu47IaARdjjbY8QJUR7vLPZBvfbQeJytaf
5F/KXHFPX5Jr8MjOsX+Ke+8Ykwe3Argg/62E2GjHxTZRFBF5w6X85bivwRm93HPf
18yYLmskz/TJ+d7uksbACYle8VfyAyYCygDZ0qo3aSigRXqs5vCUgrMTX6AwE831
zsOHpnsKJjQaAyIkAlE6Ci+r2Mk7FaLMAyS2194MzJma4wXKOzYC38AyfvoODHbn
6MWzii3JvRBCShsgz1ER6b818uBRrP23PkT1XjPWrY2qNXmjL3G3x9feS1rVMrZv
fu9pHHwH5v/11XsEqoCSE5r93LYKaNncvdvj15UL74keJr0dPSGxln/sRYYnC7Jz
oB+OJXeB8VrahkPYpDR1QsnFo3Eakcq8/ycNJYHY1L1YIuQblVfEOSNoXX2VCb1Y
5k1BDyi6MWPVcENkT1fbCgGj0Mac46VhUCPIEGkqQpBaWDwYUQhLeVR8NQffqaPk
b77FTsnk0fU9rVDY7QRVB8U7IlWtN9giYIrLSHx9ve6NVmKk5o2MkZM4alGpG01K
HlzkYjsh739D4LhyebZyQ+9Id+MMi6/XA2e3pzq8fJTt9rwgyxylJ7XfHJYuMmmJ
wZLtLIbQcGlnm7OuEDTp0K56r7hrQsJb95Z7eVCHOBFs1wBDGkIHZOB2BIdHz/i7
syU+ssyrxVcghCsf0LfgQDFSQICqCFZBve5CRZ2OxmaPDnQW+E5f7RV41DjgJv8d
dn90tW7HhcahcnGOikwQOpOyKp9KPAx3ML0yfHfdeZr+f0LulMy6y4SkRQ5KnIbt
QRtmQlguytWeaH4IBdP/O8aZUpU5+K/26lTro4RE8iTftOZcfoRZavz50aOOrfOL
rrSsR/UNcBxZ5DMJFZWwV3Kqp9qpQI8f5oVz9A/5V2QFg0yW7IKc5BeQec8btxEQ
w3wOSq7p/LZVo8ZKSMXVQvnDVvANX6XSR5Eb/REAXBsWWQk6JMQSZfWaeNtsRKOd
cfqgwQA+YmMowHYKBQiyq//cdRv+C3WywFpRjFh/LgCwb7hJtSy9XQC4kGLk1v0x
UsN0y9d80C5p1jddJN7LMIr/kIOnA2zwKOZgfAR9vta9geTHDz8qSRKtkl3wUWqF
JnrnnOtlIfpVOz/XMR53bnFINQcMNB9/sGRzphla+Q3455qFO6kkAtG1owkdEJEU
YxvtP0OFmaDJ8PpMIF/fWpU1QgvZlRUP38f93qtaGJyRDKKXlbOsv/SKFlSH7Fw7
YRscj9CUvCcc2S62/U4Mrl6By1Rn7vaxYY9RxAMIYjxHWWrpax18kwqvrHURYQGg
9F//y/7WSJV1LmV6KMQmGu2WjT4pmqL3+TNa9LgMalL64v8kP07LIg7RI6V7n+CJ
9QSd0qmmk0RKsavkrDZDBJUShwjv6B+TtksTSck4qpxKF64YvQ6fJ0GxVeX0Pyub
PUSgRG/bruPWFLSpy20RLlMk89vWkadJyJ1pl6ptp93xR4qd5dyESw+uXjD671n3
vbe8TZrUg4607eMVio914sSPgW8uEl5SpBfUHdMD0lTpZpBDJ48sSTvbdAUFXIL7
d+RfXJTZPthP71JG0mWF0di/5bbMC5QDvTcjRpJ0OmRqv8C0uX51GsYAbRyi2pM6
X/RCAimT03cE9LxT8viU5fEnvCEQFPMrFMlVQLPPHitokkxCH6MUy9Phhpk+S2j7
0kHuZRqQgCuqLKgR6VnOhaWRB79/ZfPxzeVZ4Y04aIqUm5BoCBVb5E5pMqfQLhdB
dGS+4FdWFc3mc0Tar1nLJgYvsBy/4pnPNKCW9GwKYrJmIUpsw8eMQezffmoHgeFh
sZPnlsidlEjdHgb5HoeARUyPDcriun3fAiaGTNyn67AHVm2O7tCgmGCbcGt1DUER
xVK52S0ovLBWu2SpbowNjJ4Zf4m99smIwEpHOg6pNZOFdCNYFC4KJlQJfpgOybLx
VX9/Nsf24SCLQ1KPbf1RiTP5FbteEYgA54USIHza7qdpMatfDtODRg204Uk5NX8l
YjhQBX7P9sRCOi3Q0zEyoWdXBWruEyf+sO+rOzgoMQn80hFPWxbuwuBs5NMYoePn
sGmaI5xlv2NM4EqaATn8LVucL7ciKEOc+VAXINfxQVjg/btLsIhFC1jyMu6kDGN4
UXIgnzhTllYTEmChBnYrMcVZZK0SGK9viiAC2Ybm6jqH0pOuOQugt3mr+kFtMqY3
ddwhcbcb8X8WIZErbCyeh2hdeFhHFm4gejyhdiYczPTfDVWFT9fblGik/wnT5BUO
wr76bbBcBaqujEWnFTEVXQiYrYticKCWiVawRklBLsiCB/kOXW7F9bmcmaoX1Mgn
H3AHqSdV4huUUqhoucitF/Bkm39gP14xVMWpX6iKyAYb1707TYMmZIHxwaPfXWET
bft4NiHXXNUeSl5Cm2D0Bm6R7duAHPfm74i6T2Fwkdl2ssouBvuOinmEkiSjcoPR
+64luxMziCsMv5l0wkuGp5Bhgt2I7jbgRo3Z9LyHkXwcowmCrrSVoPBN/HOIcHs8
PJuxW2rWH1QHY5rbmgh3eaPbvzqmLzAHOFtOzUhSHbw0p9I4DFq0DVtllZGQo7ee
PbiE6baisIN61ymvXVIoBhCx127Tl0znRUDERAQ9MNK/IatRWmMwAEGqYcNHq4uI
s6oJ3j4aql6wvSjAkWGK8jZ4GuHhD4yXP558ypcRfVTxL8ZXjVMzyPvnCuYLpj7X
RZ+X/vHlXNVHmVjhHywFYIgzYg155Eu8kU+WFFG2cANT2XWfmNUT1kWxxxtMXXmq
yV+Ggap3iSFnocczG4memBKdM6Ejn8G5gvPe8JrxkcCA+WNDAmbBxWc0EBpBVuSN
sD5oTYYrY4NOdclgGnQ+Rq7sLsbMLzcmTWF/hUm5n1BCGRARDFG0/zMMlBKUP5C2
7eaYGk5eBLIH843m12lTzf73MYDbi6dr7yppdEHUqBWMqKe0bor47mu5C36Ld6Mg
VoWcqJ6A6XEDvf2wba0C1iCVYAAgQ2yQifoEq30N4+sNo/MAUdp+cp6e5jk0Ebd0
PgMF7knU9h4QMPKQwqpJaJmmGpWPDfhfikFJWqYzzLBzOgyn4uwEiariMEBC6/ub
HhZXApmCsbiw++C+5h53wi5lpsXNDvVYdPEaWtxLOP4xx1k22SDUeA8Zr55QeAwo
7jD9M+VVGFj/N3LADl0c86ypjNlqhFlZWw3rla7Ynxr36RWjNbe13nIZVv7M18wC
+uz1rRxyuvj0Do6STvRwPOUNIq0KEsCt4hZgKR4br40EluqkHzrfk5ARHCFJXcnn
dolrgoMRjcDXQvwx1e82KN9Rwl5mfPw/Sl67XcV5bSYt20S/QtmC0tTf8lls17R0
7Pi1+JxzW/lkVupGinicdAYLWljHPUoukXrZS/zsopDHUPRDlSqrL53SmfztAfyK
dJral9d0wcMa3Obu21nA/UCCbqTsuJBN0WbdZU3JT69C62QksKXr7veLNIj2ZDzT
gUZDiDf1R8RZRj6zsGdV1Oetn4yZyxM6Cl3FeoLGWSYQ26GeuOLMzx8een4sk7aR
SqFLhKiOW4pumctMaGY0KPVd2dE3qWc2LqWqfauJ4DO8wWITtOviS+3Cnzkom1Fz
CavgjVq/TFdrsz3UVf1lx1N/2ukKJDjAq9qeRO5IwyhB97fRBM2lxeEzJAyylEM0
GaJlIUz4/PwHH/xp2ThaZ3O7rar4cS+qtjRaPgV8eNOgvhsSD3m/fCpHH+6Zix7a
bFPxJmPlta481YdvlKyK8wYKvQKIm3Pr6gusWdtth5UnfHetfpCziZo1wynl2UKI
LQXlUcgjvEurS3kcRVDRf+tndKz+Aj7klqXjUPyeh5qEoZr9NPtfO8Sr+NGg01ig
d0H9tH3jXvX0Hh+9vK45gPg8XA16NuntR66LNK/TQVxkJxo4vFHidWMKeOCPa9NC
v/MIEKh5Y12XuMCgvjYwC5X9lGZkd9I6DTCXJHoWLnC/DOdnqlit8oi8bS87ZWdC
Tjmik7952KeNIknD83qI+BWtoDXZuXgnlYZWQAGL/tAzAp70hKdOGKCJ8mKHVNwM
Ddh99ZV+Fn9POVd1+081aLjie29Tt4o5QTahseEZ6T+xHdwrrGGYEAHPotj1QcH0
Xv94FA8ayUSvo2QfVyisjV9AjkWITkhb9RXFawVF74XdKRRp4hTU91hhV+wiRkMc
SZPg3vcfzkB6RNJtViNM+cbetXQK4nMV/O+iIUgKocKydXS5HCYtN7SuizBHSmjW
G/PLR82qFTQIATQGSWU5FRfFsTip6oJoQh155+ZoI7Qk38tx1xTasnXXPkwHYgqh
/nkVSI5wRfdNdKjj1FF/475Ah/8CKJ3Ybm4ZGsMfM9qRbgqHWWo8Jj+qvNBYNNkT
Lybr4lgdmo9axcB+1phBE7NBpOxuyuXYFl9yTObY0nosvwYM++Pd4r2utkp871+K
ybEfhgSkTihPxNLF9kx4T1Y/M0+wBu0ef+AEPZilgSf/zguXBEtE7s5Q5bDpychD
mdh1Qr8M0Cmn3RWvxHcMb8Hy8bsd7lJ0TXydjE6U77SOQIgtmdwiBYfcJE4NdzCU
+r6V8hkk+fn/+4mmQLp+bzSHGQYNsBeV8FkT9/h8m1o6gS/H+kzNAor2v/UGjxp8
9GucYwZsPSlyUwmDw9Z0ZfDDU7MrvXq2CuPU9SOKIHlSnVrAWQpC//LSMfXPw7Sy
UaveT+Kq4AtXqQuRlxMx45BQQx2511kEOVbpuUQJk1OLVjqGVaEU1D/k3yo0zaus
JbrsMt0pV7zkycBq8zYm/gYCDXsVbnFcFeRqQfAdx4YCqvYEUpJE6TY38fuDt7BH
4IpHDG45zZ+f+BeeDBNKFg0Nu1jxUT50sslVBHDHJpByesYfpo9xaR36GA73EbaG
mTjpd9lJerIygCa7m3uSN9hXxTLYXr0YyfxdrXDGDWC9mA2mrPjduU9HgfuTp7DQ
gShcIXdHt5+KB4Lo7JMTiG+qRXWa2BgHZsRrMozfUpDLfHIexhigQ6I0DxDneFa9
QNyoUpqkSeRX6KtD/aA+/uBKA0L++/G+1WA9PPAPOoQr3QPidWI5Xg728JKI+v+9
nyVuz1cIyQXqEjUgUjvb/hl+BKmG+WNcZSHY1zlFlksDc0+43c1f/mKUCtadJDsQ
C0ExueWN5bp9KKDSVz0SjCnsiludjSi2fnzkVOWRX+keul2pRDUTt9pXY5OSilFY
RSFimCcfAReOmojPbr+gRB9RN0lXEInO8UsYbl64ErZoyaH79abMg6Gsx0+PrgzE
HZ01HRoKetdwOHoqY/uE3l1ePFEyJwk7aRC8EKsFqciw3SXacbW5u065KGQoTWZd
CZzkRl3Ly/nNzOl2YbStDkuyMROfNALLfmTxEL8Y+zY3lsbsb94gzLOYDWQCkb3a
tMKFQ7Olh8H80TNm8jOr17LsuhIqMyOQDXIUh3qxmbA/IzFxEiju+EhNHTLB2jiu
qqXP+QqnaFnfabtbPMJsIEaJevzZtw9KB/JQoB/XWllmDhSCjCS8OhLJmdrEchlX
oPQPDNe/kgXIOQi4gtYe27Zh6MP6YbUgsHrL7LAgrvLZRNxz9VoeFX1sDEcJBzfc
RkyZ6h7esQ6AmjN8hxNd22jMq2omCyW/oUXGK9h0175nXwFpgHhsThg+h4sxAING
pDBP/xC3+MbkFJXJXHnlBCUgI5hG0hWSQvhshQz8Nz1wXRe7Nbnmf+HyTAHcvxsA
WkMxEgssqr2B0z/0A96qGEAOfqAJqKEvY9lb02J0WTuB0yFwRGwA4jWRsRFX6tc5
XYvkDoJHrOUtXJRIRCGrXutd+kYFU0dFOkXSAeTsvtGsK8nCfgtqhk9EYkDnr8mk
0ea0tPIjfQmv+8qPdKx0E4Y0eIXIwvQCnYi4GJzEOry5Vqy6aTbBoXwLfXLAIK66
k+bzPnonygBP09nZDS4YmbsdlMjmhPohJFUDUN3sY1RVsLL3ANiO6UJepZk5fUzD
HHrgV1fKXuJuxOP3s/suUjSb1bUkUhpPZzfQ8m2wJ69xsstD6mDx42/CCta+3Yi7
ZHx6D1u4KOndnOJhf2rKaAXuafv6s8dqLhq/Yla4lqBSIhBZyXq/LtY4Ngb3zP+F
1PodmKPBlCZ1neDEdSkp799AdaTRLF2a9WapU6nk7oelk4RLoBxL3XXH2//zneO3
TdpGmmSLry652prmrhfAtvPJHVwdTLOK0T74JPFhvdaPIWMH1JHb9nsknHE1hLIb
+3HGJn5h4u9XN0JOfxLG0X3IVas3EEOBi6uUZQTbQRPBWVqLhoKRxXd83ddnGeHM
aCoZjUC1l3oJpOPhSPJ2L0T0amsEJRGY59cYrovj2Tdg37rNbnYgBwYj/DUseov2
ST9m6B2/HO8msE61Pu7k2PjKQw+7tyOuluJ+V/LCS1H4eNtCjRbVdRebeG/xy8sd
Kg+UJQDkyxu2SKes1ubCP0p4J2woztLogWI9RbhJFWmALznF1PWRDhuM5s5+NNbX
QEpflVdv0lLrhz45+hrqie/k9OceE2bM6mis10Rg519Qf3Yd6t7dAdaj66tH9Cxy
PYRhbDeeOYMhEiROGOZ6bV542qbUUgQEztgoa0BqNK6bld8xqmt86VYLwE1ZwanZ
3fn6hoBjcZEgz1A/7wkB9HZlE4YKv2r2pE9363I6fERujAwpIn1xCRcrwrVeoDLu
YuYKvrMuTINCTLyW26WBz+rBSQt2YANbMNNTOkgjRnmpFmfbp+78ihyjmkz4cYpX
FLSSwrySnp3PFqu8Lh1vc3mff0ForSXA3Lx4n27azWRBe4oFp1ovqQlH1uMKcGaa
BpC4u19kdx8isJcg+6QsOC+GXefMWB+oHWFhGMfQ/HGnGw0ynI0kfPpmUeIbMojP
L1UREwuFPpvHbNly1uWq5v8hByQ/Y7e7cQjZ0VCwRm82ee00swM23gfZhke9UJBq
0wfOkkl5nLOmUmql8rwMumN+HtTOu3g435xtGR+N8IkzX5pTso7eLb2tz+QGZWxZ
vDkWNQvKBefAaVUupaFEnrpTzKqujCt+0z10wx6iED+6PastmUZkMJ51wKRxeK8W
q7FRN4nC1HcCLkOdeWLy89UVBEDRidE1E99PPICneyMLLJklf6Dgv8daKYbjtTCA
Fl9zWOk557i1v5RRdTr0U59SNJ2s0um+dn7RBFAjZHm3UYFTr+0JOarMXzX9L5i8
A4WLxxtEQLjHL1EKw4sQT8PTAKrj3Yh5GHiHFiG7FEy7Q9xL0xbV3zYwSUteo++F
LDKEQVCP4QwAz21OFmy34GISLNLLnIheYkGGFtM2/bBwMO17NhlD8w+mxp3TpD9Z
FndITy6p9V3Eq8mexSjIcSuFflJhZRMkAzD2coRuvhQZCT6DYKSvxUcGR+MaW+LF
pZmgbcmqMlo63TDL98Ez6c19Dglra/ftLtUutrR03L8D0uL3j4UZrftr21ptMGJ0
c1MZq3hJUPtewb7c5pzP4Nax1wEwjvwoH8/1VP+lv0rugQrNyrStRMlJCgDFQ6Rr
AymnUfCkpvGXZgL5Dj+HpKLXO9m1Ld6KKGjnoyW8LF5Ik1GDcXEtWbDBEko1WpPi
er6PYS1uH1zPBTaYv4RTVdNajKWgjElcwth377FmFU2xXZMUOytVIope2z6d+juW
8r/TfKgPDpWIw/EFUnPFNcCazYauCBUD6/UVYB+TM7eEtRWfvJm3+sLxL7TSi0a6
wQb2rtjUUD9hu44jeGz2EIKpugD7rI7NizVXx30BfqjdL39m2A9Og7QWnlPGOaY2
I7+PvGDIeNW5kWH1PziVkqT1kE0Xj7h6/SPGQrrw60ZNoGnA6ESKKZAjbHWc+huR
s1FGQUX/JHnh5ooP4l2J5Ug8X9SCbk0f3t70PXxoexJPVB0Ux/z6fOZ2lMyeUPq/
ygnR1YcnHl39kffyQHpGFHwn/jIX75BxmsLGQ5oaT4hvy0F9BRXjwBobI7nisAdX
LmoCNHk5qNhfHr8++kq+Y6eWDdRBX2YNc1NTzmI7s8MQ8qxJhiE5LgbTF0mBjwLB
hBodKV3KO7vJqDCmaEudvYdc71hHciAdCQ596bpJ+3yF5+qGFFLyIA/XGiCjbWKO
JpzCxnEQuRvhq4ZTyY+yraJ7QCOmjRCCbePGWEOVZNng4bIyIip0tgdd5lRpmr2H
qryAl4gWe8EcTURQtm1Z59/ftULmqvE9sUzdxqCveUCwUL3YrAmZ3Vsx/YEhMDJn
c6JLs9rMaFzgk6h6vkVVL1v3hQFVQvUcZ63sqbdyToJdswDIl2ABxkcfb81U1b9L
40BBjbmWs4VsH3pF9dGp7OeI/Vn4ydudL8k2UCvfWG1qgUtZgkbE+L6IGSN+cSn8
XxARfeQd9DgqMBqxcQ6MiodpDypSMOLbsmSFyBhUVCEtv4Lr3TCMbO9eFa4dAmiD
CP/0kZy6UlJitUHiyiWoIiWQGBSHZ+4RAaLZ143DQ5jureFqwz2I6JvFznrPRuGi
WVWZruMMLUy7tfcBGUQ94FAQn/O/Uw3NdwHwZc4W6s9M7whYL9LokR3Fpt4yNj7K
sVExGU6amlVSs6Pd/gc4HMeq2qz6mg7hHPHi5wSPrKmzHMBoDafLP21Rrm2xx8uy
TYnW5UF/CJvetRILbFklZRTXoe179PvS1vOfG8Ki9cdoERaU8E/wbYRG6VRHR49/
1NUuXd/REZ3RKbSepXNuR7dVMBBJL/QYxdo5Pef2aZO9EWmL9XCUQvqmz1Lx+cT4
4P6PrN5kZRCxkuxZcT0J0Q/0P2QHgTHSRPF1EK0p+bXrJqgxoaaOSDS1ww+ig6jk
4KVSCwKcScUNlbsKjEO2qXI4P45qMGMqQ405XlTSwTwJKQUZyclFuUqrDiuR5ZIS
IjlIZiUF6AsfvL89f4MZCtHZqjW1shmZNa0fc9Lb0sH9mXtJWX5o4CVt1flURBdA
Xqv1NnbVtPgLympihiaRxpsgnqvx4Y1F9aO7dcI3jXDy7QIbHeGggxvGqsebbTRu
wzLMt4RFb1EYDBvKPTx4kIG8q1qGzF533recerwMIgj9qBCHZLoSdheZrhXtNfKJ
I8qkdmMarB/i3rFQh4D2WJ5E+/rjeMZw3yTCIl0ITe/WcqfjATAgwBKaW1D7aQ7W
QD/oAXYVfTPP80BHpnSqABy254WxE/7JHVV+gYjMJjD/5R198G1lbKFgU7AeVTZH
BGKusB5lM5aUtSTFVUxZ+iJUNLUUTfv+C0SDH5adx2rfTbFfy21ZPObyF270BjKI
M4Kyn/yNU27aJslrBX5ucGwTD0TwsGtNL2mVjqZG/K1Ks65cFUFUmHs59J8gHmPl
vCB0oggPRBhF2XmxgmIkPOFr2uaarWtkhHpkTnu/Q+kUZ4y+Gqx3qyqCMuOx8RQU
D99JFstsWR4adZvQ1nNVWPxI4lOcDhYBu++UnGa+CYMtRj7mMcmazDorp3C6jiUt
gZRKjbYAzSe7PU5AOencpCecMItPng4nN5q2eVSlywv00F6lLkWHEmmXvSJ/UpmF
hQ+eKkcSFMNBi4jBpCKoSAC5jINHXYwls+H+L52IPYUD/Lirf1SUzbXMjDia8zT2
1KMATj1WcI06WXtVVGDMh7Jo7GmpeG/GTpnEzxrK3aatyScsk8cVQCcT8UrzydVL
UD/hfp58kQFbX85WNphsv4f8SXZwxvYobRgXRxBMxMcfMwp6zgKwAP3YmIEW+RYF
XuDFeUOba2OfdM4sOOTpzn3NFx1TY+1d554r5bN/+Rdd1LKt8MJfb/yVFIcauBZS
yA4+7wjNNSFTFRTAgjQIQHASi9VmeIiNLS3awqQaOK3W8ktjuFEMuZGjqAZXGNXW
nz1B6EO7QmmHQ9VR87Nzn/A+B8QjhT5Ir/Ij76ANMTCYcmFx7Ez+Ug9idbpg9kTw
DM1DQwAiTxxj7YjzKYhGqsyVURoALbXCtsl5pT2doM3M/hMXGBDR5xoLSA8xSIF1
qZc7Whyu063m5A64wOZwuq+0WGclnphk4tkB38OUeTFbeS8Fu+yEsqt1PDAM0i3Q
SAaejDW8PcA+032F53FV3iL/ZmUkNWPl4uBjn0v2Rm5vpGwqvKQLPifUNma4JbHx
bfdoBIQ8etfvB1rekqNX0dExj5lCT7ZvfF3okaNTn/G5oRJtINhJGGfz6scE2P/1
vYuKP/Wu3mo6c6kU3LkN0XtY5tamhDsnAdR9DP+75NYkjaSPHcirVjhaRUQcvMW6
jawH4d9nJfgjF4wTJRBRyEZcAVyR/Ks427DRcF/9lniwh33gl3GGuloqCQny8+a4
AItqZn+4ThuoAch2w2UY4Sp8QEkmDwGxJZMtaqyCkevdYVajqqnyRXd4MTTH/un/
nQYtdH0YSc7xYwNnrecJFyEyl7PSF3edWv2ESsztB2nPN2c3pAdeWhz6wpK14ZJX
nENpdpj5BEpS4jxDT1KiPUnXiH1wCJI2Fxy1CfmzEYvBTBm11Xpwr0UDBKxN+J1M
tDXr7hGtnXcl5gZZL0TG0jhHdSwt8rgHAKQ2+t2TbPE5gw2ulQ0553SKRwYmqv+5
YZV2/xzdGhy0pU8KmP/b6R8KaDC7UQQzjQSMtz3TeId5eUxPl0CtL+F9KRJNxJ5U
nJv0LIWVqoZN08ppNbHAUygi+ug3/AM65eLnYMh2Hro4hztii/uINnxKo8JbaoXL
PgKK/y4sagovSriAa7BswUSGHl/9Pz1JkXQTj7pvd2/k4hKv4kV0kXdUHMQmp8IU
8tzm0lcISUKc8l/8FJTeLQ9RlbWKTqk9GvlqgLQGd+GuLpgoaJQP/tZ19hTpCepH
U7bST28TrevxsrOvctjPHDX3GGYgKjehOOO5j2TAKjWaAfeWYqDTtX7vOeKX7aSR
1IiL1Xygd0VdJJud7dK37rUHqhpktoilhgj8oE9JnrWX690MOH5VYaPUDUNx8OZF
jHNOxYB2jN97HGeCTwNl/LDfJxt9D5NV7yRqFNkvnvXGoY2q/gAt1bmUETo1orT5
e1c4G7GGmxXUxgUiWs8exfTkIDRbfdvhePsrjIQpy/q31LW9RGKSYzLs3EqjMe2V
S98BSr2ZYrDHfPRpImOY7nGjHLSGQGbS7RRAadWROPVmRSse73lEmeLSqI47WoUm
IfXV/SK3QSfHteDFvpoz9ZRQMoQHxthNuZaQMUJ2yih8Xi56LO2v4Tidrt4SLaKz
LxKzqkAc7vu3SIVKN6POa/LwdkuV7bbzPB4oYTxUbZ58KLcaBlH8EvBYFoMpu+bR
V+qWEU/yA+tS4fnJQEAnhHF2456//ZUfCOvwiuD4gFkKgaRtJdKBFIcSq4kMm2/Q
YKVNWYlW5x0tjUn5A4FMPtLqAn3AyV4GDyzxsZ9jXSRevrTtlhQs7Jzqs9wHLLDL
i+3ZIBFvyoJmbikIr3ddcnTAo+veCSXLKEXm6Y4WZvmV3+Mj7sX7To/im+qskTqa
Qhi5zs9d4uVPB9KINdu/7YDfZt76Bdh2nVW/HdB+5ya9Pe7MK5/SaI+67Dfj3I6h
oj1N3ZHqIq3o3xpSNlQdd6H8S/PTHRFQBEfn4FoSfe7BqhGhtIpQEy51tcw0QnL7
ahZZZyPhdl0jzJyn58Byb3pk5casIL8ojWZBIpmkhOg+vog72eR+TqrLq2O5LvY2
6jAKib7DoQCnOn+DcSSWHAHT49BlAUEAFAEclbDCGFJMCas1L771Epbda4e1AkCh
ECrf/IxuvaHK4XY53wn9GXUDB8oJPZKDCRbmcSp97JYE4uPf7FkE6RlZnrFLzLqe
DZbNTe36Jf0QreC8QD+mu3R7H18mTK8tHpTq21YgYdqdOjrgBEWBYaJdZOD8V6WI
CKLwsfG5TqtDWWVyKZ+kPXGNHUu4iiOPYNroMwb2wBk+nLsT0UCiCXbr4KvdQYMG
MkKaOHo2X2HyC1nOEJb22jLpRezjDEt99EFjCVU5iAiUBm4gTSLGxLgMhPIfgpMT
+B0UL4eHslyFWIjlxnbpx8r25R+cF1HoNI7pyRu9gZoy0DbeQ1UYulvkr9wvHUko
YlnGQES3fBs82nFedJDCiwT+nX2fwHrW6oY6Y/4BBBu5QlDoYc4j5vVOV0KP+v9v
2ILpwTGVEIoar7HUKUq6n+Qd8Zf8WdiDH0oJdZIUivzL0n5Abk6CxQVflcJ1ncF5
xyOYyh33JCu5uxdV3WH/IuX6F+QG+KuQABmzGFF0M8+Jgyc26qM2BAnip0/C17Xy
O8YV3Gz3hE/R/M3CsBV1dXu8iC8AFDWS/WrvRWWekx7fv5XDSkWuTs2KnEm3FcI0
s6E85xnIBmKcZXTdSihLVjtNYCb4qHK3UY15HNU8KdffAQ4Sz7cWsWv9UP+di9Hc
TdfyAysaWjMYZ41MAJ4P2CDMpNflaqYNLsDnrSOjZAzVRAxpfwvrgj2F5u0GaxHy
JltUUTWfkcMTER24RVno8t4XeJ6jIUESY8mmm/bFImkZp5Mg9asBp9BqO02ydnTp
TQCJ8qkuNh8qNrJ/EP6j8HvFp5WCamKnGRaeMxLaM/801CoFUFOxHVofupYnIeAG
aFJ9SdfKhLRZV/be4sLN8ToUF83uO0fF7fsIEfyuDR6V+d6+DlEu3st5xhasgxdt
J2uDnAzXaV+InXuWagWRltB0HAUvJZb53g3ai4x4C+x4l0mDiGD31ezn+vukWZjp
EwZxqlzP3CkYCW4tgJhnvoAO6iDi5aYpmFhgUsItZ0f7L2lw/GIbHtRw1tMtUOj2
YguNBPITT/wwmEaaKCA2V0vMnE2duRG/11u2u+tw9XF/h9bPhxEaj7freEj0t8Yw
vHzVRB7Sl1FwLBNLU9S2NARigrZ5rNMq+3hRG8MKBV65Mn83eWyDnFhYgdZTTKck
JPNg4xOXiurex5FOg3lMfm8fbKgf0KqK3JTqyLyLzl5oJ35PkOUu6k2Whss1xdX7
YUiFc6w8q+2jixe8CL6LqZ4eb2HWZ6e/Sts4M4aRNiplHqA8rrmkmisN9QsN5OyH
tPsV9CaUJH9rl0r7iz8MAH4ZkdIyQUplWNJSiFjMODONiwl660v95zksYMU1a2Dt
pIfI3nzf6FGfCKEhQf6CHV82jmybWKzKK5I002h6X4GTsvJRd9EFDPwCCqDke4kD
ZMlqgS2sBt9ZH7g1iQzO2jSDsWPAdx86amDk36Bx86cYy0k3TvV3Qnif6U4nEmzp
ijvFGWloyAj9wjbPz2oyn8V1o6gB1+tnbnd41GDbW0czoDJfp3oRs8LgIjH2dTP9
lt8f/SjqSPToXecneIX7xQNa5v/n7QhcGiGBeoC66JGpYED6jX+VyIIRJecERgwC
szgjDpGWhUuFavuof286pbXU8dhAlY/mk3wFyxs6oNFkFMMXNKusywR5QN6BI9Nq
g2nRLXFA3zFutq+hTqBWIWOIhCuikr6nDMlVk08+WytLKM5b1LBoX+/n2lQQLqqL
sZM9On1lqhO/sBVNKrZ94lnbElTb+cg6jIVkdvbfnqj6IJiwQItviXaS/DcCYaHZ
3J1PBRPjP66EIxNLakvUxWpbzdpmmOHIkj0l/6ExBWdTkB7UF0zxlvroFCOWOP83
CxX/gjgNk5oPrut5so5IxmNYhNXBxbWayLXv4GTJDQqnTSFvezpwhYBiCepR/Uhz
hmpcUh3gk4EMq0XH9uVLK9f9UaV7detUfxpbvITFGyNr08jpAq9PDk1hZ+TjXtPW
owuDZ5MiTZ7fIwcsSLlhxPnrnNMfaXeUMIYsAoaTouVZtZcmHGkoMt9lSGUl4uwK
2T9pMnazxFQDIZUmISLwXKJItKgbry1w7ZnKu1+Yxe7r7hmbKy+ohuVMk3INxbOG
0ZljmnUC3Sab5QycCYbTmHkVSLAJYcbpwwoobzB2r0AKEl21WyEQj2IFXJGrxryU
Mw0hJSlBsAopcdgDlegHHcc+FXr0AeQtZV9JDAbSHzrO9cjxducumdA2BPkOGVRU
oPClNm4NGBP1TA7ND0LTYOGigBv1LCP/uaLr0bicOdIDT+aHtBv/PfOqORNFmZD6
b/cXbtt7xtOn3Kz/R5EbnOeu/fOQglCnkOzbDoJ1bN6SYk1pmTefEAUUAbR1ja6c
mRyLYJavXLNvVSB18EeLb8R0oooI3DE3sfAgxfUQXbyhPD10yrbSnZvaBxpLdVNW
YmKXp/gw52tC6avV5eA5VAzZEsKYi2qqd0PiH+5WeHzZjMicSi+A3dKz1xBlUCyO
iUKwE58MfgRN1JfI0QnKChcbB6mRUVFnqvd8YtowHKXta/Ewrx2yYsh7Y4AC5Bfu
17JEhePvhDFCYGWFSAcrFwj1hjenpJtHz/LJA2amWPm765NY1mpHwh95MR5g5FDc
paFCtieLLILM3A8xw0RF7/0xwnEUF3hkyG3WoXOVq5v0Va6L3GMCZNqblESXDoqm
qXZLg+1LbGXZJjPtpZYaCMJfsmBs5KwmmaSkF6gWYJQcayJARjQgur6AK3afSibp
76FiEc+vmEqBD+/zLu8EuyoT4YdEzL4DH2fa9YAKJhtLIiE0zs3iB78QzhU6duNm
aKFPihXQOHhWNqHm201o2VxkVNc/FKEMnJr1uavv8dBNFSmtMkuEutyV/oTXXUx2
LF54pgKa1rMQM0gcJdiyTG2F50j/OP+u+gM6wTKmX89ko1698fEi24zr5f0EP6xj
sNGhsTs01MAz5Tsdx2ZchNL97HCTleYkYOyTPgkQJluUAfgTi//8A3d1D1Xdo8gz
EkXHHLxRHPUpXz2kraCffJESLJMp7P4nW6GXZvJvvVJc0WW4CpNF0kmHnTHMwrBd
U2heXGmAzd8rj72L8SP2KsWErNkM0GKkJzCSGfeiFMNaXe/dC3Ri7PoIWF+GOvYt
Y54FSGMUarHvwfoW2EXGiLE5wbcKW2BW4OPKWqZIO1FnSYhoYIJXWO/z2Z+A2aqr
GvGuEUQO+tbyt7o83imeXwcYRZMqO7Om8bguzuNaBBXe26xmfMWztslPwb0WIhEs
FW3NVcTLhrq6psrwSbFqOIi/fropRLcGxeq4ZuhiDCbo3Y9ZrfEyRkiOmis2vXcj
6mxe/GfL9g3aICcS/nL6CAkgp/Z0/RUKvQEILx1tW7309iMpcb1BWiVUMbIXwMbn
1c47y7wBSrFASraox0You6raAMyShDvcqPkzPaRvwY7aLijhdQRcsRqAQ+dzt4M9
QmLyLLGeGASyt68SKVaXw3F2si2Pn+E9wbz+8HeovHGTc83Si/rc1MYtuo90187v
sRNa8oIKExgMw4YgZ8yZ8Mwq74mjcCK+Rfz7EiDHcQEDJC+hsN3y5ffHn2TV34Pe
CodClqW4ifeatf/8Wo1d+FslDQ89mH8EwRRdg46eRgQGVoUv5EQKyv0At23rW9L9
AeOGiSk1dbuTTF1n5zi3b8wX1qNF6lA+e5EUAFcbR9/xj/IwQ2KGBQovL1OTGkI3
gf4cy58mbCAQmVbsP4buie7kfKuWjB+MNZ6DGpdpgN0H19tVgaRUHE+sQiErNA+U
xZ4x1QlHssrxmYbfz5wJ1ihpShaggg5ZXs7mqPOHY4wXw0JOmNuf9Wo9o1cu+/1r
tl2yVd+24da4f7Y68y8CNGsbIRz9Up4L9fkP5gIcAUp5tPpxbkkVL3bDr8Cr1Yij
ZWHKvTmSrr7fgGviRsbIieOmWXqUqWBnOUce6DadbzhvEVWQ7CdloBR6LpGQQb+1
4NJSPO5lag+Qx/upGiZvY1+4G4UsURE87CVSWBqqU5J2K6QNiUGtL7AYCM4sD5F0
sWtvFlBzyq19xx3ad7j1PJ0SI27XX7jevyEpH7Qt4S0Y+18NdaHFKvV8cZ80+a+6
Q/bdxJZVjkxMrmApuVEfLbwM/Lztr99Qi3w9HrFYaw87adKO3KfOKzGS4TPO4a3j
HuhTrRCBUSNSzeDCAIOu+jNE4kir9iE8Fh0djxNS/WgSgXyjZCwA1ZWEGTjWvEVL
nTIr2lXzus5hJTlsQhRc2YYD5GBOSDO7lYyn4KkK3FPMBEjGHs8aO1ccbKr4bqwx
pPWUnyYmJXmXv0QAqHgPLjkvZeBurii/MahvmTD+vAkp9SznolTKq3yxBRb2qvt4
MHbiG2CLpgCVh1YqQEMubfqnBpoGHvGUyV6Vv4qKWSQKiqqKnWC+ZXohZziO67G8
Jp530rDSNptmk4eFKyrseERSMCyX0F7dlzmJ2e1UTS8HQRNb0DNaAmIG7eMbNB5g
opeaKZ6+lXMoNa5jP8QrcAYtR8pvQFvG2qpNIcEWhTuXVH3jq3XM2cm+BCuMBz42
WSJKssfKaGA1mvrhfj4CuATWwio3kQ9wsah9YA1VcI7tqy1WDM7jTxoiekMRtlp+
kkVPchVm93UcCHJ82zFBM0SK9tkpgdke800PtJuLc1K62siTt/64JmqpjVlUuOcP
ELUgWPWJ2b7SluJ6lA4/YmTVLYRdf5Y16Bps4B/C73wjW1zwixqYiAxYM21r6vh1
cXyavXBlKjfJ+jg2CRHFN17U2b3u1adLzo5gS1HeAcyfD4in9gZNCIBIT1tiXz8n
YM/iMeFgvaHXHvB+v7TqrQ5LADXgHj1QsEg5QHTQIt8AFkSlHMCrW03ml4b/V/+X
pq85OAGcu3OR04dRDIehPmSmf6ijjeQrK7Rf1cBGs0tLkZbc4ETPWaT4dFQQD9Ka
qjQrYmPlp/yry+pC2tQDZ4iNGAfj/yirRzR6f+WlxC7apmKwQOgVbiRFM8V/dion
g113u6vk/SzINj9Hv5hiuARbb8pwfFajcK2H5xpwpbKamPY67cyEyvGy3KBGKQLd
swHIzM85/NLkfCnFE8ZJ5w08bUF53F5t3a2F28gWiL8hBmohRWnuxFtvZV9nka8e
PWGLcuW5sCovuGR2+naOyRzBNk0qWdgSKWXw1nJdGHR+fBirYqkPGoVNhwXZWhSB
+nR5u/ENo4ScYw+T1gPkhidxKK52s8lR5Txtv76MhIUS1drinXrgv23RYAaOV2KS
6+IHdYkAaR9nhstMvCb2IWAIbaM/SsyfaHHLzcDox7r643rG1AETqLSwywJQtDi+
0itatAiJGgr2MZGpx2l2layqInBdPFXUZSJLcznUhW0XpwKEmRoacr8KGwAZWjWW
C/MREG8N2ArsJDlAdqLe/n6e9Y6O6LjzX4TgtOHOcqd+CyfJ09A0zYTGNiRTh5ER
QU4YkKZlC6Lb9UUriY0Bw9Gej7i6iISuQkgrAdLY0WOBs4L1MTciO60z8ZyeN8hq
aJiBs5xJG+pmjhdAb6pmN1roSL29+f2j4Yt3UEvfbzlJISxcSW1OzBPX2H0Jqe/p
pJ+5T36mxFsKMbv7bvg5Wx1vjXHiBq/jU59sJa0CIIAXPkLJbbyzr5YgCZDcCdRC
tdW85WiBlxRf0R04rezJ2/b+WJtn7pJAx3KdqvvI+C58CLeqU7YnjCe0MDng25mr
Jr27vQhrV3Av9PvnSgVc1fqKcnprVhQV2yElZtn8IPGCnUgxeel3Jt19PkNJ1v/v
B0c8jktCpUxMKIQ/cMND3eE80LIRkBkd4Y+wsFjwO4RZhFEL09Mut9QdqHahhhs5
0u98mywG/hfeQCg5Jf5rvAYUQSOR5mVjuvyICt+KLCtgTk0j2mbw0NVzfvvJy97r
GDuOuH09Qe/wFTnwCVerB4PT3DDJ7Ayl4RutwGX3U98K5sSiPoq3UP1pjWwOIROa
cprG52GFOq7LcZdB7dsYk9JZi4kPlPY3T43cpXPx7aZEGg3FZdWLXGyFZPI4S5gm
/3CsgMW5/zcjeLWnS7sVncRQyRX7rAq2/Q1Kb4l2cow+8o4/Wg/uv9MigKcMbscD
r/ePXjBamJXCNQWBxlClZ6X+gIwyZ1arsGyEV4X507usRhHdS7/XNQ9SAGKTkioD
vEuNDh65mPmo8kZLQlnIo9WEYtMPF0X3n2Z5mUhZ4CrXH5eiLWUY98dWLVCeSSax
6xNKxHXWKUgzNaTOj1v5z1C1YbgvRvAGojVf/dAhdhz2Vokob/6j0v+2nGBwA+mG
5Yb968t6bxkCi+6bneMyYzkehF252fMkxeqGsK+V4UiuQicdTKqZxEtu9GHUtwQc
ymROc5pAzk3UPt//V0o7gOsmFEkpVM16ViJqGvPeQY4cJchlsAQoB2+ABvBPrWVX
oEY48v5d2au8cT07Oz117fNCklvyvTlrcklih46biH8T8/tqu4yd3AE//BZDbqu/
EAgfVngNM3DXWBdo9Rj3iFOLuG+RlkdALcWH9DldgCQzClZZqkqFwPhsdvSu9wN9
HBC5MFFTvEXUD1oTH+183WCLQcrNmld4tBd6m3TzrOT44bCbxRblPOEe41laoFBo
4le680rfVDhpKqc9W5TDPxPopPEanh5Ae5r5/+03eb9zKZTeN8zKMm3i1y7wReaN
iYkw2tCAHzZQdYdQAnSPbiovUYTRuL7ql8U2spCjuqN1bETjX/l61NNxGV1rw52v
rHlnr+qRNezTI8eQUMwhO7kPFfhtiPB1PI9fZ2Z5JPM0zRFvgVe27RjDdCSl4p3Y
2VmqxNsbakCn/y46dkCVm6LOR6F/yiMxozf82l5qS7mD82PzXl7ysL8Tjj7e8MZo
AXsbd4FINmxTT3uCgsUAcxwAX/apnw5SH7CCW0qQnNdIyjo8/LDKKRwRXGcVyY0h
mirvDxuKj10XvMJM/0li8fsUjiiflTBr1vTMTk0ZhHz7+0pjYTx4SluEYbIp5/WK
Mx/U36KRuhKBeQGTawxHNHEcZPSLFCuwYuoKwIy9zR3oaG6zTrpkSwYQ4t32gxGU
KDfAoohj3AYi7wZwDrCn5XjfaIVGkmHCJbaKfD8eaLmhdNy+Ztiv/jY8U+CfvJE7
amzg3E/RI9aJe+Dhw1JMy+nwy00YuThA7IViqcTMQ6aRZe2xUBg7ulc9wgw2vxhV
J/glBp+dnsk8QrIRWcaPx8SJewDTig534aZs/mdpwfgluPNrjHmnCOSubPOvPdgJ
YbWUfS69wnAb5lZoiJJOXoaRY/iMi6IeGYBDVxVhjg+EiQE5IG8wLFA6tmNCEIRa
OSiDEqivFXC+V0JNsMWk1xUmSoZW3OxInmRr6DLZYkFs5KCoDmep7MRtvaDmNq0r
f7EwVZZ8uzmroEhd2KwnUq4+BchH5VuoMgzjdwhmnxoU7SBR5YImFh/wgj7zgwcM
R6vi6xuIcvJc1A42XWliRwkW9XfAoeQqB+L/BKJPXDhlzYoJZeF6pWTaCgUJCCtg
BqEWz5BypgUR4S3CsUUALPcMrlbKRI1IIogeik5zlPmos5ZBPbV8+PiXQyTu6mup
8FYh5QBH2UZ4YwmAG3BfPygvjcCpf1rLVX6qjIjAPo+NJIA+hn3Dur2GKye3fiv5
b3vaOUY3/r/EFN+/An/v9VMAwumsX3TZpC8tIrAWRC+i2M+A4mYsdTlnzQ1LMsj2
K9cTPDLk50mhQ5mMC3CqpQ+4xf7ZYbKqI0fRAe9FqvOQwQ5wzY26LO3GyCmAQVV6
sQJBinQo3VjEP368RdqzppkcbZSwczOd1CLyH+DQFL8+4hB24vh2p5p+Awbk04HA
sv5D1Gr5oD/Ekwj9oKOzB1JnY1lWHyql7rKwztkF2mjDC/wjgoZFJaPobDXlxfOx
j5iXfE96z6qiVdzQxMwJ2eZ4lK7ypE4rbOdmgZ77FZ+ijYLWDPVHGcHV4zmJRAt+
1EpuZha+5FongdwOLt4AlSjH947tfuy/tY4LPdRAASiohNFKD7DeiiGOp11/O2m8
rKF/XkSTGHN17mmInNn1B21AOS7D8xFyvyl0LY4tKB4JKKlmYayBFqi3JGPm1I4J
gOtHfsoUmr50aO452OaD4otHGvElG4pkY+9Ylvjdc5bh5+HHKCdC+Scf0NVYw7w/
L0sjenxVhoE2oKc5JLBxG1UQlgRXuCBxKQDk4ZsewI8chMx87b83/Jvof0wQCYCU
/m8Sl3RF+9014STTLQ5DLcgAX4/H5VCgoqI4VO36REgOuIusmavHzeI9+AKaG6rL
TCm/vy1Kbp5DuQDkuKV1s6d1qr4NAc8kr4qSu7AABwhjmGIYqiv9N6GONjbW1bdR
usJWhsDW0mG5y5d95sRpaI9Oj5VgzIieCVwueCNmvZ34qaBbCIIpykDyZLQYS0jN
6gsVbaYa9YHVWrca4GLZKYE3L2IuuWSaaPM4FzrXdD6EDyzFJewzPXdaEgLoBEJq
n+NG8SOwsq18q5sioGTaZQHP5rurasT58/35Fnxf6aQhTrt/JQc7nstD9t9hyOq1
bHATRtcKThrrC+xULouaUnVYmtuIzIATzJJlzU2MWoF/QxsUPzJ6fMaPXSnS0TLP
grIB9II9bvCHX5TNvuIs0wPvDjH00x+FgPRNxjNR2Vyw8PI8aPlYxL9h9RVNqhDP
DaMLub+LZrBJjTWducQdhJnJFKNYAwyK+kYjTIk4uqG6RIPv+T6WcBy4cMw9mXmI
dieedhPDYXvckAmwGDtDOpU4zkJjNJJspoikRKYuWTLImLwsAFBKFikcBcK4XJDU
gwYAT4BwD6wwze4OIA0vgpsIX7iRmmlTxfIcY4bUPi/djH/aU/OZq1wgM0Ta4o8K
t7BVb0ocQCAQ7pTjz1GPAPJGSv3/L12pa7ix0/6cRboHdUY5OuTyQebLqZDXNlNb
3C1luCl36SLBG4MTQOACPbIMJ3xn4WYRVMBUJLPSM3w8edgt0ugSLS2L/9DP9W5e
88SIkxDShOOqFIegFZ/NQkBYNNBlspLEgap91345JoFfSotz5bBoBVz0r6t+GSCn
S8eJQ1LUjt3Df+7zdwRanUAOLBX2ROnumFhQRAUnlX7n5SAusrnSENKMrZulz4kE
/HiJXVjgE2jAuoXSsTVwdHaIRsnpClvYEy+5GYTw5QrO8k4mhYruOYzqtPDiJP5z
shq4IwdeQEPupcB5DMVQ5AGs4yey96SXCJSz/bj+LofUXqX3xsX6x+JP4arlsK7X
9d9Q4oKAX07rz4yj3SKymH8MTnTMXS9C0qhL1TzkXZQ8ZC3SeTEUHNSj3SvflGMy
c5f2imHDpCT+5wQxPDbZ0VOK8siCp3wcikZYOmNTOMhgpSk5urU5Gy1JIqh+4uCK
cXd2XshA4/fMIdJvcnprd6rGfJHd1Exl/Y9O7oUjRBK/kpq82Vg2GATxdWKM4m8M
tPYpt2XgzuRTqe7LkZW/WeUCfQhhAMtr6MqTbb8xje5ncQ8h95HLI1KyRiZMarf0
BOdAY82LUMWuKgRk3Vr6SHPQ2CITQlXH6/LjtYIHZ4vGjgtFO3Jvjk3OjWjDKiig
M9rpDr3MbJiPc/JcKPaP81dGe4TBFQEfkZHvrt+OksLW+l9NKOWJpCsgroaDKD/X
4kmdM4EXr+xwPwPKckBYaj61tq600WXqIcB3mC0RPzi5QUnw2SirnVMcLQI39DDz
mmnZwq2P7dAV2IhSIAzNjt67D0lrVl8MEh63q/0eFoGoeuMBVoz1WG09+xO3WYxg
cy8nqEfhb05zWrPBNTuCMvFSdYDF+/BXc18Sf82FAcspsl5fRk0Ii/MLFYkjdMj/
U4hofjk3JI/oY2y92UN625Jleutl6Z4dIXtj2HlP/l/zeIGDA0jCNzTAyu4M72ES
8CCG94pCrrqnnvgkEJyf11iTDH5WNa2E35rS7+knoHiG42z2SkH0Wgeu7iZ9mPOD
o7O9pagSM905/+GVz0cgcUS/Vp9hdD1mXdp6ObKNCoL56QhinTkZEcPVZjJrY9IM
lzqPT4XYlpD3LxYZsmSE3Rwox45l9VT3a87/+6ZAIMJShzXPrJliqSUycFqwbzZh
HtonFkvaY5Qo52ogHpowrhODljQnU1H5Ra2bI4ferV178zIjTOH2KMLl6l+ZNB9F
Gqjs/r097FeUGOsOXjtg2e2VTV+oZILFY8VzNBqfivJICPLS6sHcz3mnnLhmMzDF
gnYAcQdNJRcpdhbrhUEAJAOzTsUp/JNMREFKVizzVKlheNHjimobRE/XW0Fg+Ukl
vry5j7tKSzpHzoXJC3YFU0tEXwmdC9FAd6EPSiw1CyKSL0XgJirRJ3/Y517JwbJZ
dgJHYQWKDBzPUCSXnxJD8pnTyUHWjou1pc7QngCi1aSbe8ODVckn7MHzBjgRpCCU
OL3qkQgbZ5z1zB7ks27jFiXGR6Q6yhx75LdNXNLPxLiRzjRKLWV8Q4EDe/SqkW8q
k5tIWYRapWqRFzwg5+rvgpHMTPpwDeiZL/fHVt3CDDxM9/6KGIHTWEZwjNW5vrTj
D3jWSm4qkRywX0586z/2IPoAokAqiiGnKFwRUNi0NvpUJ+WajEhbyuSKxutFUxg6
0o85UadMMzV+HnS8tKO5lImUZIENC0R1ZmF6msAFvBSm1zD+d5fVKjox1lntaYBv
oIxCI6EzNm+vsF6XvJLIxtgGONAJXCM7ApMyHeeQUoqo1byNT6uG04EDughiNdm0
pQJRScvJxuWqxk+lY+DPFjw881FA+I8uJzR9i4TvCKLzkssJ4BOs9XYGWM/rLEJW
xD6CuXXdoBl7gOrgJgy0+NSFi1yBhJZK2nul4A1zQA4pNaJwCE4bE1scg8eRIjiT
pHiJXG2uSkCmlOrixDs+wdacPyN/wmlvIqDTiSDFYFyiVsun0zgaUcBsBxN4ECET
rrkZCv/d4PpdO++YF5Wr9mZqZgUUnTGpOmzFKqrE9LBgIrS4E/IR1qEwcCl0Hzi1
BLS0zU7eAo6DiLKb0PfvCtyBVYC5SWUr8Y94vPuJwvFmgoeNb1tK19liREoHZOdQ
b1E07D8Nex4bQBX1kCJkP8WM1Jf9YWA+Pw9Q+rzFdOa7nSHlLTgHpZkVj70ZVgsg
JMpnfWqNJUs3itJRecs9JlTcpnWMjQ4TqS+LfYqg0fpUE5fOBan+Y5hRq1OqixLR
A9EFFy+vvyzCWHRWk6STayJOHt0hqZnMoV6/ZKt7f/1S/vr3kLNUhzP/yHS+dZlO
BV8LohZVD4fQGIhdEyy+aJZQs337hZbOfdaZB04w+mi3lwQlcoziKedPF0+L+ITI
YYuG751NsRa6R129A7msf02w44tNETMBiwstnUjPFE6jbrupunAXFOEfzNR/Eob3
YsBCNkKmVZAjcsHHfl2Z8qxe+2/jwo6WRuRkCHaAfkzUY5k1ijvMwR+Dp22UsTeA
Xc3rMyTIytjsKNUpy44J8NkeWilrQNJh3lKf1+lBK/9Qu5QcZrFVbYhTrqcM9I9K
k+pQFKOxAjKHftO2G+wVNUuDUgCmhrVtD60EyvMokiSKKdhPav3JryAOMlVAhcuo
pfGh7pspI9GfoTzDxTCqfKM7fZNgf1aLzwAv/EbDZ13qk/dz44Yf2uDDrNeZ89Gi
lgoqt4aSNkjacDP3+1Hkay1CkCu3lt5WgAaUIdakY2pu6egyiElV3y1v1tyayKF/
ItgeZu+1leGJzFac9spxLXGJe3oTWxSUkfABszfBtKqTmNuMc3NNbSZ9uJxXrgWC
5RzuzhSwk/ntHKxJ7rgUl8V7LcXjdI5MOnBveGYz8uDDsKfVsQUTIb/ORBZri445
n99EXsPe1rKVvfoxEO0kJAz0SOHISjs9zNhz8tNrG4rSkG3G6qSSHHzbsvfnIP/D
9FLZKty5CD5Hks9rlF/1INmlwrQ/daEzsIjP4lHWUo5fFmMOCRm2ARsRa9lUq69s
KHpeDTPanJqP2pR95zrlBO2y0kEziJ6O2USKxppnlZ9fvMs4j+ybCiKIeBONu93e
hpQOKb3nwdu6UIvH3MngqQ2RBhNjQ+a3w68fNopl6CAVEvQJYE7wGoylQM1RA/+N
/INjxqqjxaV/gOW/6z1OLp0eZu2MLfZK7R6apfn4nu6YpRGEMzZQFW83ZojjX7ma
950E9LOq2xF468kjq0FbLdWyrlV803h0dPY4PwdpbVeAAS2W8dhK2xNtgU1BMETw
83FH8KW5f9dY2vk7lpSdPjlIAMp/ILes4O5dWfc6Bnv/a7AVR7IQkIzXipRUm0wj
xKtjj86o/ReZ6GgRP5SLOh8ybAWFYn5E2nmqtdzhXm4Iccb5k4uGkSGijDgaOcKl
EiFET9iDV1LQ7K+ANXCkP5NPQzKE874yoFo/4jfKRWlNNhsMRcvLP0TNM7SYTB2P
xqb1RGdBOuK177Pf7R2/02gvyV53iAf73fyxva4AsZgN3G39B0vOPqcJAwZZstCG
Ef7UwXRx0jZB5S2vwLmEeeo9VfJpvuljohZK0GuEGlr+UaBWxU/ikzU/fwY0/Ypy
xn/sJ2thBr5MLwvqRkTzgXRqXs2+G/EsQtCf2NX+Mz33L1rOx+QPGBE1BSsMOVH8
bW2E1jJaszx+sfp+R+gxiBSCUn3YaEtKbUPTPyiSnXclD0+vLCrIsat+GMkjwOJV
US395kMSGjcTXem/iTsKkMLKWiu3OEHq+Q/I9ushR8ad3cimaqEnMoeJK0rDn0cE
KDfoebRTEj1dsBwZPbq9e2BZO3eFthjLGrNQNrKhx/H7RdBLa9mgCpeSZVYCcpwe
30WIwM51GONdFKnipp/b/56acE+cjbmpfLADO1CLGkyhaXXvm+5Ce/zrISva3dU9
fOGWKQF4Qk05I2eryEpcjP5pZWV1PfxvTsEsUgoCKsPl0uMTzKUbvsxgZAzk7m/Y
QZ6e8Qu47+Ct0sY087A5G5FeQUHY2QJjKoa5Mqrq2j/a+yBICK/mny72VAakEniN
PG/PjeKtIDXe8PE+4ZiqNp6U7tD/XRCjixYNVu45ktPixhNc6fVnSONF0jVy4+eF
P5nt8r64fIZRcanO07DCH8BvcGdx9hoS3ZGF+MZPPjmCG1VdOfUCNz7yAMmgmGHC
Ho8RNXO5I5sIQRc5I1xP9LDy2PRQ12Q9vHCrG3sW65hYS/QAQ8mg4vYROnwBNHfb
dEQA97vDmJHszFiXJKxfncnT8qcOjvY4Y6hQzSqJ+dgLah1xJVeEvd6rLW3w5yrU
paaFSZsZhe1Cn78C1C3tgivhQB/ofERxQtEd57aPBKkiXg7EhHlfHlzfUQkYOIn8
Bt5wbMRKN5CVzH5hPSSrN1ZkB/o1sp4DyFLftq3JnRsWid7fgIa/+PrKUr2wFTXR
Af1YQChrvtxhR7o5MpzgDMaStiPBwwzqONCwOnpBev/kvbPU7Jybmrof3FD1t8f3
d0zVfINUhpnyRyozExYdYcSZHNID+6NnmO4MiqXsBEWHpKdNXWh44az3ezoGfByB
LxeawqPzvFo6MgVPMp3h9xfv7+zQSmnry/jb7HC0wHqkltl6q1BPmeCKuwK4OgP0
1T+L37PY1z/AGxbCZXbyFTqcGys0fDUJqZo+Czvvn2dWhggsy56N3pva+RJjZ5lm
dSF0sYl19mpXSWZ7KgtX1goQh0LOpjsvi/PXX1MCU/KvMbmUOjBclPyah3AgFWrT
CEKhU6eWqu1RuZq2XjVwBi7ZQUvQLdrge1st4ZdDpjw+643UhyctE84T141AhOda
bNPDSEedrH0GxZgBRsC2RNkIRt5bW09/V+8OpsfNV0o6IDNb07WCTfj4hu9GvUkS
RBniEUzSiwOocCZLvD/JeoHi576oqn9dwCWvZHm7NviV5uFjezLNitz2cD+nOKxc
qT2vt8RfzGrT/Qj+TT8FamkwjswLf689P63W8Gl3smr8JNMQ8Fyt0sOwkgO//QjS
ole+vJgnFZWm1PZdTYvx7OtZDTlJNkdOZe1PzB8ehJg2F5HHXutyQ9tU04m022Bq
+mne/8+VpRYQpG4JQKwFIV6OGNRlE1l/EPwKBghlXwqSbVkytfs69VRUJjDKSffW
ZsMG7QDRQAMn+EGYWMyCI8n4l8PK/PdJFILxEnpZ6sb1MTu9K5WLa8IzOOM+aGGx
qgEFXNmkeOa4CmRmioD1MOyZ7hfHIvpUZioRif1NwayJPS07DM0EALsJnpN+yAHo
XieValTubAEOsewV2v9FuygFMoJjbmkhiE1SYocCR8OoKpKJABvbcu0vc6RKEK90
OpyRFerWXld7qBGXenwVJ4zQtyCVgLRAtTMRS4vlFU0V+JZjMunvGwGJWZpa/niw
wR/8H338zGz4iyQuI/aplXsZHtinJRvc7SWgd6NmgltxtGlKa4wyK7PXKx2m6Pja
/uJ7tqOJ3NWtF+4/ayqNxq65UKRMh18fNoY8p2bLTRRe+sUOSKoKmwrxfEqboRTx
hT83dsLhdzI7Jor51vRcfBw1Rlia937jJlXPc8zDBQGFOrUgjaB4E344OE1Jg/HT
SpSDxkuIqZoRRrS4t+LFl+/RlyW9+p06Vv9zh/1LFrRrCSgm+7r97+Y8ir/4ByO5
SVWJ4L5r8TLB4zErMs0W/dIAN+GmtewVNWjzUe3MsGiVf2+v4tPgCfO4jz3Yq4wY
6OoEICiV83oiWNxxa4C16JvHGLjkpr5BTNky5IAvAwKbPHlBtBewJ/C/ntIqQpN7
xvNB/S5jXIkg+p/Il0MSylIlv5bJpxTLzB02ewJ4SS10iAIVljRoToB1q79fO1Pb
4fTDsC0PfJxB1c244TKpVMjRRJPfQ9PoL28Ep+YnsEDcwnd18lSbZfrafnRjYjrx
PreGOyRwH1rAJNme2jJqp1d5ooPvQ6BdAEfe04ibzVumSTZDTnsFi7fy419lwl9d
hz2C+OhRxIkJwm4vedhEYW11d95MD/sQvFdT6AzV4xh7Hic29XbRaG9NdQ1aISMU
CGUzAcEzqJBmiZz6Du3zAdlks3C5hE241a0TKv0jiudeiD/HiaeFjpo2AjckABwe
rqCjjTr72BJJOBIw7QFc65CphcLC6RbMuuVmL6oER6svZqBjoTXJy2RBFkR42gL3
jhpiCXA9Cq7SgZ5pgiGJIXq4dOewO5jO92zHXQjYitbOcJtR72n44bWA7a39aI0b
b6Q6l/Jlq6jcHGXstdnNHE76GpFsO0n4At0w3e5vWXcvKXEK9zNFTJWXBQrr2Yo5
/38JjxDyE4jPPo3YxaIadud1cxVxmqvPBqiytj8+baQ/1dSRjlu0OtQlVTBq9VpB
yZcPH7sUGm37P+kZRnq8pw4+4tVeN9fmOdN+7n83Jd44BRtyAsLn5wW0YqGCKFw7
2YRWcdRb3XR+Kq5NxAbeV7hDUUv+ABxXqV4AlhxOvFeftzqLiDB6rPUrZaqkYQb+
kHnJvnRjUJKVjaKLzAimcru2kbvRTrn6pioY3s10IoOnNSDlxsOAsxfirY+v+im+
jQofxWH8DN5RCeNy7UI9D+1jLdIVkOPaw4cXhGi0Goe46NeZbC0HSseVNXxjUQmY
OWLwezFR6WaPv5QDZ0utZEoZNc5dirskmOki4Pjwy/6bw7b1qur3uLkrpvZ05F8O
sZPnd5ZjEHbBiJMQA2zQ3KaRstFoANXmOG7auo60DJG0NFzt1olhNFiTyvT1KL26
4NkzgWtllGVVf6inYLw/Y38C5a6d/Tm5B/Shh1dZziEpEg8l+kpJ1owRXCDLUVEa
QpPqg7f2k6qKINAU2gs56xPk+v7TcabFLyIbHYp/EPM4IFzwZHkffBGA6lHk1c/8
/mBTW2JZng0PG6Ox5mMbLwU5GbcxUZww1paafN+KgtvYTkPcOK8KxSTJD7iPY+TM
65On2ieSmGbcebjJd8W9J8RlXIBSsHGy/15Er6sUfqs/C3hikq4scDZjm63s1MV8
gwYLMhHaBChK8cc2nFLfnxzZOW2/Dy8wAluIN0n7GclPKyTypYPdpxim9LwGk9B4
9PgEi5gj70pLRreTKv2aq7rJL6buhp87p5fYjl7f8gLbISZ6UmBjGQdZ6qkGDmV9
GgUJF6Kwx8GcpKzzHXJSywGUWjtXyu+VkR1Ys6Pkhu+602WTSgBKoPkKIYRf+y15
juZ+YyWmODhlTyh3NowNb/0kPDinZmSiJdoWVznk+OYIgGlgCq9I3RCvCiyRlahO
Wj95YAwsPNPYJOEEdQCHROz65eh0HFuBpqxBfy0x4J2X/h8Z3UmzqEyUIdgVBn8z
Abzy5NzF9Kvu9OqGik98iaOcqLQujcHWFRSSHTeJrkoXNjhYoD+jZKj6Uni8kTEH
IdlsEbo+mfjfVZ1nqAyd9EDCdrYASrTK91/PiVTo3Kmx/2V2BtPGEUIBglT7MfD/
pApsdi/ky5UIIM5qFP9gAdohi+ABGj4qQyePHETTM4OmI4VIUz0FZ0HfpCOlrmw4
bjrzEgLLiInNiQU25/JwOu5TEy3Show5SfVjk9I5dYb1hHgQ6T8FDOmjv+z9q2J+
Bi9mRiSDJ54Mvxdl0UCzrGxEU3XFxoK9E3+5OjtvZnA/56/g3+nxvxQ1d8d8/5JL
1nCmxqkM4sZRC3MHnqzjx4HsCphyHjQ2FVTaug1NGx4ws9ErI/sqUMQRHsYVVUNx
SBZjvSGparXYSjZLfSSz54rY0h8jL40yHk5QnIl510SoxpH8bDHEc31YCeYszRRf
trEKiB1PD5f2wT87I5SehxIiwIkUHLnjTgjiVWfjeSr4afLb4ITdLMgZfE8i0nu4
/q5RzwydxNePWZWX0/6SkZoWalfP+5OfU8Zsodq8BCzvF3uGIz350pUd5QRvAcL7
Gh6ILGtMgT9qPX8SDuytF6cO7C3hmCInSgz8ROibyVTyq/wV31khrNpf5IRlkDpZ
tBdORZgdUqgDp6ipqHI/IddEpO2TDSlJvApUNle37EQSd1O8GmcvCVaZevFmEai2
6nbBZo8osHsPnLr8L6EVxEf62Wf8PKb3muN1tE5Ot7GnGP8IYmM92IuUrwC0ofcN
/cI6XDGAgf8+yOYW0LGEHeL+LRi+vxMjAVqxgycKZRFawfycsKGbdd3qSaGpTiql
TeUX3aXmTSQYaU1/46lcE1OtMeJBW9bNK4V3r2QvdBPuUEArQx7jMpeZ6uw795EC
Nnswd96Z3EhI5kfzGez0jyw4jGgbSSSokX1LogBkB5dSpBCGa/rLa6CjBfmS+fpw
jV4cUi86Zw/v5Xk29cHrLU28rSw+yVEi3CUQLrfA302dVdNYb3956xSBuYmu9M67
E3R0vyJ+FBc6CIodEqhubdQ03llGTF55aXoTAFkbOkI9FUjb75ZZvdPF96cnonTj
QHsPeHGyJeJpUgsoI9k/Jv10tULurXNSH8tGAnnyDjRJjf5WJedaTPIxy3cVLDog
MDA8bOosiNr2K37c8p2P+WVUw8P+6w2ZWaKmXep3sjintle76zI6DQrCrrerGNvK
MWbC58YXC2NxCd4tI8vMSRyK8j337XEE6rOb3KAoSk6K3OhmnKlS9GpQARy/vRLg
Dwt2Wi6CDRgo4FTN3zKrHuPqaGeWSjQqxfYyEz+1ZJAaQAvfsPwQuob8FTW/3PFg
JhCTW79hOISF+0J5fKiZ92T6XY5U3wll8YefbgUoTPAkfomOpQgiCICA4kU1yS8V
GQiDJc2ukDpnEGVwA1T3vv4rmPnZnV6P3Qn4JLKpYcn9NIjiKH0eyrDNH08fl6Rc
xSpYjsPI46Q22RkrzndPP7rAMzhokrEaFDLRcRCHqHkLK+lkVCsPRpZvbBhsGrLk
mQlcnNx7Y01+i7yAZAmWoGd/t0zQDmvP2l1VCndjTc/ng1NmdLxMnzqbgBxFEyqE
b+zoafHLp11O6GRT/jPr1OEeVn3d41AZnABiTkpemAcGKgFoPoK43//nbjZO6ImM
SE11qJx+kJQTQHBb4yImHZKusVDZrPV3FyulmZojx5raZ+UWN6KuiTlpQLkir3M8
0RoCzQAzXoantrwff7jhq9KnHpFqMIXuJmhI+h4Pz2TXUTmBXR7M6GSwuZoz4JUa
Szlv2x0nzQwJ9JZkDFiBVVikoYJtF1z31xgOelvxBfdPA2D++4HVRU/6rAdu1Zs7
NIbYdhK9b0YEwu/oowywY7a1rJHP8pchqnpyzPMkxHPGyA4nZYnQliGv60yDXRFd
ya7pctbAF3i8ipnC0ddNy+MjJU5/q3oyXml6Zy3OWK8YUXmqjG9rKYpVETiK5WbT
c51HnhOACyFmjDYLEv78akVQhJ4sO/ImJMZyhdQ/CYoP78pGm4JOURU3CX+WPJFU
2vkRYK9syD5cfmnMJKeuv/cSazAaSiAWc4mYdTOdUI6NYS+Sc5jyFhzLeojoTXFa
6W0rZsCRpliWsI+I+LbqqTM++hoT/Zr8InBZAGpAsVoWnkbjRjsMoO5dhzMo3ZmM
Eh+uPRKyvfTcRT44r/swzPU/I9tBJKUbNEvglbL9brmSYC8v94S0bUcQxQ0i1a4R
zk7pMgQZK0/DR20zlD1cVcDDoZ45H5r3c0ZC2mMDHkfLbbIZAEFPHki4CD/ZPoFX
i8lWxNnTPmtuHkBmWgcCyRwmYigONJoSFqtOth0iLnF/URQ83PbsbbJeLRUBEdko
hJz7VuGb6+2T+qnkM8qcu0/QhPkIsKBQu8sZ32SL37P8Jwc91qUZl8PIMgZke0Yp
ERc76jos1LttzXohvX/aLXx6YOEAGaecFQ8PdX8V09wEGUy8zsblhIl5ZVeAdI7w
MdFT35hclkjhrne+/83yC4Ccx6zBrciizrogk2+TzI58ze1jhqX+eXRBjIWMpSWn
3Z7Q6o2oWALI3YvFcw5eUb9hWX7/T01M5XewRsu46oTWPuIwVpuPUcC68XUdphHk
gTafELcvgNQYKyt1IV/4bkIsAyTl8g5+T2byjEd+Iw0z/VmK4N6ByBF9WZaKGlzD
xFeJSu/K0RcelOMLA6BxuID06rCtFGrFJTZNWo6sA+lBCsE4vgMECXHrOc4XL+11
hFzX8nX+7Tr6WbL1IDZQp7Y8sGSB/oSdz9zA/xnVCuYmq7/pHsEuGWi4LwdTbW68
FU88uXKDtBsRqSaAesKOVKO1McG1y8N3HSfxyrJYXJnzHxGP2mPWypOHLHTPClzq
2V7C0rXbTQTJNfyP7kXYypDP7Y2/B8nnH2oJKULY7U4pamX06JGjKy4m3jRHIW+V
xkomeddWWUv5/WgHFVzJRm9PlG13sQ+IbCTeHaQUxdkreuCwxd6fdY+2yxaXgjsx
sqFD9f1pjLm6BqsxlnAV6MRgL/wGSidrD5IiSvDz/oYzU4H5azPUmpXAqU8u0TY6
CDzqCbssg2vTfM57C8UvU7gYtxcReBPTAnIgCyG+AP2a1OkYm3qDCvXkxc2DgpDE
y6plxvyyYD/rfjkT08TpA08hNx/1Nk/JToOAiDCVOMX5iJx3fNhda90arMkPufDL
rePWDDgWtYD23uBN+gnEDkdYjtpvwnsvDI3iR0IAVrlgMqKKwuDBAv3k/NO5qjtw
oChuav+uiBrPjckJjRuE0edgdb2INQK6sp5K1Emd4G5fSEV7L5uCz0jp0dXHW3Vb
gUDqh13DRjaCZyIp9DBT4AA3w1Zs+3VgSEcdYuMp3jCCY+IROwHnUBTXas26smFZ
SudS5o1bWOLxc9mSkS8K09hcz1fNR8uqG4EIn1FKc5zdXnO1t9NR5IhybeHgRW5H
iEhfBB2ddSI837YAmdL2OqrjaUm+feU88GhTySRlA7DH1k/YECqlgplyBa2zaaci
1dpik18Tx5JqDJpIbIYJpkjvndgEQr2Ns6okKE2CODjbQSGdl1j7RgAU+vSwTulf
U3bLFvXtR5d0fMKiIIiwElFUKJwzMR5frYIycTczgb/qDAV31Wr76MrNrcpYEyt4
d4LCBbSLuoOhkt2VMqpKbSwHyu7a4b0ohc1YolNsF5tVjMgLLuGa+sQJL3LWQxWr
8/RBL2Q8Lf4e6RpI0EDDoFrWRcirvz5hCEdHNvby0mDZMu7H9aMVdIzKrhKCrIay
tzeMtFWdrpVJX2Bx6m4tGxBcqRhcfLCEQJbzWfxjXQOtzBJmq0oF7NlZ8OmJklFL
J3M6LNw+PnrtXSFh4/YCx6MzqHzFz9PndlQUN1zzPQQXNlrYygKkJJa2gIgAblto
JKd5LM+KbeylALblBWyVlufLDt/m6InWXslIEyDQwR9VgQVx0MCroTwFfGHgYAHb
kjAgcqqZ4uLhUiAd7ebLF62l855xHEpJcRNv+N6b38ZdIHBZ328J7rwARuf+6ani
GDcj5HsoFsyLgUvrtQMOjzBAxb8yceccc+M1hXUaGxQ17J0gPb1YEVX5oTOfzQuf
uJ3hVriejPbazbluvicTvXQJVHEpKPcdXV9D/kO/WW76wuTd6joGeuRu+lu3bhDB
PAZn2xpPZ7IF+E63M7d/cl0gO2iz7Okh+Ac88B6AoyB0fuQQFRc0K9Gimm/9KG7W
dgqdTxovW87RO8Y+3jXoJB70m5uTHq7pJrI7hLAfxtIwxbNa6bnw/YcvPRFO5Yo8
Rx9ErKm9Uv1VjckBQJLGS9CzQcTD21iAuLI15PWwOvadVxkslu47xcM4a22MpCTu
IbrUZxwRiQ0O0rgD8/Xk4HuSotBrVwRNxqaHq03vA68xR/eCd6VmWQhHaGKrtIOl
wS/oF1z+LS6ruGIoGtqYIkhOOdUArM4ILwEpDlQC8O4jlgT7/62jJ+5pe0vfhuNq
tkpZy2n8vpSjcCjcvcVlE9iawsRubX3qVpWtao/4OJsM/KGSggmLCEAQzrfuDgfX
z7we4d/kS1qrrbG8Maa01Od3qbJ+4G05kDUrPNGyU5bOan5fp5eYHU0KIspSJdyP
1ncp77gFsTsV7zaVq0+9VXcXMNeczfIkKJrKU7xzg8YgMeBcqdUCyGPDRpYSGbmG
OR4sSsuyVUe2c2cP0Vkhfw==
`pragma protect end_protected
