`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
i54satHlwmTmHC2dVMr+0x/SizPH8hU2MEZan/usx6TS2QaiY97oesYU5VZhqiNq
N2zAWmn6HTe2STAUF71AoKQ538sKCGzAHot0m9uD0iyM3XxH+UON28tLQMcQ6EfO
D1Tnj370l0d+n9nueOEM3LyVhFlbLBOfjTJCAuZyxOU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12176)
aybmekTV9QlZmdBEdscAGcElEV1zItw2b+3FVooZ8Et0t4MIBcHa9AasLYWdA9tk
y3Wa15mIB4vNBol2vlVLjzvmmIGCZ2gdKkFx84Lbpa9c99vu1kimi2pexYSHQkNs
PprSkaCtYruo4C/C17YuHhHZV22SODA/v1JKjTrYRvKJhRfCKCFGL1FKjoJKRKvC
9WBQMdvmGAzRq011zFphoJYJk5ysWb+Li4ko9xhkh7h4OTyDSvD2hj1GngvKZSIx
Zg3l8ljPv1ze/GQM2fxuIjfJyzsoDUW6LeOu9APck994yBJ9Hrqq4gkE1cADCL8j
QhubzwQxfs32JKQUUQL2DjLa5B3AULqOxG6j/67rXvNOlMEKvhd1s51e69Ui7nM2
HSO2D602w+79aKKBCrlcExjjgZwJdnFiPPra4cP9A4n7qj+k4vWruA1llGZ+c/fp
G6q0AL+4/hgtaZ+2TafkeOlI2zHPMTzhGF4VYdjfZJpytfqhOgZbXeVgkQ04z+6k
Ueb4na495g9gGWXW5rZO/fT9e5i0I2ZBXaK1E7/7Ti9eEqRkDVTBoitzZqsY/YfM
Xy3fb8qYC0QQL4yRPF57g2+S8oIAgrEVJavripCiGLQKS/QtlrdHGeMXqG7URTT+
ecV/9Mse6Zxel7QwYLycZ1jy0zJY5iC4NZQkR6x6WCl/MJ+VeNnjpEEAnBlKV7/p
2N+63ilq/RvZhrn2AO3qEc2jxedbP+0p/E+iHLtEDnEL8Ho+oF71SKyRRg7sGKJt
9N3LC5W1XKQ3WoyKmN0EgSvAG9XjWGDNLjOqxzqpA+w8LOc/PHaD7dmRashi5t7t
s6Zbm7nvguL78wG/6FTgMxiAuXa3GymLo6zublAUamNSlVYPTksZP5jvA2HEIyH7
zrGb4w1GQWCuBrpXO7Iinxn/AnuKRkaCpF1MOc5hD8rco+fYjZX0Fpod91lsfVJ/
iVJ8txdmkjcMgXWXQ3hNl75ZJTU8O9L/v1bkKJcRipY3xEOxBZh2qJSD5w1/Hzkv
nUyF8qknKSbNmZxTwexKBHCkx2TEN1GUdjipvOS1fD5ITVjq8ThISEEJ90StM9SY
B87tR9MKiMDHyT6L6m3QkawO9nDaXkdohD+grhIluoSVxwNMOtyzJ2UZuVPpSHgn
njssgQ65DNHMKuQ2Xq6BPFl4pUUynN/aPdbnAxklWoLBScR5wbo7F7Tlo5G/n3dO
nQBoVGFD5p7IjBeFuk2MOPxDmB6gu8AZOQJeNwxaK1vRb5e1uBoLRoomuraYUW4s
8n/QqKHXKTE1jOYVi56KtUV/2f592w9+uSMHGBcPnYgPhg9t+BVCYpGB0Cwz5oXu
bt07Pyg9BVTMru9cvwnztLY8RB6qYGxK+GlqsjHMldoYNR4i7hKUpYuK6JjQ1ZBE
LOO5cmKFFJLxegKtOo8RRE+8RuHxPdH9yM1SgHakysxwJcwkNAwg8EqqV8lSnzG7
f3zrijLoJmIis98YgTX+xOo3YJwp9NlhbdxzxmwoVVn7BZHGJIaiS6piya4Xa+hv
D6hw75D6Gkx29Ph1q7IeEr4kj2sr7gkN85UHGdKpBI3YzhDulrwauGPzOmxIT/ad
EbUId3GReMM4fkV5LsrAHIqGAW1Ckv/wsXO71GpJy7vbAgBphv2GdOP0dbdhcmhV
S4oFo/9h/+grwYadnkxLnZ4ic1vnhAD9gYTMk6RnUt6xRssxktocfuDR8K0ZvWnX
R+hBogEvk1xMOBB0fopSKsIkqvE2fJWBubjEwx6Mvupt5C7P+hI+hRigEPbLSkub
7NL+tBU02ZjexD4f7WEwCHPqMou6+q6nt6iWgeP85nfMht0kyLiIcclOrVsUN1fb
h7V/oArsHhn5oT+W8eQ3gmfOMPqSSSJNbKZpFNcY8tie2xsQUS5PuTqzGCp73AUl
lxgt7DW9mwSpvDjN3iACffpExNSiQe1y259MnbX/OE4GlDuJdDvR+bwL33CdCryJ
VpJ8YB0wWN33EpOZOAfR9p/CvYhuC/utdLqc+b93MhbYZ/iGXz9I4DwVgpW5Aa57
esgabbmxSU6codHMr3+mGnl9ByliRB7DBUHXsLIFJ6zA09TPXe63jSmw+HQKdR24
Jtphuonkc2QqQ540+q2LoAYWKrSuEf8gRst6uChcR6znboh2DX3+1TBhT1bdNngM
sEPJb3Tpv+4v/3Dno0Qi/DV6E4tgrBOfhC+XOYff5xEL36/GzjfdpM/Bxaw6MN7l
MB3ST6yP9ynew026sSJi4Mpg1C94Q8/y21fWLqWcnrOx9Strhaj5hAffLXpf3hYt
SItfFWIWXnUA9p2i15oGhyKNUwvebQCTL9EX7ZhxwfYaygZB2d/JpN8TQo1M8xet
NoHslnMYUczinYSQ6kiRw2EWOIhYzeZHfOP4sC5LjI+IKqk8fIMudT8x+6bbvepE
eyP1+5umPg17W0mnuVtCFnWu1jIPUeIp6YakIOV9SiAJj5GKMBjcJWDXMgyeqpyo
VfZWn4aoCO2yvrtnM04GXmOj+unK7DGW/ff9UbcNX8ylyCqzr/jvEkjSqSql44wN
oxW4Ok8s3Mc5ZsAHn12B4jrpAtsy5KIsySvd0hjLQf/d4O4FdBnfI8oEgvzWL6wU
4cEhpsgRawDcY4OJXuO2LuXoGiTK3657oI9lePtgGkZTMZs1SeraDp6cAfww3qBE
osOvhqeseUkl6RHgi3PAMXvwRy4QemSkQS/OIdEP4YsGqIifLzT7p53iCasJFt1/
8oggQQOVXD3+nc1tbaPVpev1tyjlRNOyi5W26wAjF8IaZdUj3FzbLiyAZUcrByp3
dJeHaUY94Y8grJ61rRHzv+P0jKLR1LBnCT+yKmy65CY+laGvXokkUJU0T0akKjww
+uXDvr2fY6b0faBoPJUMidf1mWvFxpRnoVzSAb0ncR8frWNG13ptcWgzZGYyo7x4
LPMmZmGgMeyOjLw61mTSjNbUHFdcTJ+LXzAhuzqJ4j/oejQ/CkJNe3FgQNs1fTFI
vmDpQBXz7ViLWl2pABAzIbEdEq1f/xoz/aQr6gIPSkCDyoJWs0yJyJG0kvt516oO
o8HIGw6wMw6kyWCdXFWcZbsik2ZEdzaxBmUq7Qcg1awa+0e/Z0g/XIkelgtFjTZJ
cRgybrWH8Zi4fmmb7feo8n/w7qihICa6z8bT4MREs7pwgw7Im12LI7/PCuWW9PeV
iPUXzO6sUVEPT2jixkzWowwRrtpbwmCFPnKJTxv9OtmHupEV7MHsu2BQq9ZA+GqS
5+W84TAXWRwfdNeXB+nlF1IOjjdwypBJKlH+GvZ9wJEuYWoDzEZdePFZ2Jkr2it6
1OLmrwS4+eCmfh1mW9IQMBLUqCCfZABWbZhqy2U9bmsZXQ1xmWEneuobGU3gCzVw
9qKxjyEKPOEiqnhNumx9uH60warJpaEofjyEil3h1X051BumhMcODp3VEOmfnB3T
10OIVqZWaZSWJvyAqndHjq8qsB5tiXV74oBfKpbW7dDee8y3DHAQcRCmGXkZS7gr
kvz/Vmt2l1KFsTVGUvHWZtkVdYAwLLxjz8/oluLXnvli2iSVIjtuJuFn2UFBajuz
H6QUny9cgFVEH4WGYHcE46Tj+YJidXKnMDuPcTUUjuOAWYd6isN3Vmod2uz2YoTZ
sFFvTYibk5TJYvaWWKXuTPedz3P8UylTHMoGjzkEp8a2Jm1w9yFeqSOfvrjBRY4M
x/oJG13BcBi6+2Qst8SAQMULg+zd+KYytmX7uv+JOQgSL4+A7kHNFElxTo5AlDm1
rK5ym2/zlNa8HDrjsfdnJk9dH6wrHmLNWgSveyQsdIkFtgmZV5+0JEvnLaP7xMaO
3xAAXpK6PA6/PdUMX3Doyg7ZIDCzGJRh8HFUaK1EJdCVuMCDnCyVRAuY1xQplj/e
gMKiw+bqQn30kgKYmz8UEV6tYtVwel2P/ilyelOHP9Lh0tUtNHC1wTpmQY8taHNy
1WNSG5IiBZ3KqfZIQwCnzEKXFD7s1cu9jeZcDsx7tBqwxo2PLMScMksZ4v5g1NpG
nCUNeP91Dmu/AV6K+jWhFZL/YGZjL1IcaDj5TTyInglKWvSvBNCrVZ0H7hcznK1M
k8CkDG2J5i1hR6x5XE2D90ZHxdb91T/co8az1+ZclseYwOatPT/uCwuYT2q2yg2v
45IwAb0RXANjDH2yZ7JZKVwgRVIV6omsMhc8rlYYuSK9/dUErXPqZCQiFk7ejJG2
UtTa7yauPyD/aBJP1I3br7dsaZLYc43wyWlIlwrik2Mk3OeZH57WnsIvHvdNsdxO
NEuwCTuZtilpLwEX0+pWczTqM8AopkoPzZufokfPmhS7M30i4kMKr7V4RGi5fg2E
YFIX3jZctGvkDoU7363Ek4tjKFVi8oDv+6N+K9k9Xp7mJuApFEYUlZ/aENFrx1Fz
Qpc7ilw3b93RERINiJBE5X6BUTX6NuKoey4nexRgAA2HjLVqo/7JI+f2bcSLNbOz
6w+hTu2w05BaqW7f038uVInXE6F0TEpKk1OxiRIe/4PMaJSbk2uRJ1OsylH8eyMI
2KC84dAa8kNWm5Q8jLSI99qTF0I1u9hcdUMGdGrU4Af02s/sSkuPUENW3TRWZE1/
ApuNBnhUoaroHHUuDi55n2LYMYyPCIV6KacXfltrwapLIwpbaqfH1u+wcYzglQbt
d91G/CvNzruYCxK0WvsTREnNSbVUWBozkrLGXaY4nvTCaC20oFEKF4qHNOCd/6Oc
Cdim65OxQ1So6z0pa1ilK1iNaqYDv6Ggpo7rRzOegqZv07nMeAB7CTE+aIp7xhKP
Uvp02eByp4wzQITyQ3PqSvFR3L9rQOlkgOT99r4gWSiBz8YQNhfArSoPlHeJFxVg
qNtyzyuWs53Jyay6l4xAHjZanp2TW56x9CjNA25ImmJVto9aDr5Q6zCpm+aUu7Q6
wNX86Hkt1giqw5brmYnxMhZPqul6uqj1dT8rSDlmYNtJoi4J5B+obmqEQ5B/UHkX
E0Ml2g6XlbXbs+Uq4Pe7VCQyCFBSBqnfilpgCxIB4vHQpv6Da/tCDaE0ScHuXMNR
xgPKKg2+BiyrXe/UqH+3CXhOSHIb8HaRc0gIiFPBlrPfs7wSYWoD76ekmYhD/Qjk
DxJMjAmsSdMLjLDBOQgBnLcKB1Zim079AL4MH0KeIu7OV/VH4vgIQnf0XfRX9W5l
OFd/ZsUahmTvuGGtVcMxdSYiIGcWKfjDTBSWqPgMouDGti1s1ty4ccCBIurYJ5DV
ZTeRaxvP/ddfFPtsY8K0bLIhbhpuTRthEg3Z8sbK2gi9jgIjZsbafH8I1THabUZ4
zfQTdd7LpHJ0E5zV6Qhie8eRohkhB00fB959f4mZs45NhAjBsGwqNa10wHlCtkxg
7BxjrSsfOoDCALXX+ZuxlSe7cbZa2d96ehxvrhrPHPMwKiCDnKg3/T/dpDvpeLmg
qgxZZ9kMv56QsPwC9+qX/paig52hypShKO/FQAccyCx0ZbJkNuwbIVTIH3i1xvrM
lj3qAO8eCot6x4OFjOmNmH39SB15jjh48y8HJY5l5b9x+xm8SrMynzgwzo6haMzQ
wkAiTHQorqz4AhLEYgJRQqPZLDRwHbBPy7QzaK0bv49BwSTraOqlEyIiSPb44fcq
paaZTJ41paGNL98nlhLwtcmOKNJY9/Omcw/9F0prEuytTe7lB/7mplSSIU8i+4WO
4ou0/cU5kM66HLuk9TM/qQrTm+F7sZqg7tYlosXXG0/ywqTcql7/2aSKtNVzPuRb
kiKiw/wD5VYsrKtRMV3VVDaI70l+S0p1dvkyO2v8JC5Zbzc/2o/1v5YsOSTGfKTH
Fvi1zLvoe5x9SanP8nOBmrlzUdB2sP5h0sVB2d/fb2o4qAlZfzDYsn2CHdisHHCq
VEEAEymv0wj2b6i7c3ZSNXh6u9HbvXYq9EGk7mavEtZR8/RO4+nBlpCchESRjmL1
udtUqSksnnZ6EhDmP5e4Y722tKq4xjxUO4vPx6cjjnBQsqsfmYfP35vTSm/spbMK
Z6CkB1BqaEE/82JqLiU6NkU4+D2syQs/EbGh+rYNx4ccWui/Qau4jOUkEKrWIk6o
k56GbDApYKNg4uZFW/JJ3IyWVrGyTTsfliwYr6djKkRze7LJ/l4FlvGWYkYX/5Oy
q9aY0XvooU78wEuNnxOg8cFF8/SdEBD0rdp5jSQ2ppgIE4GGHAKI5BfxNeALwBwd
RuVAEFbORq20DeonGMbq2SiDm1DiJlizE7lTLzWdUw271abBCLLm2TeyEPfVqWPI
PgRtP3Q1OF5FoiedfT+4WVel9QJYLS3IEIURTYyhd4ImhR1ybi4G5rhxXn4xtd10
XfqTvYZyusR8i3dW4nH06gaEy3DJ6AZuIs1Yeqbqzm90NICFxRfnGNEg3DBCcILC
xgsrulylTMff09FSNMDkBeKFsUW3je4Cb4LkipNE1xOX+/W9tr2RXZhZoraMrkI2
aoUcfhQ7HzTp82qUQ8XoeCaiHDU+Gp4CZQt7kRsTdcLMrPZ/L/HP5vODmY6WdamP
duNVYn32Tn500QvSKpxP/PQL03qhtbR9vFiYr2M1UeqQxo4mn3PuAhHuiV4i9fxQ
ZryX6hjoIrLdrEffVHtZp75DvwHsHOX0Je+T0U3J+Ia6NWi1YcGFah5B5bimQIh9
iiUAbJJj9IGVKeFD9ewgKtzkDz6MjqfI6w9H2NMcLodTZq5zJG6dRfOy52dFjBGN
okDDlIh0XA7wvLYv6UvDVy1EHS/oziy8pwh4g8qSVugcZGrg06PtxjpxicmxGabn
SjX5tMlYNcLUvGSSwRY/XQ9n6W2kKoKWvZOrk/VK44x8ov5vvmQin0lV8gNc/gLU
AHVvUIuwRV9Lv6UHgOhN4gdib5rk/LHrk4H0KsuDACxGibd8VAIpSRd/jORB/bCC
iYm1zDffph0nhMw0jSsoaPfFPm6SaWlfBFBooYmXgHDva4n9YjvHyve6DkN1S/6T
Zq8Ef8KHc37SSvO7iYllnsWUvCFlNkksRShfW9Mg4aEnT+vp8ViY023yCGVgt4Ci
5UK6SU+Mz3yM5mUqOmoFf2B+6jBAgIACBnE2VD65mZBzvMrK28gKQfG3rGqPpCHU
i3wpjeLv7IU8bRXQefrX6/mlT00WJ/o/yHkHHl3gAQS9GCEQIgfPDbJxGoeleooU
0RRquZSrrwmMWsoVrg9ogFbFq7BZ7p5++/dxGGn/9dNV+1Y7y96bNVMHGWwtK2Py
wPjxgIUTxvpSb9J5fPuwqy8TkYkQLM/+wYj0YNu4mNkBtoaOvH2UEAeRidzzvYeo
Tj9OMFSzJmEz6muxgexSNrZTkAKzkQsrjsYaPbH8ww1p0HGMLU9SnPFKsDWxnnDp
i7nPv06VK3kPk+bzdm2DHheZPyqTuQmDRO462Ii2E4JEjWlTn4Bdw1l706wmU4GQ
sAP+P1MOZdL4gK3SAn76g8lEXGf/jYfN+q2yTl0j+doROVQ3NHKEHLzmlz6R7hUG
DijQMMa0gqlOL3nhtoTD+3LfjRqGOFHymME9dnbUvuL8/IlCLxpb89qq0EjzeqT5
AUUN/Jn/M9buKQJ44A4RGmm1MRlctdNvln1oGrWbZA2Jsi9ME/dEP75uv3oNlWPF
XTSoUR42lfW6yPTHQDY+fglQ9ny6PZdRBXt+00J93cpIsz+IcOt3ok2wrBKodRSn
qsjL2Cb19+CXUMz+mjMr6b+SPu0hKfSOrTuUERqyzUWB9Ol6/OQqO+41jzWZiptx
dFzpYXexuvzSMxtGoAhUzd2JkDpYwxibja3m1CjzNVPe5JL4piqGXO6lLYX8LezK
pibvcgIJStjaPX0thjN1W0tl+1jnRW8D2VyCB8Im+5Qfl0niAYQ3TuS1YA9sWVQ6
shhVP990a2K7eZp3v25P451SOhE/hFQ9jEPbKvrsKFTRQyrdYqI7PEMm2C4raDTp
PVbbfb7ozVmle4F4eUOMVnQQ18n+rAaXImdRt44/SAcn7liTLDOP6Y6xcczZ4khq
5T8YU1j7fPA8gDM4qPF6CCOj0BGXpWTxWmH0xuTLLxH6B8AcWEIduzi3rYhnz3Wn
LTkH61LsRygB/d787wBMkGWpiodyv6C/QX1YDRDbqFUDOOsDAG35MOY2Av4TW8+5
oXHzt3HA9IAnkyvEnRd/XfXAFwcRWk3mWC9N6NlmMIF7wM95IiAQfRlNXTz/y7CO
/5BEmwA6EYYgFmdLeqlzCdaxrp07O+tZiGu0s7EY4wJtnNabONGUrFNmAiw0ABJW
FeridRARQM3pf2GWqupyeTF6fFsN6hlmO8Oz9HzGBU94kd9RayeMVInKusk9Jbb9
3IEbirsycjqTfI66uYCsTL2PU9QDlPhXZup86fEvxVAsc0+5Sdj34rop/TxLki2E
9FUDaNJGjv79FAASc+JPmLgrRFNjV/JEeAJmdQrdmecrYq3A/M5cfYf23gb7f6nK
ORlwt1xtA4gQpn3o7+3RLKpa57UmARYPiF6dU/ujSCZ4KykFWgCUmhIDiov9rcDT
j/Rlg6vqqYNayVHZlj90T5gixFf5wwSWbABza9YwPeyxhZhGQPPu8MpPuoAhP4uj
OVKOctdZHIJjlqfnec1bUD0o0anAs/I7lqPJerRsmt3blzwqFzGrIXA4jLrns3JH
mWMBEuDPrxVsZC34Aitz1bZVBl44DACYnwsaxBdVgBbRzKYydCy0fj8i/yjPiVst
pJ34ZHDf2JoNubNfV7uGIRH5A9r4Y+ofd9D5pqaXPtsh1AmRAo3hd6zmFVVCInJu
Ho/bC+qcBVtSxJtSQ5Zfoq9hlqPtINO2Qn5EYn3M4pS9z7KBFNV8xFqH6HkjVHVM
se+hJorSgGphQ6eW7qpntMCJ/eMjf952mjIW0VF1s6PoYh7yLkZ93IidR82Jo84E
DsS7sxo35dyuHZRObqbs7FD1Vbsngoy8WGg1tEuWNh4iEOVSF4/3sXCgBYOReIu/
h88cWQqRAp00zDT6vhMzh4Dx55qcJPa3Ldvy/Mj+wuW1/utmhPVqAvmk1c4zBjiw
jqKqQejuXd9MSyxEore9jGFVpqTI/6jcqNY2ML8bOL2QiFSnOFsiwCOpg3EIP9qa
0Zga3Br4hiz1Ug26sOkfTBYuMupHbU7lzqCegry3gIVs8uruPyEVTvvyrWieWGSQ
sVHSXcPKlz8BNtossrxxKJm+agCzJ3jvirHYxvUwSWB/haXX7cLBDwFk4O3H70lG
7Cj9+ha5RPxKzYZ3qOJFqxBAoPM3MXPIEW8EJn7TOYDqwTpT+zheeVhCXvOQwmVe
O9UMt0Tb3INBKWO9s5AnM5enKIH5Ph0V+hKQNZ9tbrXSBZUudEp6HmsujAEQIL98
PC/eBH7F1Ez+Ti/t2xCeMyEgokdoY827riT50e1AtaTxBLQmEmnQqIYA40BkI0L+
7ARwkW+bq/mjt6KbJJQtFnvGhJdohxyhXxaIPOoZ4cyxsNhHyHnC8a1soozxnAzw
N2lh5vMQ9Q8Kn4cQ2ou1OXo0mL4bX6AkZ6ODbmt0Z8V2Dlm5CO7K7pRTVLu1I8/4
4Avg2vMtKn304JID0mZ8uGRUwK97HCDh1o5BLuODGYn5k+fv/kXkyRhFRip9yMZP
n3P0jSefyjAm7lBOx6xsWAxHUDlW3tXfavnOzy0CB8NggpS0Z4tbolf30LqJApZL
00MlZepUC0l7N0B3NxaWyTdntRzH0Ft/qdAfSSqcvK+SGgLwDfKPwet/7uglvCfa
CEkYzDhHhWT0X8VsQ1/4nrNik1OF0SNvtFpWGjQoOcdor2gZnXX5Y0IehrwnxSPU
/o9EjH0D/SnOJ2T5bTa9juMZU8RwkpVEezJvemBo3rQn/tXD5yPKpQ91X++xd0Tu
xbYpz8STp6wN0zhT1/YVSftkuVXNsY7sRVqXLeLTTUe8Mz8c10PE4R+Xalbs8X36
0BFBSvYyNr8/7rVTCHr3ZPKXFNRqojztnzPXpbHqXTYx2bvbwbM6WX+oRsYOEeS/
AHEgAyRLBrd4zI6aavOcYdl3n7egWxzAEfH3d3IuSo7XhUXkCor6beENfW9Px5bh
sKCjV9GZ3Dv5hjfAxoWSx6tC7WIyplf1xbhPd01uP1NGIAcehai1/oikePljBM9b
C+6AMXEEAXaZ6d+hCz3gj8NCnoTb9pC+m9BhRR5zT3kXLX7eAxRGW4r3RjiKCdCL
F2HiUMqeis8AnNPz+fUrQF3j1bdxQxSdNFVbgrwstnRAISExiyMKv3Jo1wf+sAog
lEDe3JYOvK54YhUixhiibrLn60tTp2K4y/9NGs7W4x9Y1O7AKVSoPU1oXBHbcZmG
YQ3+a/kr0PoiNdfZpGatpl/73tMdVBYXq2Xsaewg9+C40lbPIWvTPZjdXxla/GN3
cie1g9UDMPKcVZXtLYYJxpDs4Og/+T0t/1lQvaY3MM4BWJslCqZhTlQ+6KtnHBHB
UYy6JdINKQErlgS3KvxTLbwRnKHi342Djx5aQKaze9yMgeIttl+qjfMDgSFqz+4C
7PTa4ZwLCBQSe/kJHhiME1GcvyQLAqRIBl4zS/C8ScOPe67JwEKuwtPh/4VV1pDu
rYPQcRe50XyNrOK8UOXqyU0VTr5IZPO5lc2bRvc0fuzwYyQmpTP0fJorUfV/vyNM
9gk9d5FjtI3kAgpDdqbOSv6PClKh2YNvndFd2FPDVMH57CxKCaH8HkDjJ94os3+0
V1Zja2JJjMI4gQT999YCF8FA2hy9RsCoOfloZSq7fFVKYBGzNGGS3kUjWzp3tGSt
Ksc89ctw+Q+jKouIwDfMJUR5xeB0zVvHeImGaGlUl7GYeN0RNGjuARW545hO1oOr
owtJCLyv72hHWIAHPBv2icJqRoRv3peSmW03/WyA07iZJayFTjKCmpwAaBejGPKf
kXCGwBj6Skem23frqO+Kh8UG6EHWE5vIgqWFfJHRCPbD+kt0HaQRtaK44JjgHB9F
ptgbqexFgtPTX1HRtYHz9PxsbMPSv6hZcHLy0cGTSESKyE4Tz5R9VgU6s/uRwKHw
+tOA43RO5fNLy1NXlBTFmskX8GzlfKu/cJvweCXiMz0BLOJSzrmWlcLP9zWPzjWG
xxQEbYGGHgJNYT6loB7eU8KP8Qf4SFk2f0HdgFueFWZSGoCeoveMxEhsGETp/ZV9
rIat4KrNtOW0QDhVEOGtglL3A/ky2+47yFte5Z2b39AiRss43Q0xCMSvp1/ep3ap
u/N/xvapobsC3sh6qnqvEf8bfX8lWHlySt5b/Yi2BojEPYv9V4j6xTZGQdePVXnn
QX3/oxzyNv2WhPqyhMO93GGpvwn077xOevVNwl8/+Mux037ghtmr0OSP9NMcfhZe
kb7TGdXmlFJypN+xEh/DNewIVviGbYnG8VCkjXCvfF0eRYRhEj+CHNinsMKMoL5H
P7VessUGefSTq2kRrKZKzGvZ61nht9o3mPF/ipGquesrOvZwi2EjE7GIsqEKPUcT
qfbfj4InelImI3kStOXdHoSEP2ROIFmfvDhXbcHrz+sUAvrw5xmog7UWET+AL6/C
xw4gv/qnlaU9rZy8ytLqTsDw6Jbu2zl8vvZijgq2lVkGCFq0ShGJDlM83MJC2O/Z
mGXoP4xgwtg2yCjsbZwCbqGxvOD16m82oNIdSuiNj1MEN6s//VktDvPLM74iUOjg
tj2+cob9KGzVWnOFV+B1r/zb1V3qz9U3qsVAjF1nhv6zRPM66VCuNEtzCieU871l
zWNwvlWIuwtH0uCJQ0YlD1uIEySORHkW1ffx7/JMYKrS6YlJ0vIjbpm07xFXkzUg
AgBchK0K3Mn6zBTEOl9pzN9NBHv+J30xqYkZWpnBPiuuhImtwrn0tILM6tGqkp2r
DrzY4JBJaflvUzpauBUjizvscp+R4ZyDjSq6qJpAxvMIpQs0A04vzvfrmLxebSE9
5nJBc3EIFoQLeDxwm3RLsIJJ3M9Fy5q4uc8Acc2TcU5h8/PkmQyTPIrzuzOEvsOP
UJoWmVGt6ss7ij2JvCYBEF8qiZY697emk5xKYxlSGIgeDZZVtzZcvY5YA+C60oGw
WKEEO7v3L1VyyIIYtQJNL7QYmyyUVDrEiHBebYSyCN6sVDQz3/ojFVpJq2YANIq5
cLqmRBoBbRrE0sQJK+gfu02rn2QvGkok0C4Jvx/udICiuoZa+qJvudQJ3yXTrhcS
Ldk48ZWcIN6mlF4DXvsy3cHLrtCjqEyyW3rxc4539rJ1QXqTLQyyxtzLXMpEHyKX
1kGfxJYlEvAs61q3g1pijN1mYy9nrWOntQHlmJON1tadNFOanQgM7a8aNV+dtIa2
r6v6706/mCEzZs5kQLTPGJsJU78z81JBoH2whIxuhxpsRDxayWZT8Ia1naswQBDo
I7bGBN3/u+L1zlg3OkS1NiI9INBfwqunkVEkPvL/eg2ZPL1Xg/AJ5EKbT22w+9WJ
dzKRfK/XMzoNtCZBqAKlrDFlu72CZbUmNiH23fiLfyz0sIed+n/FvavwMnukCGHw
S/U9oLA69srDe1kTZa1VFOwBb2yqo0ikPAlu53D4Tp7hK3LGSRW13LxNvrcDlIoh
FLLwjlRdLLZNy6Bd+vUoGw+IomPk/DFs/nfuvCQyYbLpgBUve41PpemgRktgJlKu
uAb/KH1Nsgjodw+DFM3DjrWyr0A8fWBtaU1zwUlQ/+xvkJ+ne14+tWkiZOokwt8m
1PUohmXwF5I8JTMLPUwWJCuIf0xpgLC6NpUpAti6hOB5V/fn8kWIh5RiiiFrrtZ6
yPiIpimuodEsMMSW/GT8TFqD9lqPGEGO4yuqfNgxVu8RB9cBI1D0KlytsDe0AdN9
6lWm+aNLZZnLkwSWGY6R1hHFpeFHjFU0VsTZhzDGXFpBRbf78Lw6QXLqhzWZrx4E
LXBi6lRHn9Q2uBuGXOEumzVBCOWgMNSzpbAlv97lvZusv9HqtsWG8sIVuDRjj2aN
K0Q8ox9natexXA8H0JFRU6G5BnQZDYJOhpYQsbfAIJQeguJz6APeQMduvImrX3MS
N4bwjds3c5lXL2Xqnqpz1K+jgwjpkpHfsgmz/6bNw/GG+91RaYE749h4VkomIM9n
h0HagpC9omswWUeDpEWxuTFHRuGfK30WlsxcCGOxrSFHYP+Po3STpfYywvRl3lHi
rpunOISpmZ+9JQj1hL7JxcCRbVWkE1AbqlaLqI9CoIK59XiDxMjdfk4ymLAOqbyw
EOAXR4sQsakIf9sjh88PL3QgLLGtdPYGjLiQ7QfEueL1boGFngq58QnHIFC0P/dT
ILkLAV+ztosZI4OL4gcBYjApaQoOS7Uj05QtHU8pajK4iZRadga8ZdV9pFUan2wF
yequmfiifsOu+1Cbh8Ihoohnz/JE0wSKSkD45bNpVDFZzegEobmAZgtFnfjffOYq
Xhib7da0ouE4hHstRz8wE6Y0ZD2YS2IvoX+NK8R7xrN5NaMtMJRMkHYFHPmI261A
GR35knGjqrseNdPym8TI1d8/5iH5jKRpf4h6icmjQCIH5akORW9yIc1t97SXFTPn
vRXt/dVkfm36LoaQjAi6lsP2ZuJyt9sNPlMFqbfPqf/hIjtz/xUNg4N1nMzv4mc1
ggwK6BbdaPqQcZSwgoBIa8AzcfPCD4d0MRUacsiK1ofBX3D6uO3BLlBfZx6+byTk
eumiOh5Q1txQPN7p/hj7xgptj3qxPv3buW/iU+Wa41SJEjZ7MMuRyP085qdf43PU
rMfNLYDEmqbmg30nYM4RTSrg1wzhCCTdo99zorxfo0NkBB5p9nQn46pCk+ydmqHt
pIS+sTDga5HWkIkrghAv/5XF9xan0PhqKeABWT2t9borNKTt5/coIHVyhR5RPnF9
LH/rt6DNgxWAOxXrZrZ7dYd74EbGF8CkYjoI8UUbxcaT9kLRJkwd68B0Hi1hgRZC
BPk/lo/lTT1hVVEdEsMtdWfYmw0+vU8Mtm4JrEZ7S/S+typXfd61rQeF6qIJPzBU
af/N2NRrvB/jRW7uBsRbksgh3t4925hJ0DGehkVmld+JO4zGtFeF+YPaCsf+stl8
Kv4L79PvINewz4TJecyInEyETjeTu2bM5bF7dSmSMHWcSZgsQLLxBwkmYq9vopfp
+tBoRT4D3ozUsIGJDLZmDYonwLtFQHt+wK+Xkedh99U8OwVVAgoBsZs9+wF7zs3w
ncbi3SvTzU5Qf1xaAsmJaUmOEL5fcAUE9o//BrK+gVKJJ9ZN6p2wgEHJ1oiriArl
AgoChWPMrFT0wZ1274diT9KfxRcKbDbvM9VKt4nEMmpUexoyymh6aHCrQFH6trHj
r11f9aHj6dr9r5Ky3NR+dqZeFoto0EppE/1Zk6L+Y0lBKQqd071GgB8HKQ3WGscn
cvL/BDseN1vQbhsDuEW78SCrT96kCO/rT81+VG39ydBuG3N2Qr2exAqPE+KpwYOy
1nXdONyAeeUt4otI66IU86sJbxddfk2kmMl8lRE41oaar8Sd94Ridd0GkIjj4Gnn
IVtqqawgHbb/9xUjO8RUu8nHP0I0vUNUxFWZ6Rqr+wbe7khqXFpy7TdiPp02aw61
nWHn+ZlouVtG4nQjCKa+UEsrhTQoZJelmezBRTo2JzgZF+kFKgB6j5iOdloKz2gH
0iFs9izGZPhvhPeq0T23QWTYLTFfxyO+44N0JlTuNAOCJ59yXpqNKAhVVhQnxFSC
GoRjUOQ6xIput4QAd1+/X1EM9GBpBZMAIl8eq5b7kcXFGrncWT0DbkhlpfNEg9FY
nuCFG+VE+iEkjoIfOB4qsZYbukIqrVs4TF6Jn8Ww7dy3HoyX+1DFdoulPA3KEg3u
x/ves592WyFjKVik/VwvRDTo8BeiBcpgJljBfrHF5GBrONA+nXJY068ERd9Cv6US
vKt1xkbX0GmCBb+Cp4FnNCi/qQ2QWNfAY5K3G6G0kKBceOyGSzzmPB9o3VQfkTQL
yWwgbBIsjlc0uwg4D97AU4JJ4KitcNbkIGbQsepshMMmrcGSxJDlE6ZZDw2jH6Vv
xS56l++IUBdtmE/TRkGfic/O/fgOV/PbmY5/pXqNqeco81GBxdD/sb1mxRV7HG+0
T5GaRBY6eMH+xReANZK93FgIj5ClLYUUIwJUOvELPT/337O/yuZ25jdJ1l/I7zS2
Xd6dltdN7IAPjbAmgf1Gcl9VaYQYcgLDmjbgYkZdxiKjlHqkD9zQJKNd8u/N2IQU
qMiRL58w1LfMqUSTWEKDf9OB3lqj7ldz/uxkc0Gx0v3Dhdqph+1B9Q08DVh8QM0N
RtmwdX92DugH+4MLMeXayKBzcd0TOVgh0swIok8YnPqUQXtaL2hFxqucZF2blJ3n
01mxhQfhP4IQodqD2BLWLSnzMywiPt+UldlM9tOm6EeNF3r4P6vBQhl1vlbwvHdi
QQE+G9c45HptQNV2w13wnemkYc95DOWS+hJHidFqIP1HZdjnnK2ZfXdm/mwcaQN0
QCUsqljYmnR0AidaBaYNMTU4+nmdMXHYoPFI+0gzJXqPLxAXKqny0/8wdsyhfpte
VbaZJgkl/6/f+fu3ydEKfcAF2x7LFIh+qZNeCuq5kFoPfUjpfes8OqMg+FR9GdzR
3QcFGySwuNrb5sclo3g7F64YBw+uL7sGxPyittFSVblYZ10LSGT84fljJ9/Zmrpb
rgzhb9UXw2IgVHIr11nxO/sYvHlOrFc792Xj2tz8QsdXvGZe2vyVMTFlolBnhnKP
yMV9nZOzdDAFcgGe7hdp2F47kblSgvFin7eEAHTRBWEHIIlirRaQZKUEqTBqHJbw
li7BOzHapUt+L8i4FLSFB+YFYT2QQYka95ke803/Etu+yE5FEFaUAhcc4YYZlm9S
xl69UGSPcHWEohkW4ugyDth3zRFDtFn2MgzuRPPclJIsgRf86eWzFmZFp4HFnM1p
H+6HrkZQriXZdI05Q++F3a3MuwtpZVAfo67AJGKFtV4Pcpsf/N1BDCgq/VVeBjiV
aDQSRqGsnD/Vuy/iFIGAtAivTBBSTjLSP3EqRhdS7iOSUAS9eQ7RL1d/YP2givdy
HVyVlR95u4sKSaYRsQqmeLgKr5TBrH4PwwFMw+doPcdxgvohyuT9gSHDwCqVYx5u
cva1xY2m7NjNtr+1mdVmpTWfjnvi3lHrdMYT/pq8oLDIIFlrek+xQTZiAwX9AP8J
OYtCaKyXSbMAJaQlXP8w2ZVHw8lTCJC3uGM3PxjfswY2Cw2J+0PMkHgwuEzu08ZL
3IwxM76XNKZJlcIdkyDeU1U0aF8cSuSiKYSaELfHOmY=
`pragma protect end_protected
