`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UAURpCzVcUyE+AhSd0yGTfM7X73+6GFtYCBdASRFUYsln44T6svsJEx+H+eQ2waV
NTwAikWO5TPjZaJQ1Q8x2YjwR/CBYrSP9N9JiHpVmjdFYxnaA2ddnuA12isrQmqi
wouYTnjimrTkShtxv9O+0T48gEZ/ieLx28hMjlZsTsA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4720)
O0cy0CQHq/w2ejF/KOOImO3tKDUlLLAsasyXdwECn4RQr6SWMYu7HGb/TvPsI3s+
ubEG5zmafFdQxCFlACfSZMzT5Xc30vVwjAjVM55hH1BVcCWbLd60xNZ+kxwhdmq5
M1p5VqJYteAfF1zd2FEoRPn/9TO3ygtxApKFx9lXA05uWaBkFqQW4+RYSS9mGQ3W
QTzsoDjARjthGixqZRWf4zDy9OX02upWOClpG8YEavHBUIlmFjBFvqGx0W7N/HL0
IEPY0m4LIE1xrzcQgJvE+HszMm0nthX8c2rGnBar5N2Y5yftt3N5fcebF8GLcRet
eV+uWXqW4SMyqk2ia3pLx79R9KOD4GcXfklWXE+wgUoMvpaDFaiUOf3vJtiN7EH+
IHD2UA8rvQaE3URlk8m5CgLAT3zHiZNm/SyuC7vBNC28zqz+93PFTZ9/CbV10jza
dbZfCLVrg31szXYq52HedC/3s17oKHWZgMAqX3OaW9zVmFfdackUciPpomm+lne/
uwk3uruoZZn8y15xqa1jArudODlzCvDfBfCs6YB/roHznpp3o7n7xF0K0OmlWpII
5QbcO+pXwMq6+odP2EAcpdeS/3A/zkHp5gMDM2TtVhHG0xAUXrMQTQSbhq35yXcU
buXQo8S/mSWMJc9/A9urax+oQOJFbH7JgN4LjorJtHznarwpTMWvytKBZ7OP05OT
crYU2lOhp7KCWmz0CzhtK+0Gqh7hZ0pAgkUnCMeZPf1DBFs+kMfHGP5Zx7il0uHM
adOEzeRBr84fxERwmArmVDJdQPI2g3Q1fiHxTUFKcmnlWLSMQfCvg6dFzFGfl98b
QPZldybNb9/OccQDz5ppoz8fAHz3J0vZ45FWzjJK2oeanUmNvdOL7MSXpS7bZvnl
Vbpa2HVP8jfyl1/Rj9HihVnTgruNUIdpxBW+OTTVKO1PxLd/G5HC4qdmdifaGTwF
/3HmZLQEYGuMbn3EGZhJkkGfsUwJlcufHktgu2eFXInbebww6jgx0vgqse4nAvj0
fa93RAONFSwmCNzpodMhG4Gz0Dn4Vl2EM4orwG+F3fH+wHsJfJ68oOtmMJAS+R1M
aM7GUImdEin3+CZU84ceRliM62pIztcD9lGjJMJBbICwLT6kMR7+wELO9wMgWcdk
EIVbGr54tKdIcJeYRj9T9TrKqF1ugr2BHLAWhLMqC8NokGnFG5WATlpPhTU2DHS/
RWwhfCRDpnuBP2Y/Brd+DBvRkTzOb801vx6YZYXvyAE3OL0UmyvC+3Vq5nfHdFzH
sQGeDBicGge37rlJSx9Tsf2infRlOKpUJu9WEhn9sMItl5/xVIH0xlJQgJ5qFzUQ
BuEZVRc2v9LPKsiSjSS5KLB4Kskwpo7k7+cZ9zunXUGOUgkBtp7Rm75IaqFMpIkB
Ng8migbuHa1q5uAk7dAI2jksZXO1XarKXqVrz2ZquzfRjU46K/ELxqiqdXtqsh+J
8A8vIKEpNpRK3HO6eu1GypzsBwwNUU5JZMAi0yd5wGRfkCJytQEmz7GxXpP/EJEQ
TlsHjhHTlfJwZ8tXPx8Ng6Y8e9q2ULUljdT2TxWJBkOZdCYshB+dsP+O3yFdAYDY
vhckn9YgN+wPbv/2Qoe8fJvC3GEkefTPDfmygxDF1bH4xPXNZ99K795OB5JLJU1D
jsM0y0r8go5WvVCPKjKrJffC9tzzAPshRFvXv0hGr2ZTx+baFPRy5uDpQQduPSRS
JTYC7U/e43kEsZxUtcOSx2PRVP0OzmJvmdBY5D4902b4gS4PtaRb9vhh5z8nw519
4hRSTMu3kNtTeSxEx0jN1Ejk1qPZqxobrxP1kM2QhaC5shI7Pfvzry6vsxw7ioqw
ARim8OD/IhYx2MK6AEolZL/ZA4pc3NCUTRg4UY2pKQinR/pQ4LBCuYak29QZoKhg
f7GcySHNX6nLF4Jr0YtsHZI++81EnrNBqbVbARBFmrFlLtuf56ZgOPCKuKD/sMYl
l+uwMx7Uw1c+8caqm7UT808imvHoXHYdrZkUCHe5oOxCywaZ3WXXxjezgzjb3zhX
xcenSL5sa51ieQFnnNjRLwRH4yCZQonhTfFSILNr++MFI9BAg+/COKPNqj34ajgD
DcbT9MCJ9Bf0rLdwqHPupp1jzpdmH8WzJjuXL33B3PaFJMcIp2bJCfzJHfEDH6KX
Vsky+Kqe2zYKLmQRsBk02ZxAPt/yAWffHzsoSGfI6p5Z97wytwViangznYTDhykK
g7mf+eNn0XMtBw16oQw9DtMfklr9GNpFvAoS3V6WBB6KBNbA7U/1sv2+rJC/OkFE
YZcCcpuEYPfRUebRyWIT22T54uuqSpWQwWmEpI2AQrf62fd0r0Ka4Pd19Ve8DwBN
MJ1VWwygApiASjIcaLcQ5dxypsSJxILwT/pnP/EB2DHjJgqAXsK/I7+XEYGGCNhU
guF2Dn4RX/s8ivLNHclCZeIyFNZPGjJxrJ8zISaUWkRGWG4+NeSOUtiIG4gs/aQp
utmw+NSMI7X1UI7blOIbcjK/eCSw5jdFwgPfk88vzdX005cgs8yaFPBn8Ryn8R0a
QIEnAQt+kvB5qrup+uekF8L56/MprvIM9o5znkeo9Y74Ei+OL0vUAyDMfYX+m8uX
QHDGI3jgvjXPnNgMDXv4GwBHaPna2BrmRkipc6agfHIw4sH+r/pbAA0QNidhKE0i
7hw4qKoFjDV6A2MJLsVAjrvnM924AbN33oSRuvjRwJrdwsC+qxpMVYb2EN4EAvQp
I6Wf7SpLoQ7TEmjhJGwYy+FL4aObI/tPptB3cdTlr/VeS0Ga2ztrIF+HX4SWGLCq
+IzwC7xPhY7k6gV3Jrb8zDTNww9Ok65dcCSK3KZTqOV/mGV1zl965H4XvO04s7HC
4TAGFgfRXzeZvUZ9k5g2hKBAO9Qa4F0nVE89Ht8FO9zRQqPqwRuISUTGRadwY8JR
7UFol+dsoOKOVHNdQhNf9vAdZ0bdlxTT1i9nQnn47mu7pe9C208/KpYl/a0n8Pgi
58ftr/n0sDI615vFVRNFLmhVDgrNYtLv6XX5pMM5ErFLFG0Itt8f3esAwpc9X74D
2HFA8jMPYXNJWOOET0O8gO3AMYA0A9QiFxGFCj/8I9wNtD/LYBVUgmkeKyuNwDNs
F3rZsN8ZB/nZp6W5cwk0Op4YoIlEcCHnm6+lxsFdKy/vbgNozN3ODx8yxLLhp+Bt
bhWgwMBRxSCDfQik5KgVK3mzkpB0eaI9MXCDEfY2LIqhAtxARJJ8D13pEV0gODGp
9KR8yXLlLscI66Cz90ihWajlkJnpP3bnYXkcSwRCB3GLxYVhCt5mW9zV7rzTCQTM
WHLVDetZIWdDO01F2oFj/hwhpE9yKmD7W2WZy/GnafQwpEHToz54mdJqje61yoEn
GM+tMNwK4Rjp3AamqiiprrE1PWke0hU7Quwv0JP9KW5nSld456gQkXW9uFAiCh0H
Fb6WsEd27vl8eX2zPDjMorZrwJktYtds8AHKc4X5T1YSUw46g/MoGrNM8jpFYJcI
KlOlNd1QmDz0N0R/dEhMxfrUg86rX3k80zTFam/WErdEV+3hy5MPw9z/KOx1yqjY
9UTdJrPAlKiuD51Bm6IFMv2G/375Vk03NnUa/OZEU6RQvwm2BpxUKYlNgNpQiURd
AtNCF5f1tWT6b49PPGbjaps2SDYORVqh2xvQx6AaD4ISvabiPQl0V6pQGXwOm6gY
Au+h1D8K0YgviL2I6TR+kLTAbYccsWbjNPEJPh4XigsZFdBRAlpGrIv5kCYJLG2y
4CSLdVgFi+lBm/BXLw9tjdoZWaWX9avH+Aqc1gJomW2R+HCVsLooCVMBA6qQmWNA
THGnDvBW9+PLvvoxrHMtxjaI4AxAW3F8LXOOsnDYZ805AePn5V7fBzz9O6B1JxUw
iR9DsML66ZcNvKGjP6FqTyQRq1iUT3dhmWi8HDLrQc3FvsuUnDCUZshOauF/KmKx
z2AigKl514sX/PlT4tPLTDirCrr3G7D6/HOoHv9Pf+Xdq4y4EHqz3PISlNz2FsTT
4mhDfjaXLyAfgBIRuOkXHmpc84EATKDzolvlI+JahMTk3rLbqPLcHlr6VM5U21gS
LgVUqSZEU1nw2UfS2Ohe1RBbin7HBjj+95zrrv5YMAgYNcnOluixwsPTDPv1IWcp
CnqVcI0WrtwPfNq9dhA+7+4Vj7pyAOQOnhSWzetZP3o/un9zO11bIE6cSmIjjiT3
f/FARoe45hxZ1gbfAF970JWuxsPSdg4YnjqcVaIyVpGOC6QXuxjDOqHxGr4JXXAT
itiTzJ7SKKtamXvuC/bp8I1KWOgta+n+qoISWS7iKztSMAe3Xnzn0/SaOMWz+65r
G3v/o8Vk+qFKsCYf8rJ/C6AWiEFesd9haebB6+0EdvSbiaVswGokkx8Le4Y6FR9Z
OHAoYbjT80mFZkAMEjoMdB98hGdvdkboCZJwJ31aocUAdW3HMLjgTnugvIIdaw8Q
ZcrVmEsfyURgoFusI8l7ne9HOqovrf1RT/CMwlogva+r7mq9pXJQZZVr3cKYbFRh
f89NCCk1m3uZL1ZPoMDqezaI5buFirf4Ek4Luwpw/6gv4ofMe5S6NbCKtqo98Mv/
iB4188pyfLEe4RWHWFCHbHNkShzDXdQ2BW4D/g5ouA7pSVSQ8skRnfiKmVHRE4O5
fZEez1WHvWlhPWjcWZ85P6MCcnDBGpCyT0nd9jdnIHZmqEsJr2wq8d+p3ubr0jTc
MvG4AawBo+0QmFpoR+Ca/w+5PiCrOmdJxOce4LJuO/cic7EOmd3hbnmgVSSC/Npo
h+Z4BJtv+48vuAn5P6zVkkk6xv9RvcVQ15D/3gcbul3dkQ69ewDHyPpKHkjmFtDu
MFkLxU0AN+Vp4wLxsMaZ2bA6eLCkQ22O//i2V9+Hx86NGOK49lVGxrx9OPZAUTSn
QZ3A5qZNCMoeKiLKnHaOZqfIe0lznew7nrLHICeNba1yaS6Dhcjxb1bRorFk3QXT
kr+QsuGKLGtaORSdneoKTqEKSqI5CM6ZboiaeLd6eW/R8EeiAt9QeFnDABq2hPLm
qwDeso2FSatM4o/EdNQB/b4wLK51guMsi6S5SLVDKEara37KjWvIUscGhHmyUsxQ
YED0hal2AHio7PcpN4V/xjuKdDwJ0yZIP4FhPSIo+qsln/gauiS/xsV1t0F0vPOV
fExlI1HCScQrcyo8vzlXuiyrtSyrfGGGkWRYe5p27BQIySjUqVx1J9y5gV3iHODl
CkZ3sjU4H0lFlLk76wpUhlJNjy/rLMsc+raKC8CK8UCNqRCP5WxWI93FmMyV1sg8
MHPDGvRd6c1SQa7mCQZuT/u0shsk53ovM5vHG6akpzi1lc1VdfH7lG6gfPHgswCy
dPBwmhkYrpHPm0kji0GF9UdZKKF2Csok+uFO2QzLL5tOai1VqbPJ3FrU68gEyCFt
RzQM/WWsemHAewNUjQtXp2hC57IVk3wHMgt4yKSdc2Jf7GldcZCQM4vi4UIxLUeG
bMZ6A4RliZljvLRU9/QstuRD7p0+A3ntprKAI1J0P+L58ICsoIFhKB1q23RPsAaq
QPGGpTx8l0CrpI6a9GRXPHVjNxgpMZEUbuW+MK8uplFbix6YDbUt4Hhe8k3jrkCS
sN2PMBROtZLdTMli9OJ841vw25ZYjMLoKx75uYlh0NwKZNUj9k+l9lMmmGf8mFk3
f3O3VP08gYatU5AKrAVgpjJSaichvuJI0KYSQp7TspRCfj41ZitrcnP/JD4SNVkn
WuYjKKdKbWWqmsgQWXJqKpcOhmb62n/JehMymV6EHJ+28IDsfMC4MppGPbR7V8ui
2j7syoLdWQKW8fcbR1zn1Gyf1a+T0Mv1qpdbJWw1ydMrPzcgyxrfvYZHQatPPuoz
5AWCC+hubilpYiimf2rXMpf2FbVd02Jfe+/evUXiMig6BltCgPpGZJE+dkfoEaz9
vVqScxi7W3UR2nDlBwj8fiviSsErd19MbSsbzua/kFg3F8W37/CbMpf9nkpwOleN
GjT5U+N6fFaSCVtLHPyORtNQ2qPsZgj46r4VEBq2lcrZP72Yin+4V6vuVHQG7a90
HSitWmPu0sJGXFSMsUVNytTpzSFdi2b/qFkqOPWy51Fb9NtH1ZAM0SdqWq6q4See
/zI8Faoi/fiapQekm94WZuMVmdGAvkZ0Nif2IggOJL+QUD4aJuxbWnv45gAqclXL
JGQ9Y9hIUXut73cix6ZX3nnwOsAwJzas1IwP0WABPByLQGQE8s7D22E54bI1ihSK
sZLhNzwe0qvUeqMcEzbNXQ==
`pragma protect end_protected
