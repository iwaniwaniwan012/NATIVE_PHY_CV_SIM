`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DK0j7A9SfhxMU7KHzMvmIOS/0xTnyMuBK++BSFtApXJS0CAmA+ZlxRfuvM0LuqsT
ozwnToOf1NwdXN/vJ6vMWdl5yQb4oKzQRPatA0d0gMNG+vIYlCmiBDj4bXfum4Zp
2yuOj17sSxYkvCSWdfGa5msbLr8NNIeaIkI6xOgYFkM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4688)
H/OYcxwDDtk1mLqOxntawdk1ommguJ5jg1NPPy1uhB4sRT5nidVPV/3qgJ+SVi7f
YCDs05H/S9g2Xuev6+CQ3j5Z+o8LifyfFLYPbNz2pp2Nn7XmOP1rOIw6hr7+Z13A
6FTc58UszgFSYMh3IVGXf+WyGt+ndM4mps6RHvYEXJDyS7NseLZ/LzmI9zrAneqU
fx27Bznz53x4gDh91lTwITP0WPKsRD0fRTpGFLAV/s3iEAdysNpbBiloojMYWvHp
gzgni1LWRS7f/cbdB6AWOZ5bIsxNUIGJZlU7cwWsGlWRJWr0YH+ABPWSvmtispRc
ZKyvjlnyNAsW3NsnU3fZiGaA0mPqaKtrMPQwzmrp0nGMeXjfURaaNGmD2Si6AMqr
WglaA+NTNvt1dx7JbDApm5JNf8XsSH5m0aFjSABPBg0vJqev5KZe5Dn6EpdAxG6I
QaVf8rCDU+UzJREKwN/AN1CRKgGH7LXBRiQOYMpKdJJIphuNjnZO7Qy6vK++tEZl
jhr37CUSi+RVQ47vjN6NTlQclKxCbWFGpgv065Ul3QdC5D/vii0CdNtu2LEINW9G
ZLRZHDzUPknpH5ZmRTf3xqocDyl4SOoB7Wra1kDBrSVjnzYNkJi4D+154AqPwZrF
ZIVldf+xw2kkhDgXgr23BnW51lGswt/l6dq4SkLyzikt7yR/ZsnjKG2AE0jo6q9I
LUotIj6AU2l/0UdSXm26oP6oPIP+4Tz3xGLXfigVmUDZ9l+WH4J0uAUi/MINTIIM
kanwdye7ZREn5hg3wlGabzinE2oDyagmNgas/VseX7vcvi3iwX0fsbiFuVHHfM6y
u3T3sxLqsLSb8zY5078d9sWtYLVsHYkafyO0ZOkjCy6eSQHfKC43Tdhx5k9vLP8S
onOTUF3rfeIWuxEs7TLfEG9vuvipPRD6isMBuVelnvztV+/wBU8b1FoKdCJGhXjv
0NhZff1yJmgD3pmnc4aHgqG4sOyUBugF4a+5GMFdg2NCW1bRQVY916lFuXEd5vnw
fzW/nx9bPw4rX2BiOrYmTUYX0X4tlPntmR1/xqW9c76RY1z8mMw3wNZ3SSzDCZAN
PXCvWFQwGcwO3lFGd4qaDWVoPL1l8hlauFtMHwdmu0X0PY6R2FmLWWdLV1Nvi6nu
RvMqLGfkAD5QT5Afm/vBnaGG8k2xPCQiGNRdPJLRjrd+JCUeydXD/s8UN93kanDW
uSVM6vk98xs6EAa5iELS2lunX6YhdGGpxrR3o6snT900S2iA6XQBfnYa5GJ+eSOH
xmj+2pCKF8fe+f2z+75CLg3xaCrr6zyYtb2i5bdVRv8YrjIqZ8sJZbQtReuxSHQR
IL/Jm/ZpyjYvwD2UrzEEQp3mJ9mwdQx8h83aDlRV7tYALNcZCepOUL88b7vrrACH
Y9OpwQj3TuIpL8avo5x/Nbe8ZudfE6p5QsDCu5Elch6J/HEPQPXuGTfFGiVV+oRz
f/SipPZDL/F3v332IAUCzHbtM0tGsRQRm26gqZlEvElsq6iqP2VYeDKyXcDtDdRB
37XsizssKgIZYgEceARTOdi+l3KYHC7ZVkGssSnRvnfVx2TxQcqoHcvqSA7Wkinf
fvqZl/YuYHteb5MINbRi9p7VU7/dwY2/Uo/EF5n9nEIzusQtwOYUDy6O7oougLNp
sXFY85WavKSVvOFDK62999iTMbu0yyNbEDi3JCNhPdh6Hyov4avXrMcY+ssG6XDM
3O28WEghR1Wex/6BHQsCFCDJjQmynLJb/9v2gMPBRjEAGqtshs0JCDDSREcMekXh
4OmPaNxIzyJ5zSiiA12uLMGAeN1ATiTaDuE3YhMKji6X+iazchCHAPB3SA4HAfrP
SuifrumdhpuD4KfxA8Y/l2Dj5h9X42MXJIGVyKRxqIGOdRDjjwo4IihLflf+f1v0
X3D4p4DP3NRP2gga8ZB9RH9UUlSOFOzj+Mz0o4HmRS6Kqhpqj1uFr30C/ZLeWKRD
W58CTGohf3GTEmbMFOpHRgPvEsV4/ZkJ3MFeW9ldIGQxV2yoJyVYodjpTwDDLA3x
DmKdVMs8s8eXBQMcbgnpq9QU21QboMc2/XpQrPLaqVbzWjy9uPDbnEx5XVX3sREC
FusjaUFQ4ix7p+Pl3G1JD6EaXangd9B4AP1lYwNGjQFHnxrePZ+4XOlDKSV44PNK
m6yT+oMAORgCPDiVmISGwBsRK5/h3iXjAUulzbdy3PTNhraoUj8Cp00pFTrlBu36
HsodAariGJkDVyw30J3nLZGdqpl601IVQ1rncoun4ZOEcxCodXV6YRnYxl2NMDrx
UN374XCwqmbfXiZW6mMngOigu0TGnScKAM8qQVE5LktjIDDFxQJ91nK9vKQJVLYm
D1a9QyDxaiYq0IegFXBP+a0VHkzZ5NA20r9I5XCLSCQoEwm+NN82Fq8iicHaHwmi
f3/Hyzvz07JlR70AVFYOwTp5TBL2SYUeSacuPvIkajI8sbxWnLtixlLnqvxgTxpP
ZckKq3/f5ZZtLy7gpXJIAJBS7GnGC/OoZWh0G/NMCSQAtVgJ+rtyE43nl7OY+tSI
uu4d+lOEd+SPDJWZgejquU2GSBsQc/zTHCjRsskKTkb0gyPu66rHg3M8yTKXeedh
qRg1V4nG+WpVlw4SnoKYlCq/MHAeABYH/4bldBsvAl3x9b9a31DbnOx1swB+xey2
mwDhDEPt17AHazaGqfjva0KWSFetpESTmaabHJSqwTqx419LpJVL1/vi52MFRVE1
HV3RATesvgfSisq1unxipIzL8aLRa1Z2fk+UrIf2vk0Q/VZARvlqj0WQLlTJw9Gp
sTprlUMfv5lN4HionsUuwUojTJGDkTs0eGnOm3f2tEIN5pIevSmVpKDodU6byYj5
mm6EqSehcZ5VwGMZ03R7xY1pmV6C8THRpD23gZAmM12cZ+x7eBHXvqaRnUoIW38c
GWWNkjXt2OddHomKTs5aEwuTg1u7SL75OEUlOE66q56niiWcB9O2yLojF+y2U3I3
DZ1+34H++jbD4ANYAFXnq/l1PZQSAy80crvmawNDFqwpfpA126zDKMY2BfUPW665
JlzbxBOHhY/cJEOCaKq8zdFtoxkIpD0tJ6alYF32rOQkdF3oq9fnw4LoQjIOzn08
xGozGIHavFozuSe9XbVgdseKzD9rD8BOPP/pj7HEk3X7gg8JqfvVWa5YJe1xhnla
txXOrqMJxu5tEjNVaPuM5ntyQfvQlaEz2yRa9/4QYLPaqXQa2HRgI/vItCPMBnsI
QWUSVXxTN7JMaP/gsPeILyDY9STFKokKv5HzQzqZ0PORWxi1J+vizTO+oQn5VphF
iSVxv+42pyPakdangbGysSdyHdp3kQs0t+eduOKO/amVvjwqPwREAO31yetl7hMM
BZAepr9324FEGvgy61TnEHu4yiZkGtsuVmTqLEgbIyKgjpjtV73zPSD1VoVy3n4V
1gKRiCIloF80eGgWDjvqPCWJKXVfy4x4ZFZXfWi8jF/62bjy8vQYO6zfUiKBvwWW
+7GdXldO5t5lcBBHwb8FcBzAXzv35DXfa/WBcdr06k0IPc19uwfCynY9AStn2xak
y26b8VdwMlV+qFaCvL507rsa/gn+rIQhWNr1o72bdGp2P+Hs1BSsCNoT4oLCG5t+
AEQ5an6cCUf0Q93JEY01sWmopjfnZWFP8Tjj6RVOMgBa62sRH6K1eIZPBKCp1PlW
JwsAMU1YIJ2GUcJgImMsZiFxMW1E2lR5twqga8+UnvzFfTY2g4Z3sZgaqILWseQT
yS20kjIY6pOrPnBHuA3na1fLdRJlchRv5q0tZmlG+WCxt2byVqhPjspHqREB9ZjO
KmSRo2Wem/7J4+bGkfwTobZI4r3WVKyVx/Kl8OC5bUiOk6aVzTOgrN0rmuZ9cFQb
n0B129AsQmsiyNTCzVV2VRhoTbtZkVB8esW/40BvbtfxnGddHNPuyHjsjpLHSFvx
zgmM0crpvQgRjdbM1zwLT0dJhGrXt3czQn5mwGhwZ2aQLIssygRfjfzB7oNXAwxC
j1m71ujoU7Qw2Je4eNvP+QV+r1DEkRDYHw0U3yRX4Ru6ImkpOjfA6RzZxWHty97Y
K5kIRUg/Dt7K6+nMf648eQntYHhyWnw4RYCJ5cfjrdgP4L/im9XWO1ZNT6ZZMqzK
ITCnwUol6kb37heK7R+F/MNizO4GG008OUQoEu+mLFYgVKXpXIJ3YPN7gHFs8GNg
Q+4KsM96151N7U1hcp0EDSMZbJ01puANoFDjOV4eAOLTD/N3QcANUGqBGBaP+8uJ
PJb9WcPpLC/ySmw/N9ZH9b62HaFEPbPPLFOZlCSv8t+avZ4xQCGrPuZKW/VZAATi
ZGPwi1bj8mqec+zbdPV8ifbLAzTEkhdSADIoLTyuyL3ZtqFzwGTa5BWuIRBasni5
xuv/gnTO4nBJBW+wjPQJaJDpNvXV/emXf5H+MGg20dD5CSgJGts6shDlQ+LPr7CN
2YJ46AUJFQ9fQgQ5rr4PFCCtcJpLD/h1uBRsTca3S5/pivcTn+Z1kXN3bO187CVM
g+SmnLPDEibRxOEHTYGZ4Gny5421wcPr3vCgV1YqhNwc7B+LnB/gfK3rb3cQ3DfQ
4AO5pn2O18PrVBTjcTa1Xmtk5MGtBazKseJKliQpeHWXro60byiZPpuWqV8q+But
Zt2YI0zXIV7iSBzXTy1YUytAwTgGd7B+lFoVeHnPxBGGqk68bJZbcztvqgAU6KBh
3C861rPnODyCRY1LC+ZYCNcZTbZEmh2z+RWJlqbpAZJ70j+zdcnu5LEa/ZnYsNQi
pCW5DOKDpSlLsnqefPwBljQXxK7YmJLfEZ07O7HzgUHx/N/FULjmhfje0KGaNlBx
94S1x6BHOHVUFYBAr9toU+JoHOj7iFrAQgKTQAV2NCM3T0cH1Abl5UgbmnnPhJsF
3I8+B7SfbA3XySlQS9jnlFfJZKEcezEphyL2apUa42bkFsVRBLJq+djUqFX7oWoA
EHpeHdJSw4pNfxzPknx28IDGCC2Puv0AvKBUHoqsQN9wUvBMKRQMq775E2/02sPu
xllOtfiJAiLgdBosOkfYpcKsylw44OuYb0SwlwIM71LSxTsDa2qmJ0dONeylC3LZ
DlOsNYhkWQAu5ZHpZWlJhP3EUeO9fxPfz5WzmZbf/mkQ8GybeAvE2SeOEJG26l8K
zgLafxHt6mJdXAL3WLiFCaAUsjjOvoQGvCBsJS5roS9liSUFy9dDGPtgi4smt5J0
RxA/ZeWAbEKbgmzelmzMBVxr5XCHDjkPve2pP0jPP7Rh/hZXaAHNV1+2S31kaYRw
6b9fipuFjFZWpw9sN5tOdmLdTxE1NoGU3aj8fDndC8RgHuYMHQMEg5kXWeAWDBbA
bWy+Kd/+yS/5QimOOvW+OpwPiNFkAIWSF5DXK8VoV3jpK9Tu0NX4jx4mzUOyFLxy
y5lXpzQ8qIAf46fKBH+B8zPjAAZHcQz7C7fHeLiQxSYWbivc/hdRdQPEXYzpH3Hj
JBFluz4CAqcJmJYspObzD9lHUIoTX4INNAOdJlLWcbaoDkXf28dV63wkOJFxgvF5
oQ9MSunfsWsoG3E49voEfY70Glk1vaqeZ5NLmU6kzOKdBESERxTVrP+DsHd41GNs
yTaaC8gppfyXvPevqBs5E/iTo3u8ZEdMuxf1L9FmSjWSQGkZyqXc4XWamf2UVhBt
5iMWVSkv6VG4zOPmDDvsceWWm40KXWEReZt09wFnulsuKkyhHYamTAmwXZ3ngz9c
vrpTorz9zRRdAClrMt0Eiw5VHpfL/R+BSLo0DD2+rMVwULQca228YZTfVKm3G7+p
W3XjDP3B/5RKdwitPBxQzpzq6NSjGV32YDXn/cpfrJy7hv0tzIaRsL6mz00/Ysge
iSvmmen34N+Cmh/Jm6vmVKsQsvqzTP6cwFCGojv9AUBDikW/1rh/hGey98K64pc5
vOifEv2AebWLOz4oFNn6/p/AOBoUbjc7alJ3X57CbhFjjy+/NRyP5/uSHg8iJVt7
cMk3M4GwVbbwmI7UA+35Oow3ZMHzg4LSAO7tml84m1B88BnuWec2xnQDOK6oVnPK
WBwJA32H4N8/p/GfTIeHe2j2BZZy/q6uLNvdR5XLijXMU6BD2fKDVFyI8xS/wb6V
l5tbi6AMSU1rAXJKDDyCJqRA33qTHo+H6FQryWDgZ4XkJX+bl73IOLqoFPijiYei
dJJqopxxKrHBzM9QqD/HNA+1r2t1zniqN8p/zPGvVwM=
`pragma protect end_protected
