`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OAYqYRBfyZgxiltFY+vR9wP4qSWZgRR62CEOFmvz8TaK4AWNoSuJscM0H+Ke3F2P
C0z6SIGsZqc5UInzn2W7OvWPgyb6luRDpzGIezlRFqohZ/wfn1IZ7fywtVaoBVFi
vTw6Qq2mpt7wfLD8wsYn/mVY7swtyS479omKoSdpEVs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19616)
QM3d2XrhjDA6AvTsMZB9c6ohRfZfU3qWotI38jDbVzNekl2/3phYlvsTEUYL/7/k
94wh9HAolJ1sCtZV/UXwdZ10uCBGDGDo3uiAb9KSRfXlARFFLlWGASm8PGh9K2X+
KHBaLUGgAdlYi+6IUfSkbb55PKyEKETR03tOpBoLFuP9HGD8CwPL35cZzBNjCIDC
9+YOOqK9JhO3iaHcHsk1FW5qFhE9l5M4j8aGDn7bdHgaGfn62410acPx7K7cuO7j
m8nySQ3Gc1He/0M4fQ/Ym8y1Yd/6lwaTwOSvuRXB+SQNXyZiQi3Vszn5ZnPzmjay
x6lnpiscm4PcZzDiKRV6t8KUz/CoueUhmd5p7Wwhnbe8F65Nu6mnLBpFcZsCIt8h
SlShv69CZ2jp9izHOTBYiuGgoCziMOGa4OAiM5Ac8mxGUKCcfOQDXDMTGBfZY1g0
3JB6FEyW5f3a9R6GrIYaY0NR+kr8oM3SO8IR4ZCDf5HoSWK4UGhosnn/ao7dTSjm
L1hUfsw2UQWXsMAM9AQl8HMrLDnYglPC/nu/NGaPgTDDBDPYDg9dXngE8sAEtnH+
N0HuUmvUt+J5Z4tO0NMOdlSNaoPFVhnvWeQZ0vhMmL90fxiRWsNf+59z2Aso4v+h
0XQg7GR//pe8YBtJTxP8d/8MrXQjqzEvaXZ7rG5UqB4JJqDhuObRqHoWbHvXDTfT
UluSM2fxi3z9tKtzeb+xz9fpZZ7+UKaAi0iFCTObEpIppLeBdxj3gYs3s4BVlyMQ
u1xWHkV7GZmvZJkHrRjQVDDxhI1YaoGwZsvOy9Q09WrQmL0vUXqsEU83E2entNFV
1ngjUBjEfh7ewlerus4lhDL3lgpNnU1eVSeck0zzQRxyWdxyU9g+i7i8i0UKn3qU
S+uGTwwbNRh89jl6NbgRkhJZZVT3yh3BvtjxAQi4uOCbI3ZLRACgZDQrf8ot8n9R
H8qTCQLKuoafioIkNO5nRpc43Qm1EJuOa/tckL1Of4Ri5By00GIC/ZQs7P/36xgK
H7e/mU7BWDZaQnzFARVoar4iw9VDsUwrmm6q218I/oWpn/q13NjlHJSE9DQyFhe+
r+A4tdAh7mDG6gM5kq0BK35NQjs30Uj0nkTXoVVHrJLQNBcVfTxMn2Pg6OdF0DNY
X8pnGRkxs5AIJS+9b1sinsYt2boypy4SO6MVabg0T53PGQXvAYLJTbACOLNq3tNd
CrJgo0z2kC16HKOzJsvhdqNMOY4jaWbNJ4MB3nEeWlm88S5PLLq/Mb9YNKplN0Bo
oSVYWpbi8ygTIbKKkbBrmiUmCbQ3933pUYSJuHQnnKUyWjP+wVqMO7PuOY2DaVql
L5VHoqJ8SFMRvFWSAtt0w6RrKDMjzcHUH0TBd1kHFQwId17wrf+kvQf6oTXObj3s
9zAs0506TcluTvwf/cu8jVq5/L4nZ6ibWICLltCSFSSnxhGh5jUbRSrqOr1Lmwyp
hK04ugBgFiTpb5G2285Ojnzb/68YraL2MPUqyX5YPge9Y6PKBHebpHHkNbXLR448
viqxGIBkDf7EGqDey3eaPuRVczZ/HAMFIHAx3/P1Vor/cwOM52y4SEPmm8OOAFIT
C2RspKIY0PQyoDgSBHik2jQFPJ6X+vjmiOd8XGuZw/Se0/IycTNsxUkSdP6B0+Bx
HI4hGl1OXhV6dRK5eFf7zt5Bs34+vtd0VUuI8AS43Ug7OgGQwFx4z0wLuFllVWwz
YTH6E6vx5BV/+qcZEoaYQq66tpCbaL8mz0hQu7rytCRfiQmogD+a5e2cx3Kh7FPc
A91sxmATfpQpBQnre9e6rW1113lDlm+y8nd1Ai5nVAhaSfxax8/oVBgXRuNlQ4R7
6oyO8iz5j09fRuyxP9y2o92FFoj5W7ahXXS6CRtQu/8DXZlurgdqL/QxHbxzwfrs
NxIqN4zbb+bPTVu5UD8yiGzT/fNz7Mv8f5grFZUBCp8NY4uaghgLM3JdUozfBLhc
Vhghox6Ag3PaZKOA83YCQU3uuaBjcN3ssBDYIojyw54SplT6wXJ9Jezos+P7prdi
lc6plhMp1bNCrwgqNiPLms05IWYCHAE5eboD01GbiILWN4oGKSygGXRt2k66sKNI
hFg4V3uO94lF54r2Y6XAUtJZKr1qWcAuRsrd5cq1Pt5gWfNl5A15d/x09eYvHL5A
3O9r1P0PjIeOcMzcQeYfGPb0/YdryH/PzswztGWJL8pQoEJWVz5zjwVJcLg6/R+g
CeiHMO26SEbYj2o1UUXoJWva6yQ5Vi0QV8JsjApu1HLvzBWgA5GNEA9/n9d3eij9
kRdy4L1DiG2NlXSSh24+aUVvbox52TPCr+wPBVzWtPd7g7sC+qz+wUqElw9+0l1z
C/c3dkFIfDnJVU8xMa68ZposFC3juz1v0DRpRGl6Cn9Mxi7VkaOHBHkwwNiOzDLU
y2Ydp3JRNig6t6QVYlGzuy75Zg2te3KJkCUJieFCeVkC7X3O4Ft2tIA/aSCtPUer
0XA7RqR8QZN/KwddnNciZAAeO1iNK9Q8VGhXY5NKAXJz7RQfH9jecgz2Qaa9ZNQC
s+4hLz2OAyn2QwZSTdCPq0INWVtqNTSz8kngownZtsmRy8LoRMWw3RPsXbFrTJaR
EWFpQjcwHbHoAhHshZFnwmxC/v0NCUM6KThWmzV01E1CgGJ7AFiSyEFl5rSFpx+n
NECKngs2TlOgYXnUWat02ceGh1TybEW6UnFvX1EYlPJrPIbo/cnQHUr+NC3yTf54
6D6KxjI1F3syr6FCVj/G0ZV1mwi/FkHio8VfcN83YCMSUcRfO2QEm6XigKid7uvz
pLkebE5Y1QJjA9eLJHmk8Gd7lsJDRfo0w4+WShV6NMtYnXWWydVQ/EDDpnUaM7gZ
tyrRXj6ZZQzu99/DLmxGKgv1yaGbsFXQc8OEErBdXAmQpdnGQohhAgcMpwp65o81
DfwbrSIoEu0UBMi3eMhJB8/nALmbMio3B55RrgkGPgeFhp+PgxjICkFD6ovLOEOq
cE6WX0sDdO/X89YTZzjbNMC3FrsczOzv/kt2Gfgz3ogwMPcBtKXYPKqbG6ljDMCt
kXmT/ZMkKWj4LNkH/uFHd8yS1J6MVei2eHQnoDO5jphDqyNd9MEGN77wpvPQk6jE
efuDy2mpfDjnlD0mJyq6n0owjBAkFbNo9Ij8yNTj+nbUsMN3fWxYlHK0aul+61BE
NqO87Cp0ACc3U4Py39PIJruWiTOROyrbnOcm3P4yVs14Rt/QGA15vzJ+Ods83jUv
kiCDuID0NbSW6ztrObWL7LqFj/KpeDnf46Px06aPhLX8jaDii9w5ffakYsXfgw/K
pTJ6oWAuoTa8LHWtA+yXvt7l5WdZh+WeC6BKk90KjtP1qt/mhX5zGE+Tf2D6y3IU
soD8IpWMtEPhBCzWNztKxEy31JhoJQN9Gg7LN8lGBtnJIvrqjdgTLuGST/0a0PXw
5r86lg6GPkbimme4GjvqJ0TZlGfPKVnYJjAu3ZLfEePzyyQ6Zn9ZdzcFq+wk7r18
JyG+suefMH93J5/6bfIsiotn/POvUr2jMzW0vTI9foH/3wiRrYx3tj0wdfizOf+Z
T9Z/8A2p1tpjPtyvPDhNhyf+Y/FWDBGMBnzzhRzu2H7DwLaeJMqCGF/viQfiuELi
fMtceQPhBIV4d9f7A11ooFSCBuWiKwpJn7DAmEC1Si/6fK5mW8GUJJowdCKK/7ZF
lOXyTRePeDEu5h2IIuafj/pR3DaN2tb8fFFddGytkJpRcpMk76aJqrWTt/JUIXVF
lW8lTL0UaURrBfq5kt4YWJlrzl5XX+gbc9G+rb9Eud+bo01uEeiBHTOWbJ88OTdH
/FKIxvxQdE1XD3cPBFWfSmyVK7cXq3LyB3cRJsAM9jyFX7ZAKOCW3gFy21PbOTar
iVR5gEKAjOPDahz8bOBG7sW00s0Fi27Lo+bnwcm/tqm5EbFzzlskUyfbsb7WJzJz
/nQ9IOD7hMK4tAHSSjSz1/qvk3OwqftyE80cjBkbh1KZDALQVdAqhYcsMrANSzKb
Gs3ZkTFft/jAwCoLOgq4DzNfGPMKQ+TRFFIqcEYVrc8tD9Byaydx6hNVVMVoHTLo
rfHWzxf/h74ALD+rUe4cY2p+3W1U7sFFgF4OD8CNT6Qe610FjHqb0xC3E0Uls3iS
eMbr7SIXBtNB9eVe6oLwvMpIcK4V9zT6/3x8aX5Xch9z4hD4RlY5QwRSfWFUWHMK
E60+vP2/g2BEXSSXiJu9kCE3cBRZYYKRVnDGbCz0cexXh+Brl22w708QT0A/16Qe
HC6/vDer3ShG4nr0M0rQeXcK5BA14K/uSIpTCP7gW2C4AoVdId3uV5evgYo9YqLX
ObDhC+chuaPEuA0kUCqBEojPC/XlpGkiJE4yVQJ4jReb+vAXap7uYOJIFilc6ruT
sdSG/bYkpbPhgF/1evj0CKJ9U4uyKyM04pg1PzpumR26CNgS9uH1gJ7rkkE4akbZ
wy7qa5jcI/mbuqBXMxwi9rhIXkt483Pb+8CdEh5UhaPIJTE2RTEi6CnKWiz/zEkI
kjuzDQpJvOvW7PpEfUM5zPGDbTseYBQr6koaXNjxFn72tnkG9ElxjUNDDz/rtvoo
coduJv1n3+KyfI/I09ArMN6F0HKXjOg/IKefCHQ52lzwy3CH325gtEqEqo9PVKF2
vO8h6bld1nw4xZ+fBIiFFfs6Yh54PmcNYWA12+/JMZXbF5NJ8dttwSWHI2G0EMMz
ZS+PlLRvWy+cwG8yQthq/1B74QFxWJrA5cg8hpu6g9WJClSToEHZGVMYHCHn89oK
oGy4WOnUPnVSgIbspCg4QggzHk2EiiXu5dJ912RelVinJZtfzNsBUIRWtlSTzLBw
xoLDEQvs3glicpFqnD7t7sQwbDFQo942MyR5nCZFGbWNKhkP0IefypkiIzn0L40p
6eqYk2GBcLPSe0cLg27ZAA/qnj++F0a2H28h7fpoxB0Y7duuadEz/1yfv75Mj88F
KLh8ZWbUImwAglzQAYGfjbFy+pQ+EzU3rhazBWuhlrAgiqWfYwT3XRo+SB0bDLSp
SMoWACVCAyEIdLbChQPasiCdVixRZ2OCPBvPA8NMwyAZzMIFEVu2I0qngdGa4Nvq
jQUOEf5i9q6Rhpgzg7VKUo55+Rd7DJHE6e6fUCwB/Q+Y/BIS44zFBGrp6L4mc+sJ
/T3ez+/iy2DVaW/bQXxWjxU3q5i/yqNF8AxzjqowTu6+W9QBz0SdvP0U/uVIS7ha
wxenwWAHOfRn8Qd8k0pyV7nmhCxPhuRrEfQh8AaUH/X5j2TeQtNkurZuuExbB4Qz
eSf7BMi06EOlmU5QRu5AIQN1Vbtp3FWI4vkTZLgTBwlElEuhkwYfdc0m33pcRK3z
mFpPI0L866yKVtwCZov2AvULsoDN0HEP+NBQUDzjPVPSruJw/iW4Uncmf9eYrI2s
h2VNPOUOOektgWq/Vw7gWFxG0/nAlJa17+avZx2Kw7NfRwojM62Otjpk8nTfs1US
TquZl6l49X2m68IvdbTsaEkYPM+uFYq/kQVbKwGEXy3J4mgQMlRr3glXaklBJo86
nz8XHOiyOhq80v08rfVQoXpf1Wbv6RVHBfWAPcr+QWRvRqDWVm14UWbBRpAF6vsW
gDxj0qkSYUdbGsrQD5NJ/DilDqf65DOQUTfQ5SMB2Ev4o/gG6Gmokia17HD92lat
KZqBAFNi7iKeetH5gZNC4bHwV41Vi43ELcAZiyXqJp2IDqaXQIAVmcJnv70Qm0BL
Ipc/rZa0xWMS7JjlRHeb6reWpBgq7M2qOb3e5Bn/G/HVtxgG7MSBcAj8HSSGuCAR
HvEmMNP/03ClJOZPBUCPu0LwsV078pgCPKDm3jZ0i+0BMxWxdG7LvlGRlvVH+byC
TPxTRCqWasgqPVSOndvdIZ4KB3/VvqbTns7p39PJng+wBpwN1Ni1QqMgw4PI8/WD
4XR8v4STZpg5rlo9N6/xECANDmt0Rgygdyg47LMXrOo3sT2Lav2xRdSQ1o+kQX67
CyZaY77bZTFfYobwe/15uf5uVqGmjwMoNbu4UYey32yk7bqUvpHR6mKDFDCaIAay
FOk1HhSfug4YK//XL8pO+KXfl1Du3mtx4K1FqSCA1MjhrS7wBMBP7EeUtE0ATRwd
gFBQWvhjFAO84zUFWqPjJitAJw+JoO5qRXQGpWBNhqxtxeNXxxn3Eyq3I5BOW7+J
6US1P2hETT4+587OG7i9K01k3v+VGpNSwsQTs9R/EtBlf95xikehvtXBMmaNMMEz
wMaLI90Qmenxgc2onKTu6gsG3SK4yh3+kjThT5zB6qQXb00Bjr2xKM6SqDSwylsI
Z0Z4kJQE5y33mRFNVUBS0stI26wiySVN14YH3O/jrUPAtpLuNHya3tHcKjP5quv7
4T8dc0fryViR0OfPGZJVcZKumkDBekXMue8E03HZTsaQPwCN0eJcBd+b1p2wOML3
pNbywXbVqc+5BX62WAodIzQ+8PwDYuTirAdaOMVMLgQaAIDQMVXhFosNvmpy+xj5
vYEagJ+0lPudmL+ZWRux8EY/cHXWHSSX8ySUzfuCfT1cdds2MCOXUzS77oqztfa8
/CsNLLXJL8Bz8tvCL7+nEBCbsVOLS16MST9m1g6Hqr4jeoRa4UiAdveACII1Xajh
BWU/RFNXgWoHa2uPAHxIYhOGilzBWzayzxLttVVyVtgLjuMKX4Mujg0jOrlXGEMI
hCs98YR79ThHS2tvsi/DCR0PIonKLB8KPPePglTOBvUJkne3/T5POdveoXZrK5ey
Xt4jssHfdA2YlQNs9XFON6ReXN5fKYnSB8Y8qBo3y+Tv0yKvQUZa549Y5TZkKK7L
e8TkImDNxArjQgB08K/0d5GxUYGEgNk7DOVRsDC1+zDAut3vLmtgh6pl2FQHRQBv
6XtTOx8Q37LgSjrKImxpZhhbBfRJlZMdX2Om8PjRpjRQ8PoUTzeNIdUccobLL1G3
OKqMCjm/aKIKszGbf6ngGdQjd36hrNyyk19j+eIeQ9KP+Xn+2/h5sA8LoxdcKg12
ZkKF2vHWD9rz70wiqP6BBxrVZqeYboQxaevqL/8JvFGdprANzFnzKNcAl4Q6s7A1
9ToxYuNAp3ztkirQeHuSIp4+xayILsQ5cX91coA4lfi4ywl8BfjHF69gNGqtWZc8
YTbzwDXYfyNeQvbdLFR4PMZRnEKW7mkGfLaFwpRM4y7NP2jM5HUiPiXOOzNdjbeP
InTrVF+IEvD2r2vnLu2G5q9uCdATIT+sEdZWE5e88AiLMcJ9p67RyZfmh6RWl4c4
5qSi4RU7BEOJYJ52fPXuRsaQzHee7lrpWFzqHmQYRxSWLqRUVXk/smLlr4oFtzmT
GazDm2wsvb6khiLq5a5fMdddurVnGLWgynuZDhy8XgqTXov67IdwbpwBNb22IAjq
qxolqnwFjnk3Ux9cIuecDMpCsI2tPIyeToolnRHBTjywnrhmD2NsItyVrfSlwFSZ
qoAwb3iFWhLQB4uejE0/+fL6bcoP2wtI3iJmFTTpNRAu1pD0Xoq5bwXf3Bp0hx0D
IpFlgWJkOtY/e/Ov4PAxeXGRZRgRraguoliMzqOLCL0CAnx6sgUyTdjg4qBoqasb
Do8qsXtEuutOM5q2Bkb046Wqu6h9tm/sJGiHaHBcifOFMGA4qi28Ovi9HoHr2qUL
Vt1uD4rUUv2Cw/bKqsbs/BYssOjiA+Q5TfqFVnm3Ywm11U8s7bQY9TnngDicH5PC
Q3RhT9gzkWGAPkAgk62UZ5lvJL5Tm2TrzTyToCprw4QGztB/dAbB+EwRp10DJXmx
V0FcF7HEKF/Z8uHXzzacKu7+6QVxT5188yIKuf6ssJFsFYhNwtvYLbq4h+mSH0O4
WEQhWlAF8pzgMwwhRGEyEIAPYQtg7AiWqA6/uhXoLNYa8hwV48GTa4qzyVaXL9ap
rhSQvWeFDgxY4voaY/z3abYG/XHK7VSWwv3OCOxnC9+FmvT155DLrYMABNPQqITt
9choTwvj3G9QDtP6J6hVLiTtGM5zJvnbKvryYkgwpLZKNP6o3ivCh/vaw1cJCa+U
slAFIxXzvuKZlBH/2s90qQb03XG3bnFdg/X0kgG1s15aGBtVUa/YFhwO/3rNrAXq
ZHIjZegPwzI3li+IjGNZzbeTtx9A6UGpdu7UfiWgS010ShCuXStW47hbRXE5Z2AW
AIJ7FlZbu7Plv0Qd0cUXj6mEdpyIxRODe15Adh63YwmpcGE/HuHH+0a+C50KVEML
BXWSgPP9m3NB2qfJmGtUPn9GMMbHFTq8J0uscNmx2RBvHUMFUc1wEi5mxFfBacxQ
BINsE8pkEFAK5OX6ew7ZBzlae1dqIY0EnfwzaeNug9Okl6ZyvKlnK1kciNGJh/A4
FVYikFSNj+PmG6ejokxaEOymmcj0PZFWL5UwH15lhcK2GTKKWKHinbWMSQDM63pw
5ScNXFNVZKQDXLrcX8m5J3vq1mTOTX/8MtXqiHjy0tzwK1K/pjZ3iObku4vNdbqz
/dFgy4MGyhH54Y77A15ru8mH9BtRBAamzMX/h81uuqVpAZr+nf8rGQ8nwojUBxh8
7+jO4vsFzQnG1Wa/RgOc567YCNlsa3gLbQm0pIZTmPfh/i78GCvE8bgwFa2xrXt2
QPj/MGdriUOlvXDW5zx1Xs51hAjxCOoIKdB4mWeRQUM7BIfBjqU4Zk+Yjvr6bT6S
LzonzA4zRaHbOAj/dqdnzAPKngpWPdsvWsSPNlziXE8WSf8YJsZIvw+4QBbAP0UJ
4DZjYOvXDRjwVwDI5eC+WpmOZBwzv97BpOpX5NwjMYoYjVDLf7shh4Dkr/k8g6B7
7tJrp18aj4IADWyAZltvMTZF6MuFQKgDYgsVvGGIXbNJqCB04dKbR534SIYApva6
wymW+7482zORd9/EEOdyuHv+8XZPetC+F1HflgCR8ii7ScmVCgO2/a3gWBnz59ZA
NbPYPJYpn4K0HmwTtjFLZlCCFnNo7mXxxImtC2M6cEb6nN244iF2HvsH2K6gVzeM
xc7lYFSBxV6ldyrYd9lJS3pPMcPI0L2hSuhLePuro58n5Z27aQc6IeJJue5i1tEu
gy7YQARiZaUvyUndsHcQjxO7VVysyPHd5V5yPx9AHC9N3uXuwn51gv5V1dfj5FwL
sKtGdtfyghhlJB21VH06RXrHE7D8NThTq63ADb34mq6FsdVwi2lTjSntj0yhZhT7
Poa/nLVm2Rvrpv0w823Psb5HOW/uIlOLtv/UKjNzG2M79L7i6IoFJgiyTADnfVwN
rOrhrPLyBgxQPAjANmq65nb/nBvWsRVPH3/6EeLhWAEkEYbHCMw9P6G+tOzxAiG/
n9Jx4jTFTmmOJdFKKsKUt1VBH1ltJv44Ncov+LAsBFXLe5Wk9XL9BqcdOHtaUVc9
07jfmmHoOlh11B8oA8FO3LikvLSc3rkMIXr+PqNfq+2fNBud6eCt+1uLLRwBXYe/
t6cJ9IeZnBRGNhxxbxq9LazNEkFxD71t+a7svLy4JjGshUwpfqMoKGGhLF9Cc9B0
lTwTeb+77J2a8OJl9AwjHcTpyDFbo8K2feYu0KOR/Ki+sZpTt54Z4Sm5zxLEdphZ
Fq1FIUHJFhjTujnaPR1ZPMBhNdf6HiS5jak/T5EkRwafSrPH+LVmAfe9a5gBEE+U
ygH2PhLDV7Ni95NGd8fqCUtzzjxNQlStndX1LAQWEoX7dYIKafCd1c4iC/jTFL/L
GGoXfUMjbwWN67nhN40NdzZKzNQP70FMwqKPlk7mHUpPvFpgiTvFA9+pApPXVFsC
RxtJshnyBJt5Sc+2nmVztcm0KRROEklFN0rGilsOf9Bt4Q3F4ZJGRIfD4U2ACRgl
cTiUT1OmzveCr+jyOwLD3mlK2tHMHt1QFBf6ZOIcBa6gXZ+eTaOAFqzJWoDOsBk/
0mwIuN2SLappSozCpqQPRwQAsXakdbtfMrdeH/BZ6uHb2EoiEuO6vlL4DevsUM4W
Xp4yE5bHGN8tadQhnPoxigaaHCT2vfyk0dbSKBgYu5RzWVgWEvWrCNhc3qlRDoCU
DzeUFPPjg9FTZwdqGyUzw9xHhCidLqmZ45E6hO8Tf67ncgKOm5M1l2Ijk9ASrO3b
EQZiw01d6I26ArTCG29kWWIni9ICxmtssG9iYReTyOgLavXMPH5apoyeFsaCvawm
/+tKo13FTu1xHqMmOjCoC52gH303tqSznrRONK+FLOgQqAGtbOgLNkN0BXufW5uA
Iok2c+Huw2sG3JKUIxVXMCTckAWMZgW6Vf5rpNWUVSEAk1bbXJjMtgyAVHjxVWW9
VsA+EmOeUP4Z8gZtnemhIf7OAgs4RMvo8cHuGn70gpHHbQweXHObJOYbMHCSjH44
nkw07gZyndIK/zu2NuMI64XJ17pu07eBytusi41D9pGJL8UXoxg+M2VtyVhsVuxp
4lFXvT2lcNkBscUN8EHsPIPs1JYGXnGYmz05+4Htqo2MY7j/ElJJ6c2OZVncyFeY
XoDE8zN964TSkOo1si3P8C4XcULxgMH28HJJICZ4GNibWrp9TxlzeHgURKVh1fGM
4labvXbiB7jUacNSxTi/ekKBvmo1PdbtbBX0lJLMQLqoxdHKz+tevpoBbLB1psHE
hm/ggGMdfyJoH1AzYhZFyAn14W842GdW3FJ//iJ0TpGavTpkpDXs/m2mNGBUxjmZ
hmrtp2n+qrCsrTT5XC2u9iZTRqG47c0a5JlMJjZrnW2hDaA57zEjNafFBB7MY7BK
iqKwL3ovuf00PReUuLX4j2R4mnh5IrhPPGpIXI6IuJD34//AD9WpipyWvq5o+Y/Q
XDESiANgKLnOSm/JlJM3IUr649fq9wHhe9hdeBZFKU2b+HYm0R0Nz5wVXVDOUL6s
X9X2bwrcBKqfb4IIcE3wVfRNGANqTVjvQnePvbIYFgh2azGyyxCFK3x65UEuRaIX
8JnT8Q4lNFF+EO3irbzaz/Pt2ZsJawQ/j9j382vSqlPpEOZ7KrsZNzwyHReBWANw
G5WEeMTz4lZ23fz6s7EHYkUgQoxkuhyc5I6sQ0lcwQpjtHMHP8XZpdkRveubfLDl
t7UTUdaFc4IbOYZPCv8D6xQO9/n5uIn9/WSwUwo5AvBVFIMCmi1/pA6nZxFCSOzo
oUP/GWiEGmWFEdzE7Wd/tDXgIZnAYo5VqcI99OhhVuG7wx2TJ0wQuWszoSZC8t16
l9KDVu0mNuqPPRluDcqqoo/lMVDVfSJ0b+yHntv8zBLX2VyPdcMTtt1J9vUhZqvI
fJMmG8vbKq/ewjNsZOFcM92bLdKa9Q/QYGzwI/rVJq3tMEtONduxrLg0HgfThCr6
LqwbSDmzVbA2lM3qiIntk6fpyJaGp3NFcXzu17fthIUKZJO+8cue0NGHCBFX/0BJ
POY6lkHMlv5KPlFX3vqWyziOafUOliG5LsoBRaYB7UvainN/gOt33z8cDk2cKF+3
nHQCq8wWutkojfm/aK9sOO2e+MOz6B1FV3lH7bpLUb1ukwCoP3kn8zt8EXxko26L
qUoM8hSOjb8b60ibvxnJaKpLy+xVGOQ+St9YcgMhdhSgHgi6VyMV+LNLx0CkILPz
ijmIBOM/9/5K4GepU0YFtn2SlX0KzEpOdLMksLZjDFye6RJUA0B8qWFaVr6f7h9i
F7gZ5jthfWJowGeWBrH3x1BB/sV18ki2Ni+HNTkccM1UiQsloGwhwKsSiYmWrTwv
gz7VjVGlm12dQK9vsoWUeq74fL7/MOpV6aqKRKXxs6JiiekA2C+1Ijn2+N/qFpSe
nH98rz9vElTnqlFAIvAXHSW6UbThI64rrXHd7Ulh6Z2HYIxh64+3ctne7Pk3/WqZ
W+gLRiQCaFFuwlNrnJJq9Ha83tlyIRE/0TTtsGrSK1gQrPvKHsk873+0tmndsskX
+E1cxVz73sm6x6CJV7m4YZCUQX6WWmZnaB4mkjb5L0RS2if2JE8NhM+y8r/KlStk
OqAryhdoGaneJjPUYPgG5VQFLqUvVemj8brYEUNkfDLdvFh5N29UEMqtMLD4T/rI
BmIQPus7W4bwk2YJG8Bn0XD/LJiRlbLqmNK8Mm8kQBOTWKsQ0QR6Wm8uulrmdmHA
qNmyKS5IUcde9bV37EuSqnCe280+A2jiF5ztJJntPNDvxApOq88ezuERo3CzweDR
PrqHZQI5rqtea0q8r4zwbV97NDmbKBhpwzbmB+Yv+N7t8Q/92T1jOz9E7/m4lLLI
Y5QLltcbjrKJUq3I8M2wMW/gGPXmQAk9vWlD1/9HAAp+vr1vS/pgNV6ATnP7XRw6
ZDT1OQXHPjTCwUG0prvAUNPc24OIbuASoJ73sGAffXDTdzvLn36EpQYucGXh5Q8M
JtR5aCK6EQANrsXUhuhH1vTaXonFwmFi8b99D20b78W1LCpEbBQcbKl4XShRv2QO
0bp4EqTXu8sHGT/bxRcD0vofPBLSjD/Pw0JA+OjEvVuds4UvDJSBvaE/AANjS9cz
BhhyYjAhqg42vrIRbi1FXbdbuC5kI0avRSwUXKNLcdKn4F2mkwEMbqB38Rw9yi+X
fFhnTq4262pVZbW8VO7Puv3F3DaVTbUdUa/rMMhv3KjnYuX8OwDyzRSDaM5ORWKn
kgqDLHXyuwzkQusbLB2u2p7AoLB6mgYaJ8DAJC4w+Sz9ZmqQCs2hIQ51KRsOUzPc
Lt2pH6RKAEn4PwzcIepOn1nYFhv964C3T3RjP0GGimczmACCsX3+FPnaWHp4yXWB
K52KWxgmyDFfsSJ4tx5ZXzGuqmGNWByrkuEgyJ99mKlIFs3dtn7wT47Z0J3g/FXS
ol6ok67J0zR0o0VMa1mOp2zJnPjS0BOzHL39ClnUAFthv6SBEnzGOpzVuS0A1hNL
AC3Aj2woKn/V9nX8FugUU97c9AlQ1+aEYNgczhv6hBYZgbvaUoS0aHRgQhjvlM7/
GZiJmmnvfFggiBrYckx9pc2UPuMhs/mb1wE9vTymOBracngMBxwSYCXIneCcdKVd
Oj9D/PRdxoPutLLyYoYEU6HKZw+GcN673QtVmH4J6NXQG+/SthMJzpmWMcZxdiSZ
EkQ2ZAv+H/ernX6RaKBuYPaDDMtcOH8D/5rjstG/nxP2O+Po6V4RO0xmqC4Ogmbq
q/dX1XTHSIfTsxvOOY6hOFBw3lyYr6hmQGPBrRpI6LZTJLOfez2FN/YUtHHtCKiK
WbdSBCLmj9OoGf2OaPHX7L3hmzMx7EPtfQOOG3De01v5qaGpBJiZfgaBBOR7Pp78
NZE8brWaBVtDjkLum6TNNzjcmLvw4Yo0GEaf5ThXsWjatLFxiNAKDIqiGFrFoOq/
v5BZiCdZj3HNSrTO6avhWv/WMfLjbEiepeVfp5D1ChMJlNOGRSb7BlKKdbDxHu/3
vTfftdHAVpFyAix4cz5beGlJv/XJXuTrUOvoasOZOcKU6Sq4XdtxuBx5fIaU0ntS
UQJdXBSDt7kHW1te9MaqK1YB1KCPskiuvqzt+MW2DF0j1qa+C/uhyJCV8IuqgqGr
zWuTr7TEuMQVyzl5/64zjrP10l6Sf7PdzkzDbAtICClaRtKAbL+JCboBS/xcfZqR
K1kTYAdj3mSXzHufytc1M6yJ72Kgxr63nTkanbD0PuZi3BQNA/egIvtn35OTWn9q
hYa7IRpKmRn2c0u9/qmTYvHQbYd2xCrYMU3HoU/zgbFabzCG2S18XQwJ07G3DSC1
Wt2T6w2Bl3bsInuGSmHrBWQqmYMvSIJyZPhihMx7dF6SYSQrsZeIQT4KYbAjnsyF
BvQWdAS5NvY/PtiaBqrFtTpC70yMSa37A83VyCRBzxLEt+jUzAp5JfPGBrHqFnGn
zLrNIyWNi90TQMMUrehinDklN1FqZy+tSdR8CBBKOvaAffUtxjpQE/9WbpjuczEp
N4bgDQ8iR9MhlT+EYQrop/YXXhAkid+GoU5nZl3QGBQACr+Oq+Vg+h5jD3HsGrcQ
mL8G9hz+A0F4l0ivNk6/y+fnc5Kjth6PYqgklLnq9gqjELhFsBuYHQSHUgNTShbp
JcdH6TDtui5RtB1aLdsj6s/v8TWhxJjaVvO9gHWu8I4S2Brmx0f772nWjzAr31PW
O1Y60rGu1Zced8SH33FtfR7q69oTi/HDrjc3VKi8kFAWo8cPtp17DPcdrjj8ULpJ
SzG/dlXs3h4Hvq7BCXLeFqX8OrN4H8qck9qGyV/RRS+m5h1wmyvdZta1IeTWyKGG
JCEaLd6jzLgxvWfBLQ14dstdmo80RyzceCmNZkv2u5J3UtKkwevFfqtw3b4kZ//Q
PkMEsRIqUsDQYUKK3mlaOEXvA0fotoKTP5ArSP8RiWyvn1Lu2xGInfokJo3vlaI4
Kcnlg3DdQ4gsBtkw56yngONSfJ2Dd/VS3Y1AWg7ns/FPQwrNpkzK0i04KP/wM6P4
oucu49669CodPB/r4+EwQS+/tQhMfw0Ba+1He9khyCWO3mt9kWvPzKtTUrxfF6by
naLSb+rzV4dOMBc/IpkQYUoXxEcc78tLSWW06+sW6rzdE1A1c7iIDl0yWgJRQPmW
3zCnL6PvuCkbf2E3gb7Q7Rc/VUM6st7qf1GhSjzRTcYmXWWyn4FCTuxlOTTZQVdx
XEoQxuibPJBLV6g3SEJ76I7Xvsr873f3JvY7XjkE+RGuqvlANAej4Md2ylcVaSmQ
H0z9bJFkfFuXdu3/+6ZRc8vHjf/HhrNiNEB9LLnQHSiDbTGD8bp3cNyvAsJat5JF
X9SurCMsfRvTDwOCfH+sMCj2rIrUN+DSL7AgYY+ucGTa/7SIpYtxntd5HZ+zV53w
kGlX+egSS2Dqa3CCDAyCvhkOl6O74lbfKO/bukN9BPHZEavpIvVETJUCL+JdfQcM
u0g9VwEihNBBAjQUkrmYsbXMXZ6h0/pidYAvUhyqxh4KpOE8SUPKx4VxmX+Ck4N1
JghMUOUtYWpTNZrrBPQB7WGiT91/IQFrJEc80q++vrHnCsKaAQKJvjzWR3v/FdS7
LE1mcjsAHoy8HpRjBSdby7sjrNLy2u+klqUlJD33un+XEMgxHN0I+54fw4y+EoY4
kR5HkZvbSG3QkkxHfxcavkiEflNYJpZv3J+hZq12vdqdD5cNqCvaoZMOs0hVhBfO
J9z7dRBlo+WGblUTwmmk5vYH9NUh0RA+YhIcGmigmlMDacMdJEySxXclmTWL48IH
he9wdnbN5hxTxsvVrpjx7+EjjenxG6qmi5nQPP72aaZ+8XrUVK8KdVU9AthbIbiH
3T7oMuBr2o0QYfGbtqOTBTRFMzxWbQVE+wcLuLhwJPkiT1bQTAr1rg4DB6py0c7C
5GSEcDctkbyzqhbAHFzxQ1eRGPrwCyUMu+e9lUx+LfodaAYnfub6wZZcpXgE3ZJB
k1Tl1V57DGz0Na8UGiksHHk93Tm9SbuPge7xgwoQhemFSf9QrgDUWfQXrpJ7BeDZ
vEh1d36hu0Vy5Jfzie8InU++1NMYiQx2beUr4OwmvEFsHk0pRzhjOjD2onVXoRh2
V1Oe4A/xbRLNeJeV+0KncydcUGOyC9TJfCVOlspMdyd1U1ZWUTlcc36rRZk2CDXp
F4bapkPVevQ3CPIyyYLONwZfHekIBMDSKwIzBDGNUvH45W8OpaTQVMH3unkG78kW
aF0V2F/v+8gOWls/7RvhqvW6x9H2zAiyrYo8FCUhDO044gRDnQvBVihWR0Anv4ni
lZ6iIC6B6/T5Gt0Emx4vuWCgNYy/rFv6us2kY4OjuvtW37aXU89MDrLG1RnheDT+
VksN12Eq9CE8wn1hGgWKvhuBLwRFs9kP3NrQxLyEJ0EOi+D7otyQLihYi62Fo6Kz
LYg5U/3OMOndvNOG7VWjfz8h1L+Je203fWxSH5ve/JnxSwTh8mZ0OzF3T85G7O32
X41yqW9nlxuhlz0Cgev3Cav74g9IvVKBna0nnGy58cfIqJc992IS93Fs8dKqq8f2
i7Xc4ASKAHxBW54L5XowbxgJbxHL6kRJzK4Qa6fABV2wqtGPndJgwjN9EBLeBOG5
/gGvdaKxZwN7lYsQ+5wLGTiqXrJlEg2zDQtEShCOjsWJ0Aoc2Ft+WRtnGBNY7W5P
JWPgq2Bid+d8U1XMeYh6/Fwt7dGm/z0qcM5flPKtaxKH/5w8msHSWlcT/EcXNPcb
79qBdQaGFcuNOhEV/hB3oCpZIyDkiYXMcRJTbL4ocwQDWeVUJes7Bc+94ntoX5+m
gDuvaCp86fWMSy8z1XvsJJ1x7SDawd/iEE7iyufHIfekDdwgRMkkCAJoU1JTa59p
o2u1ziipaK33ZYIsp4E6DZxOgdx2/2dvAopLX+Pj1xenNXtg/bIXrW6lGX9p92iY
sQUe1jqFVL3TX5tRlUr/B9scnjkU++R3EL0hXX42Cykt1DAl1eJFTQLxemXt4Pl3
Iv5eoifXIl0W3u/tAbToUvfoXKTrqwtKiv4JRy7X3eiXSjKorpljlbsvODummffh
iGDAPOmfh5mgwcHrwAsCHxkH0PnanOT5WHYOJ2pDzB4Hn2c5sTKpb383PZ9nM8QX
P39KTqhL5Rhro6unJ4rZ14Ktu5WImCETPUXLGtxWJ9yuCLJdhpexBcuHXD3t5Z7Y
FZyHCcl8TI+eu4Jg6GP1mYGJk7yHQQZw12q+XNuTYWw+K4QvVmAUOYppy/hvryTe
AzQ5YIkL1Up8E/ItJqlFekn1Cbg9HiphGHOV4m+NEWBZ8Meuf+UvN4FkzpQ93hBE
OEUp87q7lsbe8Wc+8gSXtqUV5ICspGyCrBusa019z1kaWWPf5FlNsFLuapcEGiu+
Ypjm3LwH6g80UYUTWrfMTMX/hEeF4x82Y7rgS48cNRSlE1BXSGQledoDbI0ZFIRZ
AiBPvatKhNCOCfKUC4j7SMBpT+gRIbWpsTmBr2y3gceYxvyC5pHjKLaJ9xFWqbai
99puT5j2gt4eDbmtR1icUyXmlLINke+vQxOvzs0B541F8p0do0QG3ytYOyKv0b68
jUYOm4h4LiubLrk5yb5KcD2cGoLwd39fjhg9m9j4gPFehDLQgisA08eZ1HJMWZzL
URNLm4ncUOENJvkQN5DNBnvrLPT7Myt4V4s1VmU4H6yEpuCBpL+LFqaKWnMIsntP
PdZfoHaNIV15EejNyVdObLI6kJ0x51dBXZj9hWN9Fbrb9MK1pZ/LZXLriFweFO/u
mXMjcK9OhQDVALp/kt3nD/1QVYDGqfbK+nGiUWaUa8hdvL766PM6BvYk+mA6hUiJ
KZgqnq6P3/q4tm7Z/lX8nQMl1ksIR3jJUs61gxJ0AT0b2ux/hDha5eSh0/rpmpnM
oiuFJV9pwxhIjbGoVECXCiypp71pCsjFgJTJaTslCWP+tmmzKYbSzFkD5hiUYRI1
X6IOLV+2ke6JXPGPHP0lPo2p+L+HVFcH5FX9pqAriv7iVHZLlL2fcgE/dhNDbc34
siLbMpmXxVmt94k19J2RbbuK0Bu7G3n7rpT2sJJzsEBvbRe1lj0sqm4XKVeehSPt
mDedbIyoUo6f/WUFsRpdE7GhuYIey4uO3UXFEyGopk2jGQrCVNHvA/emZ6eiL+s8
xImGtXyMJMjkoST5Qmt4WttxaDc0OOthsa2RukeqLVuyVI1GdcfXZXB9GZmrP04p
ld5Y7tXWMcy44M93qiirVN8SLT0ZCJGP+84iyaPAmTrvdVkKMZyhqCIdZ5c/c2o+
ygxwygkWOhAzhlFBWEW8I/R6T2zLG4cYVBqGT42H72n+mjEKxyM4ops6PeY7HSz6
0Amo4KKphcObVeXL7cUxvZFzl3QzA6YeoEvrFCCLbR3gNx2zLxkCsZ45+lwu/i+U
ytW2iJT6Fo540du5KMDhiX/qJB/P2Pomvmr4M6wS2xNv6Ef0+yf1a70hO1F5QAhg
bKcFOXIH4T7FnRz+/gwWewwLMXC3M5uXcpuytp3Cyq41gSNEjRt20scqhQJudEsD
I/opn5TsKNmYbNJ8ygpwgo9F7Y0L1OpLwsej0Ph3uqzCzfja0+DzmfghMbeGQcR6
04klL77YCTynL9EEwYaVw898enVI6qSUtKrN3T9w52+SVlpafJbX+80zdkrU5bgD
T0r99xcgOeKSyhC579HeDyDBKGB4uzgFTnDDHw3AtKS0u2NPrvREnKcANoeY9Yzq
c/O+/4jf1AmmugnJjPHYql3R36DsDT62rRvB1Bg2qcXHJ9QTm9+iHXAAR9CouCy4
7ij2ecVmw2VZ4CZFfoOhpvgUiTzNQg0xrQVaOndFPrpA+ifZsbJ52jGskVjW+sdy
C0ZnbgO7OZDqK1WONTFsYqfJFuj88GsdyFW/53K/QeVuxPvLIFpW5oL7n/f0ITQO
PshIILCaBs12q6UY2n/6zc5XCVgCxUzmGi1Km0tSRsKtdEVCB3Lbqk1AuTSXrv3B
3Iwj6dhcDaj+vNLcB8KeK037j783ziUkB/mOs6KSv6Oki20M4c5ZNq91ojXjVTTt
aM/jU9krmP59BhoDmF1Eo8f8NKS5dwhe4H5kKJDYtUeHFnUE7j/MVWKfuZbfQJHE
yG2W9UlhN8G++6yW5reXoIMktL+5AWaBdne+Otuszap9M/PxVGegxqkO/CNqJgYO
dePEH04JDzERWEl2PbSmwhne1jOA+jldy9vjAlBZ+Rr4bnARllBlanqlxUx8Tw0t
ljCjf4M6dQIXnKACAszuKQjFT6h2tQdrWldv8ykA089spqWUVcosiFRP/hbdcb/1
foszjwBi/Zp4PnWYFSovPgT8O1p3mv/xVHZ/G3HhMWxz9Mf3Luppyh9ZNMtk4qyH
yqUEm5xmuYOBWUNL8p1BZxTDATr26/YKLXAQM9baDCH2ysAE199sb+ToPLca6MkL
/tV2qC8RX34rogEgS1R+SKEZ2jAheUyVcHoxZwN5xiuHC+11iX/JNt+wJGjIcJUB
0aulb5++ke7+ReAC07NU6DMm4f7LCK8oVI5CA/PAKO1gkSgoB933MqE0JUIf8+Zt
5UPGbsJgdXIXlSVmvGsM8smuPQ5zHxdSrVPdLggCA5JvZC1+KkQgvzc+e0p9OswU
8X8d758anlx6bH9XCRCOI46bHHKJPxFOiocTlmQ9NaF2VOcatngqNaQNkjX+WjUy
CklMtKlaMCPfB7faqJvzicI5sBU6HbV19ZLZ8GoOpD6kY1RsEVxWsTumd1GR2UYf
GLncXIMfSlZ4oisoIJ/898ZNbxSKbyQ7RmVwA+ec0OgzEX+kRCBCCbY36ztXxwhL
zEXibZrO8rhgyhAg2ZHDa+k2l0LMCdztxp8j2NLk/IoXpr13DICuCjIo2UmQHhii
dg0M80K0VzPEL2oeUkiXH/lO20k+wNE/wOCzJXCggzFqDe9Rt8v7Y66OF+Fjde7F
JNE7QAkQf5sDfo0GAWJYL/uDzDxQ5DGohER28+wigAz3hFOGiYAIdZaNYhWN6Uou
j26VdBhr4JbMb0WUvKh2yIX2A+V2kC8nJwcC6YB+9ktfSd6gd+++xSDNVyI2HMtX
k6opD/UmvjbcVtok6IqM1jNf6J1FcsgIP5hIFf6T8xaq255Fb5J0vvA1eLb57gq8
JNixwx3y5vKLnbebfSRz46FVIk8gutnPsy4o4rL4jcAuArp9EmapEBJiWbTZMugz
WTTiyg0hFtkrI1B8YNbY+Msc9pmRsQXbLvEokvTGDMgjydshD7mYDBcE/oyk3bNC
92GBdIuPzCuQc4TmZhnCXVHmVUuRpNeFc9ylPyazXOji9Gm5YDNT22i4Dg2dBRsM
gvhDvbKgiGqjeqmn1zMZDpI9DecXw0eIJNVzIFGLVHe/dUsuKLTi8tb18oQtlrv+
4P1Z/NhRITwZVhntPtCQKuiwr6xrhpS3WY9C/8fqLa8vZ/uv1tT/RtUo2HIz4eCr
oZ1e12jd7YVi84RmNAlydR1H4rR6zoU4mzxOFAf4nnMUGLCGr3xQd4swLRwbsrbS
YUm855Qq7gLxWdHbGDn3lDxB93fckxn8CV+EcYVvgZsR6jkPUVFG6EjirFZSI0U4
zRsBOSR7KA6rPsYYSfm+ect2U8mxocZqx79Vtm0LWHmx/kklLDTPKHJchqmnfuvf
uiDNBvfQpnAp957O77GFUcem4F+p+KIc+lwBwAot10HwlFTU6i+4T6AcIDmCLX59
CBtqZT480dz1wilSwuiCUA/qILUg+FY0rn9jON2qUlUl7rPWW/v7FFEPKx/o1uXL
WJYKTvjSZ0FDgQ6yYume91ihSOtMYAMlNEdorhyovK8LiqkJpmovyHaq61BcPrpg
EmGMp1iGItvkBGGUFeT6b7ClB1xNHC3U7Yf45dN+tUszAErOFKwdpORrkGszdV1U
3/i5dD4FVWH9dHR4CEWy1EE7kx0/gG8xFZE268UkKUa0lIzt6fTvDd9ZfWJmppCV
WHI5pSBu/D9cXmVScTQtveP4K7A5nhezq0Lm7ph+pMMSYTLfQPKY5uUVlm7Ou7XW
28wuTzVSO12+ggcDVA5heBqENv9qYW0cb5IgzH4ENxeVm/uACnKeafmus/Kblc3l
erbRQv28TQDPX+hhUSelnwMYtadZXA9lW4l2aRtiYiGf3eGfXUbq2ot/ScpqZzrS
IqomOCiSJWlN9GeKKv5iO2M+aaS2YsgL12oaHOxDOzpJFjw0XtfgmOBBWpfXgKqA
m0EkE14UgmrrYPL6sEy+5HaQ47FQSDrOpkrIU9vMm2XDVWQxJdOgEmXANP+6Zrv+
zn5QUQ9mJ/Y6+oGbw8cF9IAKmYgTLHQGv1lWFcrJyi5pkuZqqZ9srcWaibejPYdT
KOtH0nXriWuCGQzmJSfwYUl6rfeHTx/HPytGzwGm1AktspxZ5ZSfzRFHNH5Xhrq6
xe8PcmU+6FI3qSfybIgUGpuSO8d28z/UgSkw/e0NOaibJDvk1cmajvtTurulZjCy
gqhkPm9QrMn0RbI3Xscd2HLCPU6E8GNweJr4aLcKEQsh8KfGRkR9o2CzotDg6wVS
jqWNSDD5N6G/LYXRgCz7Abf/aDvxOzQpCHyEgnENfISJ03A7WrTGOFbHR7GlaFQK
0rPip0jgQejyN1gla/1kFjAi8spCq7kmzu7FiMGVrgeeGmLkKAIU1o+sfYOgD3VL
IJgbum5W+o5zXwUSgi7GLH5bt4ZMYC0Uz5ifKrd3bI7IqVqhSDwwzXfG1cSQh06U
PRQ5wtaKlwu2wEHDX0oBl+swDyPKSG/FyXahYpN22NzvO/umtkivThamTAJrCgUF
xkluBUgS8FZ/OYTFOZvqstgpLsMqmx/57NDwsWb56MNOIK+AXIXz9mbxEdiwI9ir
eZgvSV8BMydsG3v/i2L1MO/61djWpMbEylG6XlBXjwRx60IxOJ97NNwr/JEJZUqR
AgWQ9pFRX9VlYK6dP39LX33F+tnYipY8udmB159GSbsVd7KDkq/sQYBjSgSgR12C
44UdJnprEpbZeIIl7qJexiRiifIlpxX6tf5xEtO7B737Mr7l/bnt/UA2BKRnPM/d
aqYniu0eOakI1IwLHNWQ3XDFhPtojkBtmDvooFr05VldPV2eQWudcikxzyukO80q
MGVkWxQPPtYFLIyCgETLtrlBx9aDGYiA9kBgxR1n1MKU5ek1sEk9bvBM6HYaA/1k
n2D20bWQBb7Faxcz9S3h6G5hFxnDP+Mjo+kGQViFR1HIbcD1pou0w4j7IL6FQgqO
e4syrqJhpFhr/k9ze3R+8CfaebdfOYWvNvQwq39zVyPqsRRDfMnO29ygLNbfqJmU
yh4tEe8unsmu4JMuyEU/FhiWe0eXJbpMgDzoZJ19W/koNBqSz0unyg1yxnfNDRy2
OHPd8LvKckJRF/EFK+mkyojLhfkCgSRhtPteMKnAxYfF0gpoCrGezvpN2TCHDsym
KTYBQlcMI2Av9Q0Dx8Sf+vpgvRBhOsVwPOeVWiS7nfEnOsf4M+nLgqfFv7yR+z4m
cpP2aA16lx45HsD6Qqsv+lfj0WbuTO6So8hzzzR+YZ63PzgPoX7L8Xp866OdOEGi
axjKjupsgXJmWbeTtoiAiv2TIQjBpT6bPO0WD32/K7+OgqCMASkHU/azBJlbFWQO
1/53RmJgSf8ejdbdOuRCMutGW1R6bEqFGuGgvHvMKvX0DFb5EEx9WIa1r2Tp7O9f
r/DZ94iR6qilUUdLUqKvx2KfgO7Ob+gTaliR6djNsH4oDJ71bUQlqNPbMPulz2fL
vqTZf1hq+fvX72KRH7JREq7ZVbraC1oDO8lAeoZab5zMbsXVuqfOLw9Q6R4fDrUW
TjjHi5b7LnFgAqvZGrb3dFmuUSFWOWHTzIU7eJRfWpOqycHO57qaxHkmQ0jhDgwm
HUClcrjIYJ/wshHe14tCSToXUesXfnjohSFuxtLHSyzlVPD35K4GA2PUyoppkCTe
6P3M5HGoBedfigHCbhfl21ZQfz+5AMbiELv64g9nmhxRFZs5SiAyjClQtdiJziSu
ssokELb20AbSfxDUOcEbKqJYK7MN9LiCdTzkzwGORRUTlntFZslekPVgqPYmZN6d
Htzrx01JYcEB+q37vWNhNOuHgBvCNtEAo44sOwr68UYEica+2o6vmVytisKGYhQJ
oitYOqmQwgfyZMCCr+sXZJUHN8Ns6Z6kiMiSiW5jAqA0oLvTELhkHGN1Ohb0/s04
BSX5fCpyOkW0QFHVma0wQ6x+nEwJ7FcWTOvZOKDL+bbyg64bI9rPdtEfxMHayUCM
vt7uuKR3vw20DyBZOePoMZCpBSC2B/4yNgkQZvXI4Aoy+hJBI68abdzAXy5BrZDt
4ww/IbXYJR53ivnZD5rgO86GmHdeECd5oFOLd3t94SoV7cCFuVXr8GXj7Wx7Y3V4
6plSZ/ohxF9Lr+W1I/IDb32vgLHQaosw8HUjH/2L/48nYRJXZhPHotYfVtSmfI0n
5rFBinCZ/QFSyPm6Jz0xEAHl1C1nxcXllAzwrjYlcKQQPsuG7l2rXQe/Ff3U71xK
7opw/ga4wzFy0Tot2p/fWhFLWNEhOXiWkM+jQ/GFM1MmhhOxITdYz85Mk5z8kr3G
22GJksHcsUUzfOG0nEbUroBeIOgUJ7RB94ce8M+UekAlU7lubY8K5tQ3GsZ2qinR
IpAnk4xk9ceOcIfUg3L16rYjGfd5kW2/mrgjy3k/k/BFEtZs6tlIPX+mgAdbq6ye
cHNuXHTPVv9/ppSM76deyIz0E96M25V4UYibSAaynB1k98Tkr0ivTJefhOb5f8aU
bgDS3Tu/FemNvM/lwn0l+9G8kHtN/YeXbxMdi+NZGrEW+t57x+brR3UsXulDxpJy
yU1G6zFSga6gbnrOP7KqiiUwvY6xRoAaqabvfBhuSWSjgZ0k2fK9nPeOQ1jXco2X
1BLtOyoxt7zJeoLEP3zu8+FZJ0ls1bS41u0OlRebqqzCahnDzJ4UjaZZN92S8ruQ
44UsIsgXOkR0x9R5QeZTq5QMG3wx1Iedjkz/YOzQkmgXXJoHlgek9Ujt1i3l8RnF
ZULxYkaLKK0YPfgP5mw4+gYJC+zDevs8f3/MIthaLB1JVvtnm049jWu+x1UtqrHl
NYmTQ4rIpX/LFI3LaCl/hTcSppufJDPVUs6OIZMZIzkWN6fgzw6GjzMsInnsp0AH
NaDPRpPfTxXzD5GDpknkXBVclQX60kwI5GlkkSx6l0dnqeqPQQ49z0G2QJObkyTR
wVSFXl1qxEbSjyC+5CNxoopuLnCWNnM7BsRKYnriwbEVwPln3iw7RULkmBF8DTLr
i5XLtNdeoRJIknY0bvERQ96kBjqEKq3SsnyjXZF+KjeJ8Ww3qTGMjFJ6cEwQZldX
vXgCz7fqdQCPPjrWLV25cTdSbG7wc1qiuvPaxWyJl6sZJGDoRfM7KGLJXb8dcsnJ
Cja1Q8Xfbq4K3ZOtg+NigOjLOvv0sVBIN92U318B/O2OI/PZqrw5oXZtJ6FPV1md
Ixd8+sR5gZEpWdnrFlWakSLHuSBcbcvqh+bEPRrawbwrPVbWHMf+x0HV+k0DWWbB
8wloCLnIlNZO8vkDH8PzMFiFZAIRWAWrDfjj8na8HTupGlm9WglLJ4MBDDJyadNk
hlkVjso0nsvTTOqaCmJnL0yTN3uOXAIjgU8+1BYTFegfF8HDeTrUrFIcp36UKkbA
kGGE49WtxzWUyivqcYbdqypZGnSe732zpMg1k69KRXBOgrg5z99aNa2Z0EPQ0KS4
g9pIVMNYKMO4lOcKVm9PeWK4C/hcPmZcS8SOst0UGrBQISFiRQbINlJFMH1wNhcH
Nlge66m1uBSTTiW5cPi+IT1esCStJTNrMP8szncgwvbxVZhcRfVcJNpP7HDOlLxx
0pnayK09kylt+ZM+bDpJFvXti0YmrZYPQKFO/rZIO0YCAAEocjMb0XjTkyqLLa9t
oL1QnnuwTo2Ow/+d/ti0LwnzNyrv8x/JdmNjVOLgClmaZS2WNksZA/Yu7AvUMVRb
KIjs0Vt7xyQnWrq5T7Hw+j5sjjfsmFH18QaKHeISEk2NcO3iiFeRdn0H5og1BBlU
bcZDmZbirpF/FG6rwy2SUa7RWSpR3llZGOhEjUGsBnSK9g3oA1nTwZFrdXMjYNYu
3BU+NZQjZZU7gfsr26rSvDL8ghyy9SDHZGT9WIHgaSDFzDpKG2iiOWTuVBpGFscY
3rBGKyqub2qRsG9LQPLFZhqGkbzZi7eo8l12VIVx9tYhCcfl+UbwcO90gxIN4yLk
vgaVUj+gwmoyJ5E1CTtgxvegr3JauHP6j2yYCXH5E5ojJQCdpGPn9z1vDP70hn2m
G4xLO5CsdLw+8EZ0fgt99M/OmHq0WwQwHpO2PBOFQKaLTF4o1o8nw9XLKL6wZhTL
eLL7eppXZGF59HOvdqLlLQmy/wBR6ACJCQvUwActZvbp1xGvMk5Xfq40HfnOYaY+
IbEvUklIOfykrGj67Z+0Ro4TGyq4aKmwe/CPq+WfEILhvtGnFXL2YbSqVnmhNqzy
ZBhbwuRR/KR+n7bP6bVhEtPJtyndm2qmxc1MLSYf/Qn+GceyOT59wlBotnSZAxk2
bj54ens04V2QLEram81nkm46guPMuwg+X4l3PeOMSVOU0VLCv/8Ye7/VMSSoDLQa
gKb8InOwCC+fAlQIxBWKtMYKk2yQ/7c0Z8nTg4WAzVGC+KPjCvj3OhH2FummJcrs
bR+Rhn4mAvtDXE3AlF+am7aWK7eFsh47OiXDA/wObn2mxueCKS71l7z1TvKKOxHx
pJ96JtMc/0+GieVTBujL0uWZ9rwBpQzomge0DJknWoTXKYKRf8v9gITbTb/KsPCA
orWwCuWUSNfz/8lpSkdARhYw6RcNIHsFt3JTL4B3PrzyQM6ZX/ZX46k4k1hjJwhV
atU/151PLN9v+2SWTLCXaayoj1Oci7eFvuSvtsDm/6HTo0c1krv8gvo1re+8G6Z1
LA+es40HqqXLOwUPMMRt3yCrAj1w4IHTj/anrbk+ohTFGdAd9qgBFWB4c0thlQZy
72vzkMBtioWJ/rE3aSk8qJ2lEtjQWgDGTDqJ25tkPYQaKve6i4Qnkhlzw7SIhOzs
m6k62lzrVi2cvIu1N/xqs8BTYyT6/ErS8GCackS2Qof3px+jYn0mxzbwQhLGbcPW
Nc/w58cuWWDWvmuD3WR04WBOi37JbvYUh+9QqwQBrXVr0jvb72YY3+vWCT597Sps
2pqLlF7vxjKKlQo7uUpHrDOtDwVjCSWDOGK8posvgcIk5BNDjmdAIOM2wVn/j24e
HJq3SWjEEiyx6I+QdlBpAfzFZ+6dfNDpYvE5xGhnJJwVDOokf7ISwi8/qWDAorRB
nNlfyghmixT/X+Egt0CkgrXm4uSMUXufUlGqDJ5kcFfS88s9gntC3zQHPZuy9jez
nzWXpjCTkb9NSk2p6GT+f2jywKWobfMg9bWegWuL+VXVyPaQs6uLfFrv1ryoGFEO
jwFOtdRb2KXnn8l1fsIF2JxscG2n77qM9FwX5MHOtsMJoI5iiDr1kwddr4wSfq85
xvDFGIfgXlPiio1Xq9NXheUz2thj4tCNN7+28lOHuXiytWKKlWqrlwkNamTEt1mc
zRoKvJkjnNntTe5UY+U4lSfjxx82Qcrthi0gEjTbDsoCk11QRi9vosGVyu01oQOa
Gx9EikQ0ajNyfFGpEaAt+pHWr4oS9UdgfR/IKIJ/3Cd8zb8+jy4QjGH+okSdFwPK
uBEHtRuHIuKCHufAX2HsTPrBg8xjO3Pd4VrrBErnj8I=
`pragma protect end_protected
