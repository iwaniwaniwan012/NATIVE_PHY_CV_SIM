`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PmvsCVBThzJEMXZ31t4XPuDFECM7gGclWKH9GV5aDkrc268HVKpe5HtrFy4K8ALx
FIOK/mJmGIwRtieQSjpws3119CNNnExGp/U0S4sIrJvQJBnhYONrbigCVteKU/th
YL02tylmHfSlvowegJnMIUu/D82NQPQCt1Cx4ea3/qY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30144)
Pw32DoloBPK8skf66cb6tSK2PkQPr7UAsoiUoz3PQxdbAbO7iAEsDrChnTfr/BWv
l0n1V0DTufWC2S4qg41hbVCTR3VdhudZ0J2UzyRsnJgI36VqF0qvWHRkOiNOOtUg
c4Q2LFH2HjVld9H7JZb+wBfGyzs/WL8S+HZtaDXNOPi/xZSvn0ZihscwLAtuaP00
A253ed2CQTAkGU27D3xNIXUpVJbwMQ4jwM7nQjN7oPuo/NeiQ72MSgH2R4hyMHOS
AZVMQ5V+SH/RF03gUIvsu7nlnEg6XgGxDvFJ/snlc0aHu8q7S7nPN/KJi6Oo9v/E
QxvcXRLNzAvuiOwrELteEYXcnCuRzmh36t18CYapkUaCvPDbo6h5kuzLudamLcr8
5+66hBNGdr1JF/33vMnCHfq1xWUY/UpfAXmGA0SrdqVVKMqVY4v78n63Xubv6dGv
UACisUIBI6SaRN7iGost+shSlxE1ZV6+nql4+JXp+JFZeHsIPazZZH0TedKm85Ff
qLm3HiupFeUcpKjViqyY3hOxo9kSv7NQtF+G29ctQEYjaH1xuukXfIsaQ5f9/4O2
DI3VwjnIuhv+W8ZqrkqXfiYw1P89LN7uTn21d70nQ7iEDbyffqN6bsh0zJShuaOk
NXSOFFAUOJ8iPMe19FOeOkm90n/7/5fads7q2KnQnmZmk9vnJ8xAfy6Y/HaL4wmW
vyuUChiaG5s2IiFVxLeAZfSTVguHQbmnFm3SGTk6RaOXvb9BjEdb0/Ifj8S3PJtO
DpibJp/SMWSK21yc30Xjj7fpcscEztahfG2zB488kluv4DIivcNx3Bt+m5RKE2K0
XkL7hFEmfB9Qrwdqw/Dbca9hmceTuxCioC63oGva35PTimmXtRQZirAwke7CaGmK
DoQhs7Qd8Xmx0PfTNvGt092ChzkTPVOgM+Yys0hUJqcZ0L82XmLg4P0osTYJOziR
QCSounhf4p59k9gvrGXvPy3f2RLm5rBiXUN/ZltLarfMkwWHVPXcBJrZDh+WHVgL
HLP6kRkP8yyRG+hXyRzrkCle+YI3rjTgMzNLRSEUgqL/gk5yJ7ES2PrhzqoM5Zs+
mosBgQ3qVY6mmM/fd9+6tCarf/WjUznfWQaycC2tnteWT6NJuIyemmN29sbry+qX
jA3AX2hkCwNP8eMYC8Vzb6u8rdkHGWNcQNDaBl7AaQdxhXwYsAOZfassxax9I8Vb
b7HtdUADlwUOjl6l/huWLX4A6E39Dt8OE5vMCIuaf947xpjiEqDNsPMEeYQJUYZ8
P9LwpfjMJfz6Pny3Z+VXOUxRSw6+6WxbC14qxUARqupS6oAecdPtBJMHIgEmytis
++XbO+5FQxh2kQ1JEJH2Nrvh1jsFndTm6W6qzQctRojiLD6wzBRGvUgZfuO57Ep1
jZkqITuwwZyL7HxrZO3brra+ViD7tXz+FOD3LeKhkF914PbJw6F9G1U9L2hHNOQI
Oa0q4dj1vsyDE0VvpHse49XdOeB9o7iirHd+y3EwKiWjt7Qgxf2EtVmm3KAsNmt+
DKHscErvBJL6q2zYLZ7Td7XHj53sy7jEdJu7Oh7VE9prr73//VCOgKrMnbVzNhru
azTAetW34bhuRxwheOvSIe6ncNfVQ0NhDaZdAu4vdjAH2koWa90W76myyKJ75h7r
uFhMw3hJ2Wy28DRZ7brc8OFvBvR6I2LcB7wvbo4ysDV5yA0/HM6osTBbKTqUKjAS
WU2GsTNQs3CVosEHpxcETja3sLIZHDedet4yLMzmoFMf3sknuZGWWdwkgmdveciw
EI3ecIFVQRkcQ9y+MI0FpUsTbu71fGZK5i2GJmMNgZ8kbyGBoHaiBmKf36uSLLgR
ZXp38C+ymONZkeSmUZ9OKr8k9xyiEbHldZ+yBYjGCjY+zxC147aTKBC2PVb52+sG
dPKn8XjDKtj0TNyKmFV7pmKfiEG/iKuIJIpC6Be3aIqxSjj8V38DDfFiLk76okNc
QILQA3jCkzq9zyht/je5JT1++hhfFTc4zq0aDAKtjoK404Zi+LbOqggYol1GJWr2
55wkpiEeck7lmuJZRaeA94ObRmHrlloTfs8pMjn/meVcYTt97zp78VkQRhuG8dRT
G3FPtComAbFt0Z+0aez+CjhARRbwlRkm49oa0MPdSqcGOlleld1gvUGJu/TfY9T5
6QKrY6Dw/U0f4Ra0CZ0Jp9n+yymdB/7WcGyY9fP88+sC67jpF7sj6WnM1LCXkZFe
guxtrMj+ZHR9S5lTMnmhRZJh0PKWeFznL0WA8jVk+e/sRaGvlDmhlIPJF3L0QI1z
0XcIW+RAZvujsKsHV6uSM1fjvZvbQ3q11EjU/R1CWP9nD0CCefflhVcg1O7/Iqs8
eGAFyTK74QlM0GVyTUby4tXVfnOAw5oj1POQJYdErs750XNfID1c7BlcIX01OwyM
XAfmSEIPXSqWRJ3UpveUy/bnjxZDzgiiVnuJkjyUC1kpg6nAIvUXa0t++XBz5wFl
5VMvWucfso2K5m+kxu2HUjutbFSiSlzArrxX6zoUEPw+b1rKl9pQNNYbwDkE7p1w
Ye3Jv2QpOQZbHedqLx8KdAm0cLHPEufwHPFJ7zVrX0/9GVeDwlxS63w0bky40dxd
RqHdg/N0KVynFVsgZxSC/JxBJD+Ha+Fvas1WJ1QoRZYGD7mDH0rwmffH7Tl3dhpe
woYRI5P7V9IRrOiEGsy60VOJ3GNUApBmfGmo7POp1V+ncf9Q06GKS6S8ZhS4GL8z
F+fjKFp9yhGsQ31DfdkNxaWiW8ILNLL+uE1LDB0n+Rb5/MnAwWHrFdvnEPnJoTzA
vhvsY4wV9N7Yj7+63DzdUV8hqA8Iq9I8rZSlXXQ/cr2VgUxThL5zwurTN7hQyL0Y
jUaXP70f2ghS7f2Oiza16Du86qPlVlAVVX+TlmpL2e1XhyuN6unPl6fTB0XLBpZY
xkQQ9YBhZG2WJmdHFSTJyTndIBGSNvGQJxeKZEmjbG8yH/A6iXv3olTgmj6y+xiq
PO90YXutE9Ax3+EgXs08bm7sq5cNhHsmbj04ESaSJuoc99NuEanlaRNn64iTXaU2
EODILOPLtm59kULd/ds9M1O9pPdlZRoph5xWMF+2B5s6xdMq66ceDb5cfIlOuxEa
f0/R+/2uREtf6zIon9p8HoIIqU44rf9fTEdshdhylTUNOjHF0pSAFc5TviKj9Ki6
NOF8IkiLSkVjmJTce1ZvW+SOHsCj+yUkSMX/ZiQX+OEEFiQF7jyZMANy/UDz0Via
POWnOLvOTHUBJHZRsItfsOH4hCImmfiI9MIxLWMhzUaF0EPXs6CQSDV0iMK/KlBY
p5MggWsauzQFTlUlQ+K70ieStAC0W82OjJtXkXnDw3/qiz5PqXOPMUGLafOZtJck
M4yL5bbjUeRhZyanqpltEqmYEpygYcYGsMZZuuk6LetwAtC1f3rZJ57e9l4gbsLQ
wj6eutp22iTjWpUQE5X+JEWRWwnnJTL1fJR04M5SH9NZLBBSqy3CsdMtrI6ONMoA
raZSGQNGnzZ6HI6aOqe5XhulH/hRV/HoeS0yaNXRTOV0RAJr3RchxmzDS5lVB/Lp
/QZO4X7qmSFmia53AIBGm1x4aoDXNvgsWv75rtWXCsc1bJTKqsF8+4JICiSnk60I
AYLo3pCyWYVn6VSs4IM/1Epynb7aAloJIHXhpMQjWFRQLNN4sFk/igZ1WRlUapv+
J/Benhz/J3/qiW7+TmDaZvqoh/zTzlc5UXH/6pyIkUElDsfO3Wfi/fnmVHrauVH3
KLR0X+I12mrD12MDHNo3C5D1whU6yeOU6nBOLNDFAXXpdiDDxlkEHcw68NGOzAke
tWFtsWCXG0RGCu6eVPNZgIEeB16EX1KD1E8E1QxI/QtppjuYnTRadFkcPtMLByaf
+EUrNq35uOHYIec2ditBSton2AjEQQ9KQkKeS6qYm2dN4UR10zWlf3j1UYB4R2tY
CqidCHWyw9sHe/14yhgRns0wr+9Za/vxyTlgS9KmpEqBD/nmbNNz4fR7wKS20oIN
JtXJx8g59PIZoM9UD5+RO6CxCw2oDbKJ1arBGK+FaRj4yVL3m2E1l5L44ath3Alr
9g8zFcECRxfxORqu2jqajx429gfeSoRnUncKBXctCfUSOQDuw8MbPQr55U8FIyFr
w4YYrkIke5OsiD/wiVN2Of9tuXQu4LtPsBmXm4vjrE3EkIJk/MQAXuVOkSYTCamR
ilJ1/RDsMONw0Lh5a6uZD3e96DkG2r9s859lKW3re/U+c5EZvT59AXIcSYFA+ht9
CUzRo61mkIT7dCpZbXaKJDuHs3sXqcxfwiFAUUbiznqdJHpzk0tWvGidnuEe3kXW
ihUvAYBvSADme+mIi/MkTEmbKG9PlYNv8tLFdZnXvHlOmQijibDJQxKCJa2ivvFM
ZiQO5q5p1wDXTvCv/kjq03dOgwT0eukEyxPUbN2ywColKvWOPQ3SEABQkRnj+DMJ
Sbg0aLbIEzBQkLK8fhxoyVr9AAamESJhHUhccBnaBegoJJhHj3M3DUKi+9LBi5bt
9wQxm2gvmHxR5mu35WF8usl23Gi5pZ47mXLlYIGsciXgtsU+pcjFTqiLrNztLb2O
2YEomuE4H/QcLOwD97XJPKB03sDQsKywgzgp3OAsAFaOqQFg90KLw9wBzMPUaem3
g4TdwZFZsxH+sIisCuCi36K1YWtUXan3pYGyqe7ICUQR/sQxTtwdy+MgR3CXFppN
vqPk9/pBfLspN3nGfb0ZR6Asu+3YHRLWx8Q5m9PcSvN5FmwADVUi36VmEq0SESkR
zvEv5/7YKrImRF5mZ1uGy96sq9mU62nPCL08fD0eH2NQi03vqDEDIyG5dksuuS4q
o8fTDxCw4MHXqbX7qXraEdiENQKQTpUMZlIkZTI095EdEyHnY0dWBtVJY14ymTPD
mUrapXqWthmtGPqT36o81S46tQ+eR/LN9dRiW3SdYU4nDz0SojvfTbWpygVRx1sa
lzJ1bT3ZznmgMsxqchzU/UlEexlOSYNaMPBschpwW4iA8tikagKuSzi1fqc+LLJR
5GRdJzqA7s9xzT2bSuLs26hDrgFoaB8KeIBheQKJGQ68osQfE3NJNP0Oa6UO3Rcw
8zzPrTl3Le4ta7JyW9gCbjQsyJ/k0aQU49NBy7FaSHpUkAU6yTtjfT2aVnZaPGxG
bUP9dAPphgeqfdHqJ+CR8dl/WL6RGW6PPJTnz559fpqwHYfN5sP/DkWfN2lBx+UZ
T5zAX5NhP6P5vR2vcWM9Ia6fMnGskJQ0gyfe8g+ghjblQqCJVxE8zwIf9sdEIGrx
4WXkn/Kn+JysXtbeWneUVCGJ3quPvdGQwnx3wVIjqw4S28bAVi0iHr2r32Y2qKRw
MqHZBWdYmhNObDgRPUtYAIBk10QWjAdxsPizCkbbELySfhg32sRoo0VceovcCmos
kGEqh4Cq43BA7xQ0UOs9fjwqPdBbrIOMbkZAFxDP68n0LsPRdZ7ItkI115AB/LLB
hYVO548EYZAtu8J67piQzLb0Cst3+NAbdtqwmRzMrZXcHXoqAisJP2X7nw4TTDNc
/SLhenlRBCOUUcQtXjzfhqV8h3yWWzHFhMmkoGEpcqrqdxJ3liHoQ/WHAA+yiNS8
NOQxs00VL8DprbJtQEwdCu4ixkAGy24VYTN1t1iTLejrKkqIZJEStM5F7Sd/BFVo
/oCxQJvGozIbX9S3Nz8lCgC/gZIHeOs6Blr2P3A5ZWmcmQScw9wo4GpnKvnAH00R
ScIIc6dnXvhiMn2V6c+e6hIVc9NMiSoD1JXvwhJ07pGP62YlvODezgUmUQwYMLxU
Osr8slRoBJMKXZbMJH6GUMKfgNG/BJ1z/mfG81w+AAtcGusUyyp38C378vP5tN4K
wMOKTycm7QdDrrJfj98Qd7IkpuP3EwwTlqe3aqyLCa4epWEkox+d9MoOVboWRxHv
6LjKUTPgs0BeRZzxmkcBRZ/m3om/uv1j9alpfpCf9IMLzAEiQNJMuSxcdxBNTv9l
IrXAkwuyCfJClf/rFsTRddfitUVLH2/txNC4cHn/zOtpKd/9OQWoxCyPQrQKt8Ro
hGfNspT+Nl09wty/74Iz0bYkG5SLR9aYyxFP+wJlYrmBAdBOxC+GXChEuLpq37oX
DilBbHoe6B94E3iv7VWtwulV8Ws584XFQjXotinMRp1FBafCIz2L/ZgPvX6wHtzY
27LtqaGMJbs4nQKQT5DvjdzElrcjYgQjoeWszR8fM3XOkswg7v5qpL9kCYvNmuce
bQ+yEQLKwQ8gJWqwELKjnCZV1Kmcu2k4cVUi3xIJjsd/Pkn76cvUzOOmfM5XYkFv
IqiOGgdSZhFawX/s7hzeod/Tl+Kr8NtZdRKtq/0U8GoQtcUa96fQ1mHVM2pqxrUi
zU/wE/VyYg01hQlqYSiH/mbPVCkzcbHpCdrOkmB2mCc6U3QDuzSBEJZTxNNWlMuS
gWM5RKp2UKNQE1XOtiUpVGM6IAqzrw1rMQdgBDedzPvlFXTYqfNAyhxeS39JQHIK
23zb4cQ3rOYNbJHiAxH/+A6wldOi3wpysPyyNMhVogr8zaf7NVAMnjWBZfiQGcZw
WeBuWhS5Q26MeemQnQe8EAuGp012F5jote44xb+wxP47TQSyZj4ljsruk5HeRIvW
xf+IBjL5XDZsEgcG9G/THQ8mUO1n0n2UuTG0PBllvr8bXVc3V3wHqaJgy0E/ZksP
jNJutndN3bus8vAHx6bXdYlTvPJY18T1SIOoV+IkVIz2TP01wBLtu9LZ9cmbF/kk
tzFCw6b5TQBXQeeDceoTmz0O+s3zYC2myN3Su+GRdOpQ/mDOgc/UeYTd9m2DXnGl
+0Yx9epiJOdU+2Jgwp8lfM3Z+sD3eyAl5BP2RjsGqouZc+4UCj1697qMXBd2UM5w
q8B3jKAH5w63onMfLxnZnVbQunvmYInO77vgxA2TyO+BEk7aMUQv0GduNEq7lT7T
z4Up9aGenNK6rDgL4wj5ybaXBHOeGndmcOOx4Zo7BfOFg0hcYjqxICbQomMQxpkB
4kGzx12LT9jFN48u5iZe20s4BLLw0ws+Gt7BmB/npfoAg7oOsLZgKI39O8+6w6nL
jml0PFQ0mP3BmSV3LYm0Kbo9rVs54ztB8GcWX9ee28IgR7VNGPsDh3AtYz7ZquQH
OVaBavFeloxxzSZv/lxOxmXqd+4ZC/PZoHRxJytCv1r4lCVw99FQxy7MRxSG2OKN
56co3sdK3I0Misyc7aJb++KCbtIW0rm6F5Pd9YEDU7uMZtvV0ZTb0T1PiHsormM9
1P2ryea5o4coaFSo0gAlyNMtt70HyxTmfKJDX3/wTnU1ust+NB+i91YbrC5fMYKf
MCwVH9bOJW5U6vRlnFbNvm3eTkvJhFf1S3VPrxdLCpIHQklEiMmQ1iFxCoVFJP5n
1K85y6VsYTmzcNNvjRZfYuhYBhUIkK6qHju3P0Z+tNB1u95mo7H+e2nHQ/4oNeCM
Jex9XjZmo2OwdMalYZYWiLXbujKGw/4rM3vsfZY3Ly9e07990678cILFUIQ6X/Jb
WvDq/FZdZLBaD8qH9ccBcoysOS+LJeT5tDGoBIcrswisvlNo+rUzHzSEudvZzO+/
Jy3HWO/vI+anD3H2TMne3cqjuVYunTXaHCH6+JuEZXuDP/QKfNKoGCj3De7a1Ecs
9JxMcHQ3q3Au6PpKw75wwjnSy/NR6tJxfHzJO6MVjDzvqFYpZKWuFj5Mvm9jji83
W7fXQ7M5EBcAjyojqTYiOlCKizwYxlgOoc7UJK6m6gKi/+VVF5HwVt7yjBh3e+7q
nF+jEuXafSxqHEfhwrpNipUgI6XbA8jiP4iG8stNa8JBsVHkfVzXy+dx9DA+fLAy
RJ9LxuPoL/IhPM1hfcohAqiyoZVOqAgTy8uLpu0SX94AHt11KecKjyPq8FTR3FY2
t1mJj/+gYY+NVq7ryUGGSBD9fQYXTLps7PUSEOeOhIPjON3WTEKELk6VIR/Qxndu
B6QGXNATO1wqoQqSAZGrUGIHBws+yO6hXZlPATVIfLJ0sEdIjMJnWfiFCPTw6c0r
l0DQw0lfa/aiefR+2mxQr9pHsAb4l+criBkYTPgy+JLKhTH/n5pKLxBYyww+gx4S
XdrbgjJJJzyO35MmoWpbBrg6vhWkgAWsBHXy9pXUZSqnMDhSNeaxA/yQDXSehxpM
+/8NkzFcaY+7aUVCM2X5WiPYiiu85GAWJDkiYStRF/UVwe2zujl6nSER3gwa7SMD
RpQzp2UdOUlq8G2kf2EucSXsYWKlSl0czI5c7IPfbNWHbPy9eipc1zSNhUuG/pFl
fFyW7lwhpVKSFs2LKz2Nr1+2casNG3yIFazZO0K5dzq+jYBzkYoO+EAM26umNkxR
gNhy6trvQ7Hy0p/7P+pFw8ti1158dR1yVrvHavd4cgkPydOxzc7pdoF0jB6/TXLE
DoLD0P2d3fH9IyRhXzhHSoWtsY3WAkstnd8kUBCJ5l/HZuZ/4yIDpfl1k9sLUVNT
mm07RKD2sGk0hMxVZYqnrtucs+R9ZyM1qess3opq5BeUBzjsNVH5IlVsWqj7cXUr
WKr7m7EV+6QOEPNiQIr6VUwrHD9Ohmn9lYvTmipOIKDwNAFBeqEvDE9QuC6xtHd0
+xSNvad7BLGbERFvCmLfo4SS7NIZ+tPbtBpVYzi1I/B77Xc0/RUGuCc7kPOitec9
7KVHklRXa8hkTeW5b/TMV/mIYFnFQGGHttLHgjGfX8CNtW0qy6tX7MFQknLMy7tW
FfF/sEsswWF723Sp/2gcYLqdeYZYKaD3Pgcgw/KZ/OOwYy8+zsgeE60GHSE7Ojqc
sw0U+E74/7+JohwSiYbSp7RK707fJd6z25ZPDi/UBYW+PSYuUbByYI5NqvjwZtf4
GquAEfdpLEczqY+P+agofx3NtsiHeQRmKayQzUodOWaYLLJ1K2J3/ac3Cv/7R/nV
tD2JXEeN1GMIEw28To9Y7Dr5KTa+NIuZQtgIMYHvzvqbdH+UpL/5rbTxE5wuqjxC
uEQV7SAs7TW9oeOnSkhV9s5+uTN9FvdVe41i+xr1dVAs9owbcopTAPwdzItlm1Kj
hjdNigqBZDnQEwlC9rnpwrI6u2GG3TMhFi5ZIoGa4bs5lMnLOC66fNFkjSs/qJLR
+gjqvYWJ2iyUtU3JF5Tu2P007XCv0QHGVfGuB5D+vMK5trfV69cMJAlXP3e4NUkJ
d4ytb9n6p6d9kl17xttqMyh4QiceNQKRV9YrqC6ikUpVQsFBcC9yzAVAWCnsNJK7
Q5htH8IpDiZybpKwtE44Vh3rdDSEPTdQeTaxcLlJIeRAW+kCyeQjDZJckhzx+oJW
10xoeu2WPgupKmYlnHiq+qC6sRqJFIv26zCL+f92E95pj6kOTacNHA1nvyC2OWDQ
/m2Cdr5KVAzvrMUzd+eNH0UBCdMOARxiQuyzNSl6ga6zdqwdI6lj7mFiUkanHy8J
K26Cq2EQrWKWskAm4aRtIDSiWFRe7yTx7WxE5+AbAfxN6UTMmHh5RD0vvificjsM
oBCcZDTuPmJjpedrPGXBP1zJUAJet83/T0RlsUQhuBQ11eDOv4y3n6RPodeEGJFW
+eBICOb+GGDLyIcGPpwL+HaPB7vHKJ8Ad1yriaFyYzGWa5VD/xUPAhQuRRMVYpu6
j18UI8YfSaZwUlqXTi38JFWdzEz6CIZ+HKiYVnSSSuk61s6ORSBxZgM1Bt46pKss
/bLuw21Plq11R9WrcnoO9pg7zwfcUc/ca90rk9Kui/+1G/r9QEoB3h9eAI3FB/4c
harxGeNex+/0Pa3Ul263YwhW2JXqQ6fdFEA5FvOj4a2VbPfwCW9tgqc9tkAh/l2Z
Oe6H8PARA9HL0vCCS0/lHiZOuXpJYqhEhas/fOhobWGlLVZ+Ibmn/N0gpBE4WtQd
Tfbn28Rw3621t1GskcZaFF7DVsW6g0pYh9WT+UVGfHMEGeO1lxy/JnbylY1mwtd8
rW829QFnXOzgz4dy7RRQXYefWgGzz2O24oyu/A3luaGiygnR3PUG2GF4NJCpcNEb
p7Nm7lRaJ9OJRJM5pjqMMriuxzGV+y/4oC9SDlBphSlYdhVBDHXlIRvfaNkRPQ3W
K/lw+0OE88yEbqeQKNVzmilao87qaam6Gw47/5FcH5gLzzacaPLBnoaPsIezC247
xtgWG15iVh9efG0TVHGveEjFWDZ22r+vaoIpkGfzlLN6R+j5kTW8MCbnOKyjEQeG
6RvqausYZwSzDP51bGXJBbo4PvyP/MaGhMi15X6+n6mt8oIdDLwyaOSX7ssQp5QV
x2rD4IQcNGH4PV35wiHyzko5OfmTFaP1uGeTcxaqorpcmfRhI0H82h5C5shBnFpd
zGZBGnAG9y4ePX1IosAF7ed7bl2sN0Lo5cocscggRIdj6GBrdMPwL7mtL8WBjTgY
6pVfkye18HGkgNMh9y4N2WLFnzfWMeWBhzuInXoRqqxh6qcHBx2jqh4lEWAWDKEd
UmXUgbaaRn0qfM31rPZo0jE+siIoDRg8motCGwMxVtCi/B+nhTJzpJbkWyNPGZwk
QKliy5bCsYJWXxj1kE1CoxrhWQ1ADQ5xvKMBbOirH6ixxbWd1I+LgaSbxnaxVQyW
jJ0guSoGjyjAu0xwhgdO7+CPtVO/G5VTa1KTntq4Sk1IBMFkGl9n57LEJ1sTedpb
oDreobJ0K9naiMTKDuC34EVuPEd+ab3b1j8gQKdt4E8HHt8c2gMQvocQw7/BL0y0
MKI+imXv4wS6eap4FmUCPf7K6sXKAIvfKh0FjvEC6fb8Y8COnk1NjwbCEGlr2vj+
2GLWLllVLOo8HG5GzJO8RDs+Y/OYsBtg2ScSm/uQO2rsmpz79r4YsuHtDxZ1iRhH
k9ipK4WQmRU6smWsGCJTjlaZuT9lUOOnZfUgfDqbEYLf4avhiUZDchVOdjikILKG
w7cPOd8mO16WESPRy8eIpQrYa+6rrVDHQse1b8iFR77m7RWolmdM7w+bedpLS7Jr
tHQsnaUqtLzNMVUGrN/2ppkCMEpxPGLe2tvWVNTCnZVWX6HoI4RuSWViHMP7kflE
U2rtAP5o5241mjaOU43VRcYnVtxNilWVS7e6LiupOBDzKB9S1CW1lL1XmuK0QNjl
Gzh7XQ+knKbIWQqEjqOPpirKVNs6xtFCbKy73kq5BIAtX5WlbnfydGT6cAGHKDt3
Ujlnt9+k1CR6xU8MUXdgszKL32ypnKsxJlGuOz/XZZHPofTZ2YJr8T2uGznnQAgI
/k//H35FdpaUIeHAD68/Cogfe/JtCqOlhYFMHrOBqmaolnndPr5fvkTNzZI5mwyQ
ohWVlKmWIAwZ/5eS3ShH7YdP07ak+Kwe0bdMPb9rMDSS9KKa5VdHEteeqSgGqrhi
TTd0uIUf9kO5P5YqXqMo99xcmJci+kxJY0lVSr23Bbnqg1k4pX6GwpkYS6xXP9CS
IfPqJTfxYVVI4LCxCyGvldtWOnLGs9GX4xV3ICXANa31gEBoQ4pZGXUgePpJ1I+P
un7dL/6JkOjnM75tycSVv7J9s4s/xik1+FtDvBnwLYoJ8Dhd2lToe/Ysaj3+I2Qm
jq09OeWjg3klrPsFJ3+Re0Uz9vhBmHn330WWBAmKPgJvE4La8qnybDIJuyNPYim/
IMb58YEXngr9qi8W84aOgg63tn7HYnV3cl58HTLffMn6hshHwQGFKK7tMOkpNtZs
fMZLRRGJG+m9Dc/3cv4XacVQ/L+eMmjqMJvQb8duggV9c7hJu6NDmbztU5Agzru+
5JUO+CzRRRkjdAPRufbaqFTHasqg23fidNISaTRuVrxz0+for9gVl15CmzYZDP8V
hQ7kjLb/Nxn6SYjzHIhyq6JvogdJTN2esix+BYoMOBEmxAke4TzqgbIiGLbzWjfU
jGC//r0xyNOPxKDZHX8/FU3e7a9biymvs5FC96YO7NVj0JnyxBF7zFU4BbLugQOC
z3NVK2S+LuWdGzkjO1GvsL5KWEyrx0a9sar/lcq5YlCKKW/l8Su7EJv8dOjuyFPO
3YH86zxE+Fr67ex9VhS2oJqYuKvl+aTG35DNyaj9GbJz/qDuXb6rLtuZC06e2Ecn
WtXf1YBJtKk86RGuKbLShkVVqLrHPSNhVwi/idHeT66VRMFqb4DKL145xFEV02Vf
TP/3Eik1c/0xjINV09At2puAbVGflR9sijRTvJ7EBr3KG5+S/VLsqAaZxyBUhG+m
smQPiy8j73C/e76n7zOiTMxr9mKbHpHteleZiNLXYX91wGo7uY2UD4zTQGF/mAPy
9kbRMOPuT1QUD3/OGO37LxQ2BFlCEIKCT73e5Oqg+3ZsMMgBU8k7MMMLixRpCYuO
ZDcrfofRWpfxCz1w3ZYHvzH17LzofyItCaniEep8XdMdN+dZYhCi8p6IDw7GbbWb
f9egOTsQLCaL+VsNZnj3fZJ7stvkwOc5w9ozXmeUGKapmjpfqfL5MTtpdt5mHOVp
eisRRPDDpO6NBO97izBupcmZ7hK9uLQwGi9k1bvBcC2J51IUT7oJfCkgJNeRkCGg
AbcVVbyIJ6QafNnZ2GS65uRY2QObHdO7RoshzZQpkSBMQlFPEKHwLQTPYsYvnUVC
ynv6O87rHxrdkA1xLik75C2At0sOfZMsCtyLGcsa4JDE3bdSTfgYgoYoiPbmaSp4
++SsmLYDq6XG5PgJ0meOvrJEYksl6J/E5zFNYGxRLBRBCu0sisZrMu7lsEysle3Z
e/iVSTug1H3LuegFmXIacy8McIW3mPWPcjj7PjE54jBryb4RbMg4VOrPHdHqQCmL
X32YTm7kj95/5jd7+JOxVgDWQCmnJnfPveH+HAxbN1zDA0z1dGJgDCiAUWLaJ22u
Ara/Om5ZnSQFc+ZMJ0Z9DsKuYrv4xD173VTCEkiCCy0QTDRHGGbg0npOYxsHDoI5
CS0L+zILkkXDhBVLbUr4rj/yAyZQRzeKkPAXn0HBEV0vSaWpWhk9G8G5DWsHyCcf
41/R8UVwVBCpiKYVmZZMlzfdirapKDeek7e/CkICcE09d1ZrOTsH7qCY8EhC9Vbs
C5LB+tbmv4zbAULuc28iGuVhConXszKWa+dgCcvAwIyX6KV6Vh7LtqZRF29azZrd
KMB1Edk/xdbeNWjzvY+Aw2lfkN7C7YW/RP/3dAT6dIKWgqht7xvrGZKdZyLYTH2b
/wlUJD2OGchaGGMBjjWKk2ze1z8DShAxWPRR8e8Qj2cE2pXgO7ynyOKLTnq201s4
uktArLLZEk3LFCUsn5IcbhDrN9e1QLjeg36UyPSqTSm0N8lI3GnFvRwxgrk3jMg2
70PEV7tjgi0AAu3IBplIcFDX1e+7cbkPdfz9lIMgQHio9lvwg3gBLvYDL4aHIrp/
ryEW9riGzQ89JIwXhX8E1ha5sz1rz0ZF+YX/QGZAjAoa/2/Y6PzF+IF/g+GHEvah
L+qTu+/dqlqwEkHbUWjxcoO1wCJwLvX2/PfNrsixtwBV3Yjn8aqGZI6E/Ilo844J
/kyBil61O+2eJSppnU1zaPsrfoiljc5pZrmknawva0GRg/deQFcvqgVmPmZ5wFPr
9GkrPEJKNDmDmjqe3mqqRY42DnLioYJrGL7vpSrN44VT9LBkluUJD0IA/wES9xbA
e5B96imoYidGC9+jFCKW7+MwB0vayR2ZzNMGTnuUmZUyaTgAR/tTVIoKx56V1zCV
A9UBfeM8Y5ChgM8hJ6wfyDSqR6ZozGV6RWONz8CPQpU587O6Ax5n9cxUAwGJwF73
YfUPmxr2qE7Wkt9S7jZpZ/yb/+YMRLX+VggMLUoduMwanTRjDAcR2yN2HdKIpFrB
1HoOb4xUo6jkY6X6hL6LTOkrCzDNhI28RNfyWKhZsfnGfpxcO3T8e+W25Yr5JRS1
uTIm1ZPet9UA1iTPtYSLOHL+B9uRprUN8+xMIe/Tk/G8jb+I7WtorpVqSH2tpYJR
KU30IqQKuG0V2vaHRVBLrsHCyiElttjHpabYd4dGV6tdPsYJ4I0awAEYVpWL2Zi3
bqACHJ+NR+B6cYcFfCd7UeqZe+d1oQ8NPRAl2PWAHCjQc1KbHxW4Fy+Z7A2GSkm1
9ZQYThkczFFBLYN8ZCsPFWxO4cy0wX0E9C+TcovTbtYE79yGRVdffh7AIolxx9H7
X/gEBCKfdy7Tp/9NMZwKm4LWVKtKeUrUPOfOva8TFnmH2qv1gm3Iqlp/fUAtSALj
OQGWSxu7VuEnxJqQLxfQxH/Kzc3OBGcyXT56EziFUUOaew3RrID+fNBjqfbrEalj
MoWqj2UkrhhVYzn6xa7XTIGeUWQPfVFYyo6I2vGwuMA4Tc9bamRPy0ZwRvkSBepi
tl7FM6C57MbxsPA77UXW4357USo4zG5j8cQ0Cn6uRyiuQmtZQL2JHd44ZBX9SBg2
lznuf0xsUWC5qIo2wClaOkRl8B7S/lQO77RFbGDrNKcTuRA0bRcsQ2pwwF+JQY6S
ioBVuMwIPjiRd3mDUBI1kwns0qXpPzsRbzKh2RqdQxsY4qR/rzDY7MdL+JWNezLj
0vTpX1rh8HzsAFW6WiZ68FWhuaGhtLM87mJTZMUDCFSwdpEAZa6Ywy6faHQIWSCL
WqYVR3Qe75ibIsedLY67Gp9rUTaOZAdg+y8Tqr2BsCYxH3kXdAfZcAyxuvtWUrJP
F0iEHPuMQkJC8Yg1B1b0tgTYg1q70GgN7V57rsR+MJXCw+ez1qY0r+xF4X0IcIgd
SrYWfo+G/pqAwdSBr7NxQ5J2cWAHAlsJgp7pmLa1OAdtjzVUitd8uQrhdEc/Y/tH
UvIcyDBEVBUXnxMV4+VCCrP6ajIwwPtRgWJJvt6VqwE4/UKzz5+P7eGAZ6yKRNV9
KKNCycJuymlPIzQB18o7ok3aAQVCw08GLZ5WqEdlhyaGfR2UM/eB9FZnFmzKFWdm
5r+Lnjss2zH9QyRY9EDXNkZF8rC/sn2zTMHO14VvlmsuDAZcL7hT0LGjtp73ey8J
gx+74qy7ymga4PbH20BzL5yi6CeNEDLQ29amN3HhiLY+oVt7OXgJqOxqO+INSScB
rSpTYVDrDqwBiw3xdFKJAOqFnDMpYn9rk0E9xEsafz3Psn0vdE7JW0XtNuP6uoZO
REJXXik2Oug9TNtcZEghEvZKzZIt05AsmMPC2AOo64f1JJlriADjij5Ed5UKoQyC
KfxztC7o667Y8nq27cW80yC8ODDPD98dr4XE59yvUQgUEiZQpPXAkQe/Be/TVWzx
3+h8S1I03RyYgVUZu+zR39Shvcn0gw1e+CLOZKR+1aJeNgUC/tNR4Hpj+8cWjwHp
TjU5PaMypWeh8ZURPpqFLw/KgGZjbUnc8g7UGC2aigd2VVG6cXVKm5O9keNtZpJg
QElqsaVVWDPHyof3Zv5x9pkyABsiKK6HAnaU4mZMWkNEU6C8+YVmEdY1H88RVfIO
h7OVCZJHeoOduXpcPWMlO+U8SOMcdOo/rIsikzVHb7SwPSoUBX1E1/qeXGaTg5p+
ck5A5GLq7Kk3z1jjcp9JKCaiNT4WsSkib0QlYwpWOp+HEO80FyPicBzx8Z2IZHpc
lDmP22JPErO9gndB5WYvTooIi4o5d+QCGDaectG0JkMGG8WV3VmcYUu+eH0tkOIR
JKM2VVtBKGlZNAl+D2pxHN+qKr0M9SmpR44w+ZRaZRZLqozGjYPVYd+o8fd8e9XE
28ZIRjKHzNZxFjFCBjmdG2HoKz1a+R3R6L/A3KOZqfnBAlHxlIEIC0/P862BDPN4
RYyEk3f6x/sDnt0232uAwt6oQuXy4wBmy8kfLRlZv5wfhrrZhK7MZS1SjoSOFjEX
Xf8dJHIoLNCGkWuC8MX8B8wU/cRbUDMp3BinYa62frCJKCOsC0sYknvjpsE6KQ/Y
XG/62hfyICQqfd8DUJCDwajcRXoH/vrIl74corcFLnnbGMzozeLgA1Zt+chx30zu
Sma8nj7GlS0RLJm2apOsJ/D2FVg/V2DaHTuLC+PYlJtJkZDUdsrgcVCLQmxEXyPs
SgC9eZ9aHoaFHsT+JdZX1yW/3M9z5XXWhEv66J35Gg8Cw0Xm2tTOu4GHctja22ZZ
HaeGmLYMr1Ot3qYR/MvLj/ig6xgbjbtWGCMbA4FuIFX81C197tTmShCfJk0CscSI
IMFOzqx/qy+M5yooBzyhBe/F55w/+rV5032CZA3r7pziED+ZNSRrYwnQFOFviAKO
H82I4Gdnw9w9wZDZPdpx5IRrf5bFoQzNdnf+E/qcMUzzDAHSEhWkRhx3KOFNaem/
MbSE/gL6PM/FhnTREfRgXafTOZd3z8FjaxH5iLgFu8bF7wMEV7+uJz2uFU1myEsu
W3cU2ez60NgHF5TpTsqfz1a97byrCkV4PBoVau+9LiMu0/1OAsAy/K9McS0q031U
MQ0176zg6+1g8gXWHnA3mwOn17PBzc9WaoesDODyrD5kBf0RpC2WdjaDHvV6cEm3
mMv7hzMC0szwJYywCD7bTHkoDxhU8vJsH3p1YmOI8AhSlDrYzy34Ut2j1BAIy1d6
QPgXT5e2F2pwrNI4B0vpiz7Qc+NtZFDJc8p4nQpsQzxUBwb3/Je4rMINqRXkzm6n
ucvba4dfWBkHwlbtitu6g/Z3OqwgaMHxrq+V2iEFvksywjBHvlGM3bxcFDx6JG2E
00kBc1yj4OdZhduti+mKWq7xVN/ddbqoTch6CGSlsJ9OnYp0axTttjVUpVFhsyaD
HOaKN0ub4byvft+MLqsIZCuLq+uK3J7LkovPkg5W1qv7wqRDshloY+Fbn79JNZAd
CGxnLLtk6/icyq0iusHEVHgozIxkHsAo7wtE1A2CkjqwFSZaB/s0z1BEvIOb4J2Z
PhqSHNzavSmx3tgyZAg8ru+JhlYdwE9gUnGaOrLOjdcduIHg29J+CWhbMY1cSDMA
K+5nPi5jySUhJSVwjnf2+WUnnQrDBB4V85u3tJl1dmjC5ZHAuOMxQYa76RC02oxt
HkD1gJnRheozWIBWrJVe5U954u3l2lew+gDYI9NrFKSLZJOwGB/d9I9KQgIxmlxU
NjBdAOwNK3XW+xts5ErGT2nMYP0QoKN0oZ92M68Ro+Rqkv4x09wJjnEhUTIkVHMP
O2sM5Cig1AT7/A4H8M/IxK+zYpaI6+FR5BOQLAmDcJp/WG5aq/BGuEeOZieFQLGM
uTKkRdDBYFJIIMxgne/ljqqJ2OG5E/2a1wlZ70d+HHwZKb6Mnu8lDVzzdAnYouU7
qUiUQRgDw08ueVt+0vLEs9+iXyeatQJfXt+xacmmJM7muDo87SPnqCA+zTzU0Ni3
ZfXnl7D6ZePMw76WDgOAJZ0cdQlreUMB67ySGpLmFkFZSnza//REriK7HKjeMtui
1qPuCQrhUmcQ+KpQxxscLPjRYe2k5SPqevs1E8m5JIzXROtCxDl234/Q7ChBYiU1
17XLnzckQpkr5J12WCIhPFxBnZQGXlMez07zZ2HiW/AYvu4f4s/E5z5djnT9B2qU
wYRrMMfpW7C+ws5vP9vJ4iUJutfgdrBV946KgmtatNEDd9/5MdWF5oeLJQ1aPbRk
mgOeHkeeg3lbELI2hTEt610SGN1vTWaBLCd+xcu3VXvw+zc+/u7ea6oabAxjW4Cm
z9uOA03ATj0mlj7QVn9+1eFlBdpbD6BBOmAWhkB0ZAcV5Hie8eW0RyTqyChrHK+B
p+xd/+2DvSzZK/doqNc4roLeg6JACqO2J2eWLjH0RgE3qnkw2N/cF8eSt1q15sOw
NQRbCw786yh76zDiIcEb3xvMxJwizzW/ZKv2d0uvtDb60MlUyU2J3R4ZSSjq4pyU
sZNS5iy2edOOvleKmEOf5eG3ehtbRIaBfQW4Res9YiL1r70hj7idNczUJv8PI8M7
QHFmdxhNue/bsHHzn9xbJ6PBmLwO83SmaxNdmxurYxHw70x9JOojT2hELDhuae6u
Hhv2PzJ3hscs4NlFcCJt8+Yf5GlZ0LbUNx2RgAgNMfPTbdOSRvbsFtSiqtVlbRbI
YgfMrcLnKZUnU4ZcPVUgurgU7dQZc9DD7ofP0fqpm6b+FrfMADEv9aYdhJtG/LZL
7mY9SfU2wEuIQDj3C+UdMov38KQGuYwgFjB+lmaDQN1/oAq4qNs28CtphuLeh+km
o8SifF9WNBFJ+AjwgHegEo7y50r8c7tm5n34eNa5aVmUrv/6AAtqvcysx7/lBFej
HpGDXzFH8B0yDvcSUpygqlaM7Ch1I7c52wDDh3kIgNX8+cbekR3KQIe6rb8NnOHj
d76VYXmbJyLLAEPXUwje6V1xVfIUEFe+oEx6n0JXTEyqYaiLZQxRAx8eIj61z7bR
AD1t7PwzaJwvmFK8xn60ZpWRORGFP+O93oH1775Hu7b9raQmLVpepnDK2EjNefCO
0KqJW+wRiWhoVkpbieI1+AbfmdWGbV3K0qaYsJDKUSYBdld6MMuEzTFYPFSs2ESg
/GUr+p+P51Ii/vbbiRKvjAGEiLiO9savki+qc5Vu+Eq343u1pG+duIhsY+vGAqnr
dSdn/L1H1mh75/f6LnDULBNRcu+H/QdvUyhD8DtSL2q/1xm7hiuzxQqhQS5QdA4I
hFIAQrO5/salB+iNcqeX3Et/cF1nsVgbVZGXWJkjUQ6ksX2O9irmFc46ddrleGeR
xVXPukU1h8xLUIJrskxFgG7H+0yQkqj1VukbapHCnrC9R2WK8dhQoy252Eng9LWq
gLu2Ao6RkrPVTAC7+xP6GK4Uk7FacL3G9oYQyv5sfxadQqd1ft93GZSjs3ojstG0
4VoQR4sQwKhL0dpodDHOBxAmfr5XvuvDXmTq8YHdEAIEj0hu8ZUiMepHqUcOObqG
oDrDHX15Gf/cuq+JEMZy4cwoF9rj/+ZxSBFyM3xhzhkFA4rQqrXA+1PtIVYK0W55
jA96za3MmX/Wp6kf/xEz96jPpeKIx4fo+U5OGebSL7JkPh+fKnQ70USCekPE4IqQ
xHk1t15WpCGM3H3D/3Fv4Qzi2dLEXD8ERRapZvFmyJlOViJErx2Q2XkXESJSi75x
gBH5oSfEq8lWG91LLEDeCPo486kBBDHB7AvAu8Y3UxTxPtKxUyE50+YyaB9ZhnJa
YHZt7pFRSdTuKSrV5MY4dgFCl9m6Toaw17aDKUCC0msflnm3O8eHU0Q8vOsNN5pS
pZqV04WE9qieVrKmQYXqmymzgST7ll+c+26pTOsRfZ7a8peUQW7It0TMIDHyg1vi
6WF85JIbyF4RVqBUXLGILQ87XXsGY2NQbfJe2Kj/56CLsOUV4EdXnVn/9PaJjt9J
s9gN7wo+NvRa2zIBMWHH6pTyztHQdJ89zjprWflq600rJyPzZhWQhkoUn1Vbn5jJ
iMos+0hvkc4p7x8AwHE8ztqD7a3skvJY9aT74kpxSZsH2NIWhtUPLzizjLzulU9F
O/IvwTr7hGQMOsry7aZvPjWtUOHwYeq/hl+9j9DbAv3iYIuC5W778CwS3Dt1vPCs
K2qp0ZGmGdODQwNSTnUc9AA3d78BMSB08FVMPAbt2s3ooi1AbFVddzIT4T5BeBIv
bwFLDuu+DldCBE5jInxZwKfy9Wl7gYKhtdmx6jukwLAAT9/JXJdG5J0Xz/JAkHSV
09D5jI2GRAqXm8h9Pnhmd61yiAq1YPHvhCcUfmevqIJG905j4P3bJ00G0mh4PllJ
bm5Q8bg2WJRUxHmM6ss0zlHei/KOafXsKKeB3SoI1yKHnG9nJ8A/d60lOKhNKxx0
RfwpNmifOP7vJ8WkmZxoLO1XW8cKASaOllNq2w0lnurZa0UwOqVpMeAJ+KiC+JJ6
RbdvLhriCn9T+bcvsYUSo8aqTt67Q8HjoLPRkXJGL44EtYgOuc9Z4HXAR0ThDFE4
0l31L/eYvQGPTfqhzbnUClCt1+bHXNI6CaXIN6KZwdYaAme5byJvkCAnDYb0h0RO
eXLSvQLliaZrdT9MYAYVK7MAX6DWj2mvg23nDwBdJKwDIqQuTtkQE05VB3t280zm
bmAXDR6iborexnvx0WGvxq3UOEb6fujdWenA0BpMcXWuoW167J2kGeCbf2L8V+Zk
dqyyWPtDF6nzkrr10112APJb2SFDfcvrUHqQyXh5D62tLs6RMZU2Rm8fd9Oomm1N
hSJdjvl/i/UkTk81qsTW4g0WfeOEXqBe64RQcOCefGVs2bsi1wnKHH8q8jUkxmpB
7hIVKxEEUE+Ji+J1KVhyvkeAsM6pi4+hkEJ3wrEftSDfM82xY3vkfPK2JyNmWvh3
xjpkWMQ8J44v3LsBBFVAPU5HYt0BqAycv72QvpGndbiGrnViJ1SREYwNN1Jlzj8Q
egWSJ5PtG3zViziI1k4XDWPflfG9zaafRopbaR8B7DEKLmli1SGwxHj8YUQ7yBeM
xGtJ9UeruaNxzYnieiLlbggjvxiLfBKHBDM5d/ZjhvtDdszfONlCKOlaEldfwS/H
lG3uI2TjkkeO+IK+oyhDZUqIp2jBL5OdV+nLMZW2uGYuudCSE/HFYwzw3HhmfnW+
7reAWB9MrRM2HLZwLLcMmewTvS1joaFtrX27etUTwQy/ZU/iIDRMd4cUA12Lvzxb
+JHvEu9iv7HXNjuRC61H+witFkKSlA/q/apvf1WMbw6hx422KHIfmkxi3pcwjOfL
YsEpZD3fVuzJHsnNmCRqMLLvgusS00PweUuKR+2LhqY9Ux3nYCNguWaEvd4dtKtw
TMfuihnSOcIaIt2NnMsrIAi579YWs6ZOscAWIPvJEbbD7oYQ3cSmAXgnoiLAPx3m
t9RzKeCkd86MhUEbA5oQUbviipl9gt/t5XH+hf/npJaowrXmHtAU7a1+9/3/QbiJ
qaDeCYcreD/ZEdNe284tPG72OFaYNi0+pKlyDikQcY1VIwZWB7geG64Cwyk0lDgu
8JavWTl4Xz/iwtC8oSR5qlUYzex+DnIJNrcoKnnRnfnyKBDw1/vimVTqwf+9leSB
Z2KzAIB5PaqAS+myN+FAe+bZMDc/hiEeT5odLVCppvfjZFc06OQvqGCDU2C5rfoX
gmgCA6LcXWDjNIcu1amwryEEauWjrZRtNF27tIMnpfuv9yNxrPCTMw48KVcdeD6p
wlh60ZK7cgVHp+gtZ1QSq/ZyTIS9v3vB5OPE1aBpiAONC0JPiw76bQfOaabMfswv
Bw9QJMUYGWYLaVyJdjTXkWNaNIduUpEgC7sjJUWPoMuUn/jGYoZh0M78m7fMEwv5
Zt3Vm/TfKfrI9krZLC05jOONxaiTPbPlt90NdmbtTfveKbqOPn+aLaQUfHA3+Wwy
zPRVzKWSiSWftZiS/1m+2enouz8MDPjH9A0aj7bGLKYUQFzRicKGbuGU1ltyetxz
1b+2IJ3unfvMOc/NRuhWz/Y64TN9uFaqT9L+1k5sZIzeLEobAHXoENzjscnjXh/b
SO/ct+M0tHWcuipe4bn5PZ3rwiNKaKSmD71Na/9VjcZUTEVxU3go2uqIPSHFyEwq
jXruIQH8K6rrZYAhSAlHvnhxbjIv/hQCqiRkn6ETMuyKfP9sE/q53d0UuCOGRNLu
huSW5aYnRus8cZSXHnz1iaANRHlOZyVZl890aXmny28fDo19EMJ72PRW7y1XOOyd
i/fgZSOu/bQX9cV/fx4yaHRsaR3YYjUcxA3IYBgpY9DXcrqB6oBfPvB1gQ9c+GZI
V+5xIhqNKuKYgp1muYIh9s1hCvi75D1XWmNzjCPIT8xKaUvePXBB5fpMbQvvdKgV
GVgx1DtGnpROPhQjxjSAyZ+7VnWvGUZRbqWRP0qjjqfwjqGznUnsYrb3bc4YnSM8
THfr/aD034/mIaicxdr4T04FYoHJTzgWD6ni+USBCEJd1GpEjwiIJqWIh40+DtNN
77FJCKRYmPA9kHYM+Y9jEqQ/WAinibwCtaK4v/WbUrlpaTd0W2LhWpdVASquf/qz
8ryAfzlHTehXMhCA904PvlOb6re8fX4KinGP2W/cBOkHY641EzEACG51pzHQFLOc
DJ8ang0SxaqU0faKd0G7tBA+9197dgRAqTpicaD2P7Pij+xpnJwx9MDgathzvAxC
cuFJi5eJGbAmrX48SyhySh+ovjdb3bhsRNGBSKrPx4zZUyMLj4jXDy2g9KkSn7bM
JYfKub3cZOoE9JmrwEzhCkyAFqdhcUDbqAmDhxcoxHIM2Hb2PGPdJpIEE3w6Z/ER
mGO4YP01vqLFdAzAWAETkDqMTMh4cTvFeUfKOni9zag9mQThSswQoyWlaInF1Y+k
HKz+E6fZRk51wekbauFkZ9VrUKDs/+oeSeTkBMsb7J/DTr9JjMdGkmmTQ/0cllt3
eJdnEnA5PUo3KVA8fs0yFaKuVyGC9WJmGhLKuHaDeka2w6p23lzwaAEdobb9m/z9
nZlUVLX7jKjDGrtoSPjHSIxt9x8a37kEP3CW2OzvUNjHD44N5lQiUwRqlYl4V7d/
LvlGje6/6e2NTdctt65YuCTeJ0GDokFrwMDXt1AHgUnEifaHigI03f8YRSqWkAJw
Jy6unxuqEpeStYDghpV245xICKSk0i7r6rJ/qqMETbXuTGqY/hzFgoFyY/eRcLdM
bAjhAvtT4cpw8fRX/EBRKqbASu7vgTMp68wgL0lBc/5BywTExEG07CDEtJMimbZk
8AXIRO5xzyWlylnkE7Vjo+qH+UvBgsUJ7M6YOj6r8fUHtPtRrBSUAADNTWNcRo/E
okq+qT8OeSbToH5yReffBB1GKd+APn3q1YpfMzk2ohZbFLNEm+2+4WMDtV/FOJxs
tRYTxqA+x8ayMlV2HabZEOike19e/L9E57h3NIXOqUfLkYUB4cCRrHXlg9/dm3K3
hrIdguplCjtLI+ZhpB2CZdyL+maqZprujSJiHP24NCfZ9AG4mKw3h+nrleqPU62p
wocubIHOqhMpNvRjTVmBISBs4mv0h3uf3zM7t5xTGg/QCkVby9leot1CQ3mU/rV2
lJEmwWr9wTCdGKgKIUTDOzOo5nd+1aR3YVKID/bf5/7/lPVxEogxWk7TFlKqJOF4
XiMSjT/jUHQCGX5f/ns1lzh8+nYcjKGEocs3LvQTMiMIlWWjt2cVALzIsf0OvCrh
DazOopVSM0RhN7GnIzuxFj70MiJ5dMQSQtrG7t9ZdItcoGTEx4ABuu5XLtHlRGQq
uEzfjBoDh4S5QAxah9Z5Dzs9wiO8uF47daiI+PfcOvNovb4b/POYezVeyQds+sad
QCpBvheU9yomQSl36dLHznAnMFbpTmM/U2RWnTpdkssgPfSkqiSTBEbmN6zLCPs3
JKW/wNp/x6YQSefkmJmLmluw8bNhCTnJyBY8CrggMfQUF2i7u1a4CbqnyB0KZdxr
goTdXE2izOWHYXz6A5xOIboDRFlf9D7rg86+8/YLsQmOcns1Jp1j8/+FrKjWN0xU
nCHHBWnGnsPueGw0OKziLrQUIXx+UGl+6f7uu++ATmdx7JMXO2jxmnzcM7kbNtsc
URSNbj0Up1yV3PHFpq62JgxGuDqHsp6PSj7RXkx7E+37w0sC9iv9qFEAQbgLUGo2
M9QeTX6udFikm8QzipGg69CltcXheOinKBH5jpU9oZGXB3Kr4sd4KG+vJhN9xxqa
P0oyGUbTXJWBGtVjR678WGKWINlRf2Z9GUnigqewhzUEEzpLHmbV/i/xYsSZWXkg
8BFuxNmdzFL/ROCnyPyJev5S/C7gcfkrmqXQWTQnaYOnbzlHbpb+7GkhcbHsCkWu
ihzdZJnzztRlb3pdvEY86ptags57ckojAh+SENNcJgJBwrnvw4OOjI1YihJ/Tgpg
6S5SlIJTYOGp7gecD4gpCNyMe+91mjBg3sRXCVnb5eRMapBt+wDNsoljQ8B+Uwm0
NW0IW86AjCWE4Mf4F/RtoEfk29ZaXU2Ha9Rz4ciRUhp5deVGQYHIXnagtduMFQRQ
M631UwJ//I15DdI409zjRmrV8TvbBdpnr71PhA0BqgY/AjVDFHiQShDdmg07MFWD
PyDQdfY18/sPaP1me53CrMvc9+myLC2IXAhHI646pj6af0qSdGa9P+AjiC2FJ0Zf
3OwuiKZtR2cLxsTVhaWKexCscQ7ppLMSrr0tffTiHvZjOyGyqXPdn0A5FIsKoS4W
67ce3U5bb1bzuz52X9UBTPgAwBcCGSgndkue5NNroDtdHYIOUQKK0j/AlWZkOa/k
QBvrpIC6sQJrVtXTNO1Mkl1c9R+nhrq8Irl/5klvK4mMSjbXyrNm9csQDUkNrTHm
KMACXZq0AnGnpLWz//fGg6paZuj7UnYQ2ECPqZO6XbB6gNV57p1QbqdP/h+xldDT
F6wJUcCqxiKytc30tBP0mM/98zK09kvaSF3MGw7R/A3pwSfhnOwIdFV55cOH9uOy
v0GytQpKy1D0nGCawiMf4pvm6j5YDdJ5rGQ2X6XohWelqo7fBu1cYvSBb/XY9LDh
gmvP1/JJNaTkmPh8VOWSxETfB2tGl+jPBe/ST+FxJA4fYl422uv3tplAzGE2fvxQ
Yf+vJDMCGC7fjDKm4vbmIPXmY4ooDQvgmB7e7VFElLd5IhoScvm3+QPidHA5z9uF
cxOXyFdP4OxXZOd44jRJjYJaw1KTRIAEt1UMP4MYECntHUBIfHdH2yEU6VjAvj2u
EcOgYBVNkiM9ZKmKIV12Xq/bRhs5Q51dc9Fdnx/6AmjlPvWZfOzj65xXpmEar6vM
Ek0H9Vh9Mmov7/Q1wk7NcdyGBCV6pnLKJ3B+7ulM0z4Hx9WBYFaS6RgqeBFpi2kZ
sIbpG8wU1c/VkdjL8OLTsgzeWYipDRmBEjaoKSrirzIvRSQaqREmMPzXk1+hvsuQ
097t96xkRlsVAgtuw0c8+RiUcRLXvYgJfYuyYcEA98uGmx2ZkdqANEzh9jgDYQ73
N5Hlo0UgGlXzNgyUEA9T8omMwxWI+cuR3yS7Xds4zBb6BM3M2BSX6ts08AVsyMd+
W137sNZl88Se/sOYB5NJs2RGROmhSYjw4QdMdltorJU5TrJk+wBX6bpjwTB4izzZ
7P+oNir2wsBRWwbrbMbodZRT5yixjj/i5afUAn+2VPu/lXRXtoSlokxqPXZzly+1
1N+QudjM2tUIjMcL4YiZrwQccU+CjQmio2pY8/D8zMAvtzFMXcGV0n8tzUczPAWy
gw0hhnSTGI57no8qgjQliJ1cRJm7oCv7ID7gRni5nX3gzsnDd06HQKxThm7hJaUT
/Vp3wq6OkyVvjAycgq9vG/5y95NZmfOTrRPkxaob/NZtCs+MiUczTIg0AfrG+kdU
w+8+uUQ5weZb+6dHKlYPXFr/yPmn5fBuZsvsWSCGNoxAB1kRDsSCFnRiVyPlXHax
gVC0k7uOOI97RvaVNKR9i/f/2shTWBFA2VHohmP8dP5c50CX4vQhjJPNB+ZJF8vT
QA0D4o5UV4h4uCJVk37vcwmqFQmFFnDZozdOQhI4XwWSQWvyOq8ONJUqZYmWHNjV
feaGkrxUJg64lILJAhyML/4XeBGpOTOjwFj+VkK1XxSB7PKRuQVEZVaMZE7ReNOv
2I0+iGUobl4+0rDqN4vRD8qIX6fRh7C79C6Va7LbTGG1EwB7MJQJSW4QVXLwWD5i
MkxNqCjrILtPISUxOdkKs6hSff9/atZuCDPdV30zVZSVn2m5kzjUyi1ILL/hxctm
WHOflCEKZ5Jf2xswaMUG6iu2Bfy8d7T06zr/9d0EPF1Bluuul/CDxXKN2JmpY0PG
ALHwL0BD2r7L4Py4MClHTkcLAAEcGZEQ4HebZ7ALYR1MTiQhc4zl5Uavao8Y8Wwu
hmtw5l4Ig4MEbPgBvsnBhYYZhv6ArFNZBmALkxHExmpR8FnpkwZWy0HZuU+qRe1b
4qrB16sff9QGqT8G5VdnlgMqcSoDE66B1YqyyPiFoSPImP5fT7do4NG3jvRV6xC1
HS23lrT4U/yomJv/bX1srAJlXvcNTY7lAndxxtY9cUJyh7JHWHt9tig1HrULufvf
QaODRgSJ6F8TW7jLX22deICMbr8JqlKZdLlFGJxdZbZQhEjgztF3BFZo8pEC3DdM
VxUzSurvKKdluTJTZVz4YyC4zfWaqUWAx+fZKYpAcT9lwFZPgviabgB1izzmMLE9
78oanxbNO7IlAUszpjGgLGtqRsbXw6IqJYVurEnXavJivNBPQEc3iiF6DF19e7u+
6D18ZjBrwM9f3R2Oe46xZzCeisWoTok05bD0d2HvNSsErDiAgBeHJVcN0mrlw1hz
+5GdGryTkxt+cK5JiW89TKcn7hXf/DcvegekPE6fvJGGBPCxLBSklLAnupkdTWvN
oADy4sIhxh46dIrQSSPIqzyQyB7JMskAcNJK7U9u/VcHoFxMyNlgBw1ivBDweh5f
9zINWaoiRJl4Hl4/m84JDHILP3j1ATfEFVwCIOEFRugipLYApBdhdj2IDhU0cgDE
7+I20PvXDhvCPj8Yz1+xaVvqUDCUMGLNaaG2JMzstBDWfYdstQFwqwWjk/5M0mEt
s9mcvfRsuOKSutDIoq6Obo2UUhZRzYZ58pmzBJOYjLxzPIyREXvVdLITYB3HuJ9L
hYK+X45DecEYVKGMR0LemM3Oe4Bc7tQ085uGCF7wmuwu2KEA+bJs/6K496nViIzm
LmcKF+DKNSJEnN1bCQRhKFBMATwjkipXfN4TVh4yeyavrQ4VtOdI4mSkxto0hEBS
SZL/DcuiUF9JTs/Qn8PL2JPNnWDTPTOkhHOUMrQdaKeSq0t+wak8xFGqVlPoT6Pj
eNyc4IeXHR6huUQnMqjYpM0e+fNiXS75Pl9H5RmmN9G+nBkHTQjTTHJyxZ+eeepv
nZ+Lmn//3ny5yLKV0/DaTnjDtoNd23bj2oD/Jonh5KElgCYbCXaIZhFmJlXbAVcU
k0YelZjfzVKmVvpefb40ffFXWKbbU2+QGAkbfkXun0uTqnJLois1QPx6IPH8wf4d
fv6rPBF+/WHl0JlIIS9V60TynZzvT6AjdFBw1AHLq9lkOYONY181x9btnnj6h2A1
FT7W9ccaKlRHF4sjlNg9fILlKiZk/NIftG00pXZkidZuPlMTBlCz/CZt+7ZuUg/A
jrqOyOO198cVuHw2BZAlnW6ZcPOog5QW5AlayOfnOqx7GSvKd2QOHVTcfoi2lcq1
/w49B4Iy8NChdoSQBFVNtvoYroHFf7XU0DJOnwjk3bFW50PKM7YSBtMZwNi+oNNh
HtHGxnTHlcezDd5gcJFZhpXCLy8B1K72ZKZN9uIvFH4fQBDh2mY+f/SJRnHsJ0pM
u8KOA+pexGdUTh1tIIcug/e1vwlmVg0cO2KxHdsUSGpvmJfJehQl0lzlv5vy3QY9
yVyUb8ZhpNKwnbHsawtS6Dt7zRo0BGX0TKfSPjNKlV7n3tH39RWbXhd4or7ltgT6
cwAqP9rIMZhnvkIjzf4Frtr1I1F9KHQMa2VTaJin5VG6KMqgapSq33kiUJTlstA2
m5TQ7JNJSRDfg9iZ/8KFO27r8XC7oXBQcrrDQpiVN+yFeA7lb+ay68ZlzPZiK3AS
J4yRQdp9dIR4k88K5TlNDqXPvDt/WwovCmtMI2SsWN1dEaLHJB2L+f/j6e0hnGX6
j54vZQnMqtjVBNhwx5JhjGmByUrDVGEe9cmpEq3A1cTRow10Yupze6ZDKmnnv4gk
z/5p969pzcgpNPT6pV99kQVNyLJWOr4OLEjULwAQ+w/wLjmkiRtSnws6sF5eHZuD
SOXFRcJ+AxwcgRg9U3UWPGxucgWVxbPSP4XK2bEXFGXYjQ8kRYxy1fJpfKBjfWc9
1Zax9iKridURl2k2FuCPTtEYxsWlT/k6PlygzsiQSimXVv0ai8kofZCB0E+Vo+Iq
q26npvEH2mUj7T0i7MPSkkni7Y/CdZTzdjmB8OKcokTa9Rnr1hXdnCJM6YzB2Rp9
ltQ3H2C2aDwx2yuzlt/GEkxaU/cJzC852yPd4Zvx9sE8CmVdc97oh7FqjaWntp7T
k4cY1QCgasNjT0KdOlTqMfee2ijLRXGl1BNTHn7YkgCPiY198TpYWzl2peNXfmqf
YkAMEiZaNMdQD+PoFlyd70pC7yC7esSUHX8H5bbX4wRvMLEW9OEFVAUKtzzmqING
BCxaSJwn5biWGlebYz4+Q9ddi1bzdiGqTLhZY9zy+EEDsaPD0yXznUD+LZ/mY2hZ
pN27kC4rAe1/gM82BjQi8fJxcqoHcuQbYnWx03/sNASKpnbdRSXgCKp+D+b+Mxc1
7HXzTUJ8uA4Qh5Y3FMETjvhNlob+hJDruNmRqDd0RbClo8+LfOLjHBHQHFtH48bF
v3DLo+XGadRr1gf6fOA46Nu2zhqgpp9uN32TSZs2qqZCvFG3deH5aqJro1wBuNaQ
ruWL/7n49Tk1iK8KCumHMkmKPXEvMhm+mC6spH3ISztkzLT76SKj1+gd2aE1iKdp
gxkNZnPbl/Bqe3RW8bfPqObiLrsBZ2IsoXGT08f6/cP5XJMXrEp6RKOTUV2YK26Q
h9ffVeIJKj40tRLbj0wobmQUONoGZSslIRFG0qXHumwpfm0lack1mCVyFYt+eGVb
swHE4QuZFXtIsWEwpEfcO7Nmt04tjT0WqI30luD/gfaSBVC5Z4YshjeT70G9KxIy
wnsGMB177Xwydj8Syjd86eOW7UFe0ickHEtWbMkhRFm0QGSnmKln08LzzQCNabK6
5S0pXIDvg2nY0Urms2nTdSyLPR4CW2aUVKUXbf6jksv6uLwtGk5B/NZKce4odIA8
EYMK/VcaeRYHy0IrYvY9Ajjij+yjh3DMFvmswaNCP0YbW1CzE+yDKVHon/TiHjM9
65Al11SmyOSe2n5L7ahQXOYVL66oRNFqixWheNFm8QnAnkEdLhb6FZpZ2Q1y9PRw
hzOFVxWhXwbkULQYkCMMgNHw7ctKlkUw75m05WTKpp85YDswlnlWL65yg1WNRw4d
MzXIgvqyp14XsgGbGQ9sZR2NMkW+o8BoWuTS4aqXpjV/Sz/kzaRLaFiD3ZU/WrcR
/3Ntc7f9hI0q/UuD/eXpN6RF68YK24oHdYUun09Xy7pxRLlABZI2O7X+PYBIsET/
bT5TxytKGQ0YffofZ+pYiKEzmoPlisQxLxsdFzjHomJflz8kVeP1Zq+989wPCi8Y
p1NsUG0qeu+lXgFll8dP09TGdfZpb+B6+W+ykDSRKZfxJuuoIYlIubZLrRNwX14k
850qJbd+L79b7QrqUqrr6ZK0zisUqF/JLCR3p15BnjK7L9aPVg3hJ3aJZj2KBKaU
OIlnqFQOcSXZ9o72/WEF/io0cF+/rGYSzDudYOvAB7gcYZi9UGIB9GLB64Untu3Q
uEbOvZ9lVl6Bs+cMIi2FnUJk31Y4p7oNDE4aui6pTepLWVJuaQGnU0MwZza+RHQg
WkYLJRwu5ALGnv2wfWMnSTqRA59NPhCuXv8hUHDltK6m4iXMuRxiGjqMK7SdQYLH
DSfNrEZEHlB6tHSjHOtf2RwhKvSGcaEVzL0C6KHfTcweCwXa2nD+wuCyfI4/lQ+2
FQWLmJnSa7lc8WehO/5xXc/ZNUuva4FsSXSlSEmLgOUiznDqE19cxX4Ulb55fxuh
SWd5AORPiR8o+O6qsduzWH4rxRx3S7xDgVR6DpDl0xcjrk4VyJWSpeJ+/abJcBMy
nc2iKg+Zg/ZGkoxVROlnjoqXDBP3STYDPUlkGf49YppPgMZ05JGJW/2y4xsDOhtH
GVBO/nlRsxxBABdbi4FD3Q/U5TRsn9WGSmwi+kN2UqGwE9BWvHSYJ/0a2/yQ93CL
X9VGIs3vFOZ8fUWtNFXt6a/PIB6VqRj/d1b7XEByERViyYw7r1k2egFjAYuIjGf8
/uxCy7yYbuFSk8k0mgdGpdUwKnTpZhfKvTc05eZct/rDjCoj1PeP40akK5wsNQhC
UP48O7Ce+p1T3v4yFG1nfHmp8mt140NULEk5EdusU3xN2XzAx3tRGjHh/XfTTeME
QXMyQK8HlEI+cXHjo51etQSAelBVkcWjsZqxo3oLWryzh1wHXsPh2T48/TQQQ13k
buf81yzPsP7oSHOrx8bVk/al1/DAXJb0YKzuWWOB3UXcav7Nym4dgVteIFqEWfo/
KY917TqwjZAZBI1h4HwFKlq4Vfetp5Is/r/Btq2sCH0VXL3oyTcKQJcPI9BKoYjj
DuFY2HH98ZRGtslB9WrDjK4ZyazvhqzVmbIQvt3owrN6c+Be4k5EuVjno05dpOAi
w/eYH5I6slITQxnZdcnqodSSfWymEIlICxy9w2f0kSmXdRmuM0sMWgFioM9BbBt8
pndTP668hOoL0IRaARLLiDtRvLETgUNPrk5U1keJyUIHPH/iI+qyXdF5dfv4mcT8
YPRAB26DXRfQnNyCORp/ceavTktyryjCuC1RiOmv1DX97ydFjAQmHZfcfDNw3PxO
uJZNa2DvdvXdWHmCpRMlilLDIVtFyyNY15GY8TzZ5hqUiwI1Pyz21ypxwzvyZvc7
erN76nK8JmbP1jLTdan+0T0dHi6tZ7MXxc/7IEmm/h1G+YBiTzB3Om7+BXUoqEEp
K8C4LyW3qWpr/EQke2GzNCRllgHESovEwGj/74KvmyaatncIr/tWAsb24joMwFfW
l9Ti0NuiZ83iGaIWA/Du1VTama3zs5Asgf+ebAqmyklVuyHi8OAj/+WUCy6BZhR7
LTglvoJjcwt9JlprnpIcyqhaKxM5gNJH/kIusKMtFTDPbwPlQDJf1+mY5iTzm+gw
D+QQepY/NVjGRq4zed5btWxyCTqu5IFD6oMH/Cuza2saOi8Q9umNl1hMpkjs2rUG
Yc3V65aQUE9//WKBKCcOYwM/4aQIX5WJZvfMiEg3v7juV81P6sQODi4n5iSKk0wv
PsDI5wauo1n2xy6SoeHAUhUE7OO9YU3zzQfL26LFzH8Q8Y/7fCpCkxrdCfkxZ4KU
yax7T3nr56qjTMnlLYm5ToJRHRVNCc3aAWiM/Kktoz51M2vDrnhppfA8K5I0yL2o
ncjOCjfgn1PFOmK9cKU9fQ5PxxRqeY1e8sZ47P8W2xVLWJl5q56/6pSiSSYvPJdZ
IzYAnTgvtWKbM3/n4PCM/i8Jtn6L1X2AFXDNUfpmZ4P6I2j9AWOkkbCYHrWByvlG
KV6OteQ5XvhLthA+I6YZbvySVXkDUAMWsSTpRfISWhol+UIb/4UR9Jt4B9fyacAX
UJ4gLJI4M6UpXlNiIulnDRS/+Ivzyx0+XNNWfSyrsr7eUwqirrrOa7e8DIAaVkVw
MqZi/8QyGMVy4eGRyPk9ayIpKRF83uuegcvDDVEr3fc3Z3uk8Z3AFEfPNePIEWzD
wBHV3gyfWiv1Asay1977IomxH5VdjVnuv2m3Ahwmn6v9g4lOMIgCnwCOoxExAKrz
4D5n6DPiwScketo+8bmdaqXg4FsFR8iGxO7hMAyvBqEPbL+g6iUpzozJ6RWH1mVz
Tsc/I9PSQkgh/RrSm0l4kaOl581pQ1uwg6XANG+5wgkdBlpXPzUaGnvvSKO5Axlv
nzY4WTaaNiwzhtZwqXiYX44LxzPoUDg4/QVcBUKXAQJOrDwDnP0Cdp5ahfShofWY
bPfQ6Ty8zfo98c/LtKGqMBtXsowmgy/hABLREbE+r2MDXyuAUHl9XZumS1YcBwYr
xS1vcWY7WrqAPo1k3FMsWTmOZhICwNd/IKz5OaDzkywZpEtIsR2RWX+B3Wlf2Rqb
qHIZSTBoBV44eBSXGfHvLJhtKUgrUoYmn5SzRLVgn/H33QICz9IuwCHBkPh68EOi
AM2B67/tUrVei7NTosy/s9zCB8CxRLC7OmmV1SQOYPX0SBvTmsjOunPBXQ601bWh
oaM97eZZm4vTxNKRccMixDDvzkCOh1OwPUGaJqPLY+SbiK0z7DZp/JQCLJqiPcfB
W3xS+t/GEDCkGhfhidbcpgx+DZoEnLQZSSGdwzz9p5quJHVqYRkBVe6KWxWkSEDt
t9lsnzCuAGRHyh0J1kTFL2kre7w+c3MBDKeMVxpmK0PP/laRi1lAVzsht6wxyhY6
F3TmY5FIN9giUODa2p9u/yooDiWzLJ4QLbFX7DiTOjZWB75g+bAB7Le+mgrJ7PiG
76fdHrYzxeTLA9G6cwsu5qU8YAL00WR9BLj+U6FhVsbEbDHNJlJm/Xf/Pxe+TgKT
tz8eDIb0EyP3wvKpePh2TeZkcV8Lvg8upvG2w8W+NdFDsK+nNHpx/J8nZITs4gXj
+yWl2s8BhKANlW6xjgE/mBHtjGlsKYJrd66WeQOvFAbQ4f8pdk9mKZDyedq7gfNc
smacrZxL07Mvq+o26rqFKRU0AuJXuvDRJG36Bdra1euv9bzhTIN4HzQbjtAdUTOU
LiMUPpy5j5/vDw6daYjCHFQ5D3mVbhVEuPA1nQgSOi+oy/oH1vqNZYXCLAKTrxlw
oFjGnegAmfS89/0RJNqpa1wZFpjRytL0gEmUQ7eJGx3ewxDz+9jTEnrj7XY+CgOs
2Ozlq6iq11Ko87z46yuhamKMOzLrsXxEtSuK02KEWEEv7uOp1XWPhCkPwdvxNjVj
sM9ZKx3SvWgPYQHxZv2kmZ+l8t4n2wRJhRyaiWgPsQ/vehyqsadbmbe7pV1+JVJy
FB7QIDUZHwKmzVtyorPBsWoSqxQcSDIoA6Kha01GotZ+cB+LxfkvNCTgQEkB2yyT
sEfZuKSvWvFN5OQgWRP3wxy5J/UUtEuKRE6QeZPfGr0u2z+3yZ2rrNXyesvcoZGp
z7s35taGPR0wThtiqrItE/S1dJBhbH1jJEX8Hq8Aib2g2sgXfVz6M/W74SV0VLd/
sjCzbcKGEHpYFcfm4wF3zMlimdHEOwNr2mkhMvU3SJs4dOgfVHqsGPsvvcDSWP9h
ErZXQNtpP+1B6sr+HFRTPp7++7Z/wsF3pw58I2OtieR0YV2u6+ktjF5O2VGphEnv
Rkvmx2GH82p9wo71VnJgAoPweRTIaFhBhMWrVrzLqQY8tvs24aPRvFAcT7pvXxtb
kjlybQisl3qmEceperDDjuWAsS9QcRQ9Rrz4dNanCAALEgFrvPoacCgHOT5IePIb
xmtkfWZg3jpAk+iu1prWLX5MvtrgY1eamzFsmGrQJrlKfvTskA/8UFE9cHiYADpF
1p3VNISkVcOFQw13D6neY3+mE8Ds3jEDvYukBNVCtjENanx25FnMnNVA/4zXiUGa
k62bsVSo8MGepGYpMZcJAsVxQXdTRvQgbj1FZrGdldsDCI5MvR6kaambnXdiR+FQ
F5kbNaxtDUUNOnWFAFBfOLNDU96OfMOHaxSpQBwE7Jnblsrzq6HOu3LJSQlMrG7p
6xCPQ6BDtZvXSaqadkmsOGdGHdMmzlg4hRfbdeaX2usztKxC5gE0GT4v2i4E2knj
Od8uJVgLDqQj7vi9wYRGlGZd83MF/AELd8hHbCmhKmSu3HVV4l3jTJ/Sk9J22zzb
DVUokluO4h5nBC6XDWfJrlMimin7zYmGI4CObTxl8VBQ/aqRJrQD4lSW44LIsBre
PgJ6snD7l8CHw93RYgsc1cXTnRHRWKFOo+89yGbm9lEb/Q5185unkym08icLEtqK
hP1hhMgXfAhApo6ljWZmecPDLnxLUzhhZcwt1et403FpWwt2MWUA5o5uuQ918uWh
CxKsgLHJ4/tNEynvpL+0nXWdCB6odzCi5cy5UeEAgSI8IyWLCfQafmcA9K9HBWZV
Xe/aDsOFQB3/yAeD8u2mG75SxjEC6nC1N2PFOLuyaqe1R5u+0rfLsjMN1NFpsHt5
EfK5R5ffZBxzdZP+gdSpCLlgsvSx3SvzxpEGkRlkR58CPquIfkxcCEmvmTcqcos9
L1g0EJycnIfBG1uR5q8YT1CpRGiIQqhuB4Y/eDIl7WIc93ptqXuIC/iLUjaSzTFr
60fN2WiQnNoToJrZt6VssZtHr+1u2t1kpgkH+l0niQwnMHlHF3G0m6KDyzzfb0lA
nUYFU+/ljVNZXbDU2jrSn9G2RxyZtIBkkxGnyXR6c2Z5TY2uXfHa7cbOpu7a2+9M
PcZGtt7xZA7NlA9Pskdos9VHb/N6x/+giIEgEbH06woUCUSM2MH3xeRAEUM2NzLK
01maNGbqAzywwX7tBmNE3CWDb2gacQD+DYHONQ4GkNRcAUgboJxMqqwJ5svttuy0
M4QTZLZc7KmtHF6Wb3wcHP08HPv9Eu7NLDFq/oLEGcj6A5wne1E1UM9TYKp6k6aE
KyLD8kGyYijLEQNX9j0CUeHFSefx2jDeFpGKjfvjOWH6S04XW7Y3OtJTrUYpP6yu
K/kzzEx3KoxdZKXjz9wandHhOP9lDfBD1Mhls2mkaMRx+Fz7ojX9GBtGFSvLzebh
y4Ltk2EwE0P+985mzkR/34SAdmYQzoC7P+4HBNyfcUmMsiXLaW/vQRD8FYD5LQ+/
KqEZz6nTAEpkt+0EFX7uor/KJA1DieCR/wDMFN/4qWr9y2wxTWC3nuib8WhdITE7
3G2tjW5VpPX8UDgcn7+rmfYXD77zHIV/J3oWMOXgUIekjPmSZbcfYow2k/4JCqL1
0lHNJ6h8t3ypP/Jy1nH78h9/5e1yWkIkJFioOVWITr2pxdJ/tQpQmsbyv5ZEFNV5
iVKUPPEQpt+h9Bftkx5Tj7HUSCub+B9XD5GWJT503K+d60tkqYZET3A9A9/iIoAf
ipPVVVho8yUYd8CL+1CuWMC4liZKc/Gre8gO/0XU3OhiNwPIPFOk5fKD4ALytSMp
YJjICZhnU77IqrMCNOpA+T//IVB91lBA1Bv+y5PTbyxhWlwUprXHAB17xztjq/hS
JwsxKqoyPLLkFgcGTLnwCIH1ayMgNyFWnjVbkLFytD57O+eA7hc5j3nsYZtoctVY
WQpIyLB/YAdX2ExkMmTJNh2HpdWBmjZpnEev2hYSFGwfA/E/w+S4JXeRvBRIDHU0
1FXSIULxAXGKvvjjCoLSxjwt1MQIiqC2h8Q4tT029BoiEH1S6PtTpCeS0PHiUbDT
KtnQv92LzzW8fyFVbZtrlnH1UiCKcRqIwWfYHLX0gS6/8u4JNN2z9sVrK7SN2+Mq
S4m3TcopZQnsI5qoEMpxaYX5nOKx1Uec5JV4Y9vlG2bW8BAlF1waLZDMajqZRjVD
LikeM1vhuJUTph25LlPgmSUmslQGnLCcF0sUiunhNdb+eq0FhjgCXXxLXGvbD28D
hZMhDqi96mtYnnOT1VUY1rRROXZVPPLopxtWTkQoHpqlW/g2J0q2ClXKlrUJLuAS
LsKtmJqfnMGlgdFo+GiM5odWiVK0DlPkoDb6GfG629ivMwchFx1BCcRNmC1YWHNL
AjUggwvTbYQTNWHfRjf1WVxQSnn3Br/ylwe5rrY0OaUkJzDPRMiLhn+CSk0DOpAn
0Ku/W3amJROnFk5wPQ3GcPBVQlRhJDhpj+L7M1GHr/TiHj1mDsZKciupEh4E1kTB
/vxwqstIFzwQhJ/QxVvprRAgGFufU+pb33YFu5K6Pdl7uYmrW5e5fV39byRRAS59
bD6JQUYanxf99ChsmiLBXSS7hTLkIOEy4bTndDoYp5yxw9/0jTDZHr/nws+b4P8M
1sMU40+kLvD5kE07ZFQYow5mYNd8kwuCuUMu63eYv93OYLX6sJdR351CURcfyRcp
etVqLGY/CaoBZMIjbIYpXGsQXbj7co8tXt66/aTkd/QVLtuBKeBan+ip7hn2xGjY
7O8R88X4xOc7/TdYU/qQy3LhQ5X4McJ5C4cgXJyFN1QcJaWwfZmbA2pFAxu0a8K5
SZe9RbdjAY2hwQICz6kXGmkltGi8bwiftI2NCDiBJoiycqtCYCaxI3lTp9hfiA9C
9X9kVSBmaYmciR6/memv5gCcPvTfCXJ9pbvJdLfe28/xzI/aM0SJg+1DkjBaNqfC
wTT/OjbIhxEa29VP6TOwNm8CC9WW3RaQIDoexHBlUdsmTIVrsD0xz+FzbNK7yFf9
ExyHB9iYkdEWR1/kNW1jiKmLiHYqUrBjBNOBDD8AjA15Xt3OMQKmLOck/3ey41VL
3Io6lqDj4/Dm3SIhn8+tXpfr5jdKoqIZcp4rH7g8RTzAU3DAr52v1XQIO/4hfPP1
CJ67zJN/NtxOJ7IC8NhzQKdJaq2feG5M/UIRTFZGaOK3tfcjvWAWmN6/U3v+Ub3G
4dAHnWkc3KU4GtjpbvKTFj/xxdFw9OvfU/lB7gN7wq19qqjJD8cA7iSLSkUEXwh0
aHdwIl/d4f04yipUT4goPk0FbtBiyB2FuaqEiS4pnlOxyYYkhEhMq1hr5LRVa5cs
AogwDHkvUgISi9ywSP+3M06qPb/1F7JJblqCiBJLqWJRNQALedQfxCj/skcBGGJB
kl+IrgHHxiNaOGm1NDjWyy8OVUvL4sLN6egN6O1+oHVxGdnJrRz8+62mjKbZ2OGk
QNwWoBjQN0TBId81wJSnm86utXhj/t21b1EnH1HLOILxXnsNVmstzV+ch3JBgYXz
K/i5K29ir2GcHGv6FTVmWSnY+hzMDNxGdX/kl6jyDGSE9Ls4cb7ih0gHjGd4JuDI
s7Vyo+LFMRiXid1AodcQyU9JjN9B5KYRTZS0/8RnHRLF0Z42Q8pZGTS70qTiWrfF
5FYFgtLUuZEdk4XtM9XmBpo/QwlSZmzA5OZsxeimrCiXpNGMFlm6dkErM1aCHqbe
Dm1LDaYQUpy1JYHdpzRX2ZlpoQORwR2rWnYAZZIB6GK1Bzmz9q+ml8crOjh5/pyx
sNLhyptF4Ffn5qn1d2BeSZT1utdtqKqeHRhO/sU+3EEr+ozC5OWDGCfMzFi1w+2z
yYXSa82Tg3mV6MtBwxPiuRXHU4Ba3AzLGbtnxaOyEin67lZTriPWEBZXMw/IY4iT
lJ4DSAQaDIIW2hsRS5isnitXcW7JXdeIDyN8yY4NWPhe9n1AB7cF1ZkCRQg2sN4F
USU2cTTcFgNFNoMcSMD/10J0zI3XdKaZarkSAHrSHC930gQKqhzhn5tgJbZWuCeJ
icXKeR1syNlFtOMuuKaivRQuu4jLS6wCS41B7XSQhmhg27jNpQknOUIRdcD2WiW7
HD2MU8flbEztluOalhXaa2aoFtndWGIu+FVLxtJmArjR3RRTNygHULjdt3F3zRri
c1r8lmCOiVOMBF4MDLyLAJamJNRkmCTWR/lkgDdksftpSpni6KkwJqsENYmL2Msj
sdU3JgqBeZs3nPMtC1QLVIIfWt0a9QfLlHwcNrrBiXA8Z//hTrrd/6ge0aMnSneD
MvOCi40X6olO4xlirlA7DqG49jj321D36R34z3uUVX1Xt09KiNO3h0xWINBHBhW3
mMR7PJ/k9tZiNdyFsCxcup1ySZHQXke1OcBnA0S2m8vqRpkWFleSmVmzh7/sFOe+
BGLyCW32sJvXixVBS3sBLgp8ttSQnW7CFQUFzC6jcWNw5JxUGDifWb6H0JaDPcyK
6S+vdblXvwKglQd9PF/chmmjo0z6E+c3yiqylOIaX/fRDA4B1k2JklPD7dAy3Kk/
FwL3ohJ4atCloWWFbvrM97I36KAPszZW21J2QGnIfRqJYNZyR6o9gXg0XkOzv9bZ
Qeq4nc4rJi2lURj6HJWRG0iLZ2QzJbqrF1QdFhucrPE6cCH+qSvNFlNcROUauaT8
Dcm7/JWQRJcxFj33OVtNaoBk+yU0UvE94x0kfi7nrE5Mayywt0Z7eL/ra8NpVc/9
+TGhiLXJaTIefu8mIhcYmt0+tRwHtQTmqc/kluOqYYIFytJS7nx45ET/9Xsw+Dbk
BmYQMquVGbXKTUV2jYQ7u4k0kZxAxB1xfjGFzSp+JLzRBBWV8QoHLdDDrh1BoFP+
B7bbeChJoiCFTul63rQPDmkhM2CoNMHlOLWWTeR5ZXJUWWqmqxsATMiT4JdriYPn
h9445/3HjZralIkVb6AdoyVQIfMtQxXUxTow+tSRSwTqiaOsVulRwAvybgkCz2Jn
rcx8hbgjO7ik/wkBiQgdvLQfMjbFbqINtVzALtRb+8KSy3/5SXsmjM8OMkfjIiEL
/SCVN4KjekNRx3dVyDMcCb/wp+aVE4D8mUkHHjQMrJfaPwOLKpKqR/5FlAhfVl+E
OiTP29qjc2Z9/YNZYH5VZiW+M7IwReXh3XivNZ8qNSnExkEPceFLxdOiUiZBsS0O
YOUJzXnTenNkLHc7chl2oME7vO55sm8iK5mFFvVYmYL7rj1nKZmzTbnD8MwBnfVu
hP18D/DaEQdAnW+hA8GQTvjC+Z5ItYBu9AEvOJfQGxcshpdsgeTcpoJK2qaViyu/
ISqz3bGg6C8JlM5/6j8zAY3wMawVAjSgqtp7RBi5QAK5EwshjNDAQrSHldMnVFCY
kEWYKguCaOu6GUjzdywmO6/LwOeFVSP9LejDnY06fv/CaUafuRjXpEsX2F2mffd1
CanVVU04PdcQuPCkZygxOO+P1HUCPyNfFCxjoeUKn0X4WD1ciXO8C3zVVMSjHS8F
DJXjEnTIdJUv+pY7+r4+MgQ0yfXRgCkteWeavxR80MuLhnNxrw3HLg3EGj2PI9Xt
N6ptoPq25EFWV27dkHhZAXAK17bxw3YOZA8nqpqpJkZYCNp3OE+XjbdRbvW5mXFW
i7RSah0h2wTlWnu/E2LEYtXZRw7PqNbAZgIXuJbZ0/YsqPnh5pwrcCJB+NcNLSEv
/IW7p7Zs1c3KxSPW1YaOTbQbSCVIota0TW9L/ZOhU9cncIw/W6MHJt5f4p5SllHW
MsmimzmGwC/ucW+0w5gY2MXmQt42AquwWcBM3XfrIaVm3Y+3UrDDDkWDQlEdkoPn
pEDpVVuLOnIWOb8SEjkkgDFtolUZrObz16fU/s+uxMh4erNJTWDB9uYUacRNSt/O
oIMJya/9wE6dmljipy5G+Zqy4kJ0RaPzLgYDEMZUwDZT9X2GIpYKRMYlG5rA7Oll
/FLZ80tuw74i8hj3lQ7Dkwq3c77B0Z1oAj1D1gJcBqqiPr9z4gL68N04jA1ENoHj
ALnT8egQcsOjWoTYaY3G9rXCh8nZYRnRIsGEhcwM5l2HU67FUv70LQmvSGUgV/WQ
Cki75YXRCu1GzDtXADz8qRjPY8VABW/e09yr4jPLAPRdK9tMlgwE2XTl1jDlqho8
OnoOl18sGG34V3t/ORhIE56yWSOsdRid0P5RtZ2q+AMFTFjSvNG5Nl9ip6i0Bq66
LDB8KdER0NMQmAcFwNYDJkU2YSaQ+0i1j6li84M1kf03UW0/Pg2Uj3SnRK120RhY
ljfElJSPsnuYgKDdDHiJvdi7yDPkt81XzoJKjw50dI1zHbI5sMNQxOGuXF2tRcw9
fNZPorXiM7lqnwIKR7/Akz+0oYKkH4nva7NQPqXt2wqulC3VzNP8w/GYKJffctAv
aGlhiFUBt4CIZlKVfBYpiTre8jJRwSgQEdjz24ipBli84V5lRlixF+ujoT6Q/SjS
g8xHtDw2YOmCWyoBzXtw3AyUbs/TSevaDiRpxzYQqZm2bR/RYv0kR+8atewvek/y
5YCtiYsfjSd2rVlk9FdHdV/OVlashP2GjhT7QYSJ0U23vyAxhTBG3+yD/uPxLm3d
BYNVWcFHGvCKX7c3nitDdUhpt77P3NEyFngttPwJKQ26Fl8agL/ekLkiu128bD7f
GdKGJ4QIMFGtfqQ6kKOwEha8AtKrUDZ1wPPngT2UZOxRx3b69kD70Su7qAIDRoy7
CaLX/+Wzay0D/P6FCWiDdJKDbITCCbxrSSTN5hG70daz9qCWpWakgrVMjnbZR6Dz
TbqVO/h0ACZP0HM+EuhdcGKJnVD/pHDtfFG93fLzs2uuisqE0NZ1j8zIBHr3QS8Y
tMyEOHBgmKaldaIqkFVZI2TPofibruigezkXW6SVl9m136mySDJCkvyy9+m+X6mA
hWwO7B3p+mOOuUQK7bGN6JGuUa2TS5WFShAqk+smxxCapF9cal+ZBR40nWETXVGN
RG9IxYLGXV8OlIZsWYCRiKuEC+owCqC0iVw3Etg/8l+kzbqNQy/fOIbzwbDRK+Dn
u/TYMzALDl0h5YHPTu3GsyxFG7hch0uc+Fwn8u0uLLrAs966Jd00/EJbQ9flr9fj
FESm9fgn8Fgfha5g/ZK7Pz8cty1wrvFlJV9imMd1AboL3M1ee10/lWZNTld8Cktr
FIs8J64OmyhSqMnd0e3n3L5mQfPGvDd0/+GN6LlptwR/E2ffT0VUI48cEQ1zFUqI
jPBich6jOPCi2o5AP0eL67KxpFLyA31gwj612hGvD5CJG/i72HU721ICvb3r99x7
828hjSUUU/j2pM014jKv/GZMd1WGVU5mzw8h1k3ypvZZH7ENGOsAR07HYhGUSy32
`pragma protect end_protected
