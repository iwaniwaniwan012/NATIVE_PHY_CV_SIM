`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AECKSZ0HnFaVmAmvVLDsklJRyggyJ5t8N+4nOyTK20AtqgwmQRt54B+olkq67BA/
wcSk0z1iqgah/PEDSC6qdX1Aw9Wi3Ee15aDlk2y/G+vPnLpx+3QIiBDiDz/XOla7
cYn+fW+zB/chmD3KazMa5RNJ94GgaF8ZB0NDg5chnqY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11152)
yMEn/HnfKL18LTiYZjDZWxiqoVWX8zj8LajERs25eBWHZ35P7yhPQvcDU1AI0K7a
FRaAmqnFnhZsduyWB/lCHY8nIiJoOlMljpNqdzn1ScyXa+WnZGDPakGGeQpBIovF
iEg1oeTPOFSFPFj2Wnw5XRZcy3mCn2HKlhGvoW4CfFFu6hfPAO/26q6Jrw9SugLU
vpFdSSC6XnGnVFFy7F02pNcWURIZCWpR0cfFloYX3+7VipZYEWdH4UWh3D3xp8AW
f3/77Llcc9vB3cRDc/kY3+cn0bBQTyhhC9cdJABoM8n53IPZ7xdik2q6K7MVkUMb
a717HjGhIy0K6Yrud1acyNmXrainDwe/bzr7kSg07ZfC+F+uK36es0zv9HOBbevv
u6oyn+8Nr0KWtw42H8Y2G1S5up2B6Bq/Kx0P3LWETbmrIGuoDEISE7HdfGORYu4g
MtSdmGGtIuEYe6sv26QXutNrzqUtN0C2pzLYNfqgQxn2J994cBhZX4jXGDGzL5ey
zmExNsmfYpOVo51RXYQngTJnmE9kyTkhN3DhJc/bE9ok/EfVUQrCwgUvVdXsIJe5
EsazymeL3sd55zWosBMbiY/NufLgFPjfwyQIz2LZ1m2tBGVdkZtjmo5e5NSq0KH/
VXUApzB/ggfqOLLUkhDcTcNGjlMyacL8wqJht+1QhKFm9RQSkLq8iFyFR13WSEKl
3h+I+aZjEch/LkXJP0F8vTZIAzjA4JNZtVuzzEDFHxDp+fdnK+HcZVJZsgs2dUXD
RFNh5jrh2Uhi2BcwgAWuBdGFXMejQqwu8G6Oh4VnmwzEf7lSr+Szk2os8iZXEyGW
52VUxzR8Tr0QqPOwEMt+oFQrd0BkUVhuIL8zcMQIrW7uzTgUiDzH+R8EQ0vEIyYt
VtagqvZdtw71QFAqgtl8Ino5wB6ci59nW+AfijqTUMBsldX9JJbEzkbJzcEbf1sh
uCXB2HffpaYoUVbCKwW8OxIuJnNVECXqFhWEHeDs3bReTtVMKt6RWpO3LzEyNJ7N
XCC279xW8mpoKvZ6ADMgrm1qRnzcF5K3NDHsoPiPaWvuh2pY7LHpNyQ2cNNSBOt4
Bhczxh79IfVdgbkxRYttTwQkS6nA16j2lDJKrpCySzdAlQZyljp/+D3o2iO+2uE9
DggHjJt2XWnXSdIlj5ZZPlFtnHAv6OyC8t8W4YlWG03TXRDPIa4ngGFDPZRxH5kg
xPd8P08xTGyfEVSKOB0HpAdbMDJ+2U5On1sYhNz2wFX1H40+Rg4DuAT+ot9nOYqP
no5IqmBH8A2rl1+msg00e/IpwWtNJgdXXG7QmurMXmrxVfBuDU2hRrLDnKnpRSy1
Qcs/4uIhvIYq0G1jB8oYJEF2xpHnw9yZ7zEQ765QQ/uXP0EYnMM3XNFPIihuKEaF
qT6WHoQjkEDext30McYvWVQott35BhAHb6leordC+VXoaUVKetxGWai3QZxapVdY
17/B5GDiTNHv6TF1IZsWTlDE1hdTrJ19FfQw7dAeAQVUwjlfUsGyUmyj/rV2A+jb
JUhD4rZ+xWYz+C42vySBx9IrifcVTI/U1jiiGA7+Mi8IBymNh4CJKFIsPCNvEBka
JRTAxlbeBFvBFLNQeBZP0MKBZ616166me18qfkUXhZutIx3wbQCymljZ4IT/weVC
1XIj2N25ijAb1rl8MqqfuPwuV/OGnbfcAxrZLy7if6RwXE7++pJ65L5Qcp1TVlkt
5tJwU8XVOt9OAZFFInPmv1FmvIgtMSyKlWjHsEijtpDJqqzrAvWzAsmPv94STkII
5iphwnf0egiD/VYnKQN6E5vnSSJ7+FXOV1/BZThMtejRyc02bpu6QzzEgOD6jm/a
T5mE0Y02dkTKtd+V5aj9vcvjwkprSKzFBWAzvbPRbEkkiOcfWOP/MPR2jVA46A6+
bLQ4u9YfkeBtnNUiVLzySurqFZ1te4K/lOndkSYqVnympYIJnm/eUe+AuGxjMfu5
E73IcuaLbiHHdg7qT6dKj3yv2qe3FCkCwrQZHR7yqIWhbqABGCdW5EEXLMeDipuY
jAMiuuyDm5/374MQ/1CEFLZsZC4FxwrfEePhKAYskaBZKPToPVSOZkUVpLxN/jA7
FkFnjWHjo3JwwpYFqXD/x7AaMV6GjekypqJqKs6qQKDfO8KqrZeMcZw0EnUwdNmr
xk+I7Nu7uwwnTXDqbTNaxWwg4U516ydyPgbKau0tp+7fCw0hZ39PRdbxyehjHpRp
C2QsuA45hS0GONApgIncxNLBOxpLHU2AOlNIrsS9isobMZjqgxlzUy7iTCtTcCBt
5YERYga3rPtme2fxJRd1h9ri+w6k/fiuRG9qBRIpH4Uki4CBNYv9G3DcxcTvK6oh
XWSEwD0rNfD5eCKIjFSLZF9gaPmnrVVJaZkafveH1uLgywfWKJk/QeDLqcMn7WYq
bYn0rNW4Clyw3XewPblRBNoQD3wgsehNk0QIu7Xg3LxsX9HhnIXrmMMX5STZ5Cyw
55rxOwjwPL0Me4ilhC7FUL9ckqR2IkWGKePAMta52LPAi7+oy8mnEj1uTErvlORc
8BmJG7tFFdkZ4ez+jRf4UfoZoDEvuSp30kmladuS6wgg/Gt77wSAyEIaxnHI82mx
4DqrDDAq5D9YNNYl9xB69+j42SNlgcEHzu9tBaDJTLfJ66wxmv8UuTvLrRM8eXKY
QD2N3zvV4bgeQc4I3j8Fescue8vv9SMfKNPgi4Rwkg3m5sDdw1Zn+PAglSqn3Udd
UkSixBqwIzvQZ4RyJqQugDTvBHnzLpDf4zmh/KGZS4lcpyPvVMQ4FjiZyY6a7SK7
zkC0ibzTCJ/WxryGqaMCPIntIEqJ7pZ1pWoBlJoALK5Eix8J0vEO8svwQXOn7x9z
TruRNX9qBWRahgUZwDZNEDK0upqjlqLmG5XdbPvzGPFkllNpqmB79tmTjpLLpXuu
yse/9mQZhaGc+6FDx4SH7E6XWDEOEBqAui3ZETWenz0emgthkwsROsxPRPp7f49+
nHJnDs0QKxgb9NSypVy2JDSGPcQL681ojSZsuwRYUkJY8wewvPM1Ebd4uP9j6bEZ
GaQ9SeKXx6vqwvexdiazB4zpSuJClyw0yfTpKGAIIEA5YlJgc1+/AgHwr+GhX9n1
GQ+wwShUwwUtQq9C6Jcwy5eLWeIqKgW6v+1z+25kpAbLqidmjBvdb1i2xQ/ocbqX
WV/lSqO6IfG26Xhp8s2b3bAbrlDn81t8+KtHzWnBrmlf/Sjx15aNAfdPulYQ2bwh
w9XPn2+5fq9ryx3NsjbUAtPC+AeEMC/rts+5kFpA3TNzm0tQa9uf/XqWk/rJaHZQ
kqZIURuqBD4OjgffK1eDHxTDNDXazQhRjdnl1WnDn/sTQOdazz2nrSeksNhTnO8j
oZiFxHq4Wvqz5MpgVNKHPK6+CnsuAO4G/ZtxAciaZPMx3wD2l+Gf47MdZKVMko4Q
oFBRRz9AJjJGuFgdU7/yQyvMH/jjcEdxFk+KzdtdaFHRhE8JvILe43/JypHQ/io7
XwwyRC/wwJkZ5UcB7zQiiTirnryt/NuSD+sHkifruNUCefD9wAI91n9S1pYEv+AH
kaa5gg9G6SGBW4HFCDkngIgoZfGlRpwNczxgoaRPFotKYGQHoZOeGeEkODvA+Ixj
dmzvxMAJHdnYFSnZjF97ZEpbPufXVKIr4WT0XFO6KIzO2+xbSQinlkgyKCsrZXS4
oFkpMeekLPyWZdl6mZyZSi+88bmJq4Q0B0wvfcFYKKxOUuX76IRZmaiC4W/M5cOg
LgX1NiRI424KJq6VSTEwt3hkwCtJmizhawwSvS4I6KCtO+N0sGrCuZZHlnxnn1+B
ERGOzTSd9FAk5GZoKvZFXG9wxESNhqpg+RfizEMERBHnsm6Y1NEx1a6+I9iSd4QA
uPzC8FQ/rbc8yR3vCvrwDxPrDWGiudbv3BZpzkNXzMIOoK284htVjcSLYNzQxV37
wL2zgZSztRE5yQzAvDDUNeMU7Y4kViZyTgewm9zbZSrkquBUuITU6WuImH59ZqtE
AsapAMEQh1EFldC3LlK0qJxqfJSI8lNO+NbNwh7xdKECKO87e8qPEA57+VUHu+1v
soJqQm1FhOxvT4HdF4jzfLvnghCMNRqK0Q/3Zf4Rm2NgUeuD2PQnzyf2FNzTRnJ2
sGZL9uE4l6fKJFqHy317NFwyNuINqeqv5p1qG6CN6ygkzI6VRnHT3nmUBXI+f+Ox
7ytpAWq/zCNj8eHxMzJR5HxTjGj05o+/BbmIslgc50O6RcQGOIlJtHX1wlBkOtYO
7qWo7scdk9t4iHQYWP+FBeXogBa9yPPtmUhQhBTzAyBJAudgcRSCo+7jr3QoYc5o
EV2TTbvsmgb5eqQcWHbA9IwJgFRvO4RYh9W1f4VhzRHYgOtoWrHUC4Qn4HWZq0MY
IxgyNV5fGnhez9etG5hpoi2YBd6IwN5W+wu87sZ/EDMeO3S2Do78U39FOULEtYZJ
9sV98L1HdoaR/eKakP7rW8NcBPEyfH6JNNmn5SbNAMJywWUxWkium2htrRmk1rpx
6qzbNfmjaMTDibRAUz0Nqba3wFYj08xBfYzO0fJxIUYqE5HU8tjC6b7xwn3G2vmu
ReYK50C0IzBrbznAY8Kl28B6460TqXqPZoJtZOHZnJ9J+72d8Moq8C4JflUaOxI0
xC3MTqtZQIiNR0Ub52ezdafKT1gTx2HRLJRfw2KBSrlWjx633hjQ6Ph6m0Nl7iQ0
trT09ZIEaEvXbxaaWRWg2NXNe9BqTOfsKF8Ek5+ja25CXBsBXAjRi3WVE6ViiXWs
iI0phSe3Kc6xwLiKNM1NU+JW+ZYoxdnwdT9uOLPNhlzt58rZlBVVF8jDZNIlDB4o
cCVCtrn01NI23Y2vR7ZLNhB/PdKNVXLtGfH2LTnUoMS/YlUocL6/xvwppLMZLdD3
3o1tQmO14BbWvjT80MhWiQ6T/ScxSZtLXWdYrG7h5SX2e+3cN0tlcc0lKAtf6O1W
3fF3fa534vpMjRuPpimTmqza+GNfarc+WsW1dyelnGh/MaRok9tALk4kq5YOjBrb
D9Q05Vuy2bNSTUQrevWlJtJTQ0/MlCbjqQBhEXVOIZNRxI7RQIeSh9cEl4DdjDnV
NQMMWANQ6sava8hxeibSO39h3+zTbIQ+XA/Fhsfd5z1A9++xm60aUwKhU65vhtwA
LKmFnskYr7KlpEG26r+yqGjyfiBDX218kyU49vsbIclWdV8OEc75ee5zDMT9wV0L
/6n8bkH4fAQn554Xsbgy0Tzbo6Qnw74VYxEZqtVaS4Rx4DG3wPxs9FuU9j2beUsi
ICbckGw98aEDbnrNN8QR8t5+NH8ijFw8lv/ryRaOHalTU4w37aHpV1QgccqH/NTP
kK8wLcVuvA/2CCHIU4Ku0l+p/1i+sK4nT6nXDd6Jn0s/4UOdy+eTvl2+OeGr56Zt
4nLp640Eq9peG7VifLiezPbcYRMhtyUNaAjgeGsw3dkJ2Y+bYTtDFV5dOoWUKLOh
ewUsCiT2+T3dEADjtcsdt7wBQnmCFxgx0BZsaGMMx+xVcwF2LKbo0RZ1cEQuEoFA
P3hBesqTP6aUvc01vfRAfiSFiMpfq7xZ7YQFJS3bGdlC440dnLbgoUh7yuJiRAmB
B1wOiwnWDkviGXLscjLdjddxjNIiUk9pgKLbcqtT03kvnui2KyDWYC7UPuanzlJ7
iXr1/gbRLE27EseB6wT+pz7mwTowCBIeq83iw9l9R1evsh5ZGa24pxMakFREV8GF
W7vJz6rzTszMVBqHQYj4EiL64/T6IRoUq6D0juy2dXxGJGXGPLeicqJhCyJNZSK4
O89DhuKmN2H5w17pnih7kbeL/jEeA7h+pZ5RhBbWvdP60tY++yOV7jp1IMirgGcg
urgpjvHHerzx4TdWQgdsS6L1cODd4uG+BWey5cTg0fN29WIPJEu1wUi2Yd96hcQO
Zf3ye3i80qcmOgQcGSoOk8W5mGgC/eX6ZTkjzWxQtPrYPzyMW87/2JmmvOwy+llK
M9eoEMg6RTxdiYzsv/uG9buN/1nlpr2NRYhGZfwn5liX+xMhBwOjWq4hZiXKhD4x
NswNykXnz1PQoOZaKM8VssK6OnRhR8jlo5mBlP1l7NhHYpDfaJ/B3AucmQaVekvH
ikyhMjqj1kJy3eX8mhm1DYqSWFc9WQK/+5uYzVqpl6SO7+J5jaLm+N76a5ELvUeW
kXnWJWV/Bhmca7c99bcEU3+F2oP+D8QPYwNCs9VF9eynRwqrphaD0MBg/Pt8HEtu
HK9Ce365eol/Gn7c436hvcxGqIjV8xuWLgOrTSNICufbdgNgNBauOMomcUvz2bFO
Mu2leoipPuGCNbgnKnK4A2CZMTmoh2ZLGROps3uS0bxC0RCO/TSaunhhTIQkjcXu
Km4HAeGcj/8NKMt+03iY+VJkz0SFCEmpUjPmCgJyqWU+cL6XHZk2ObEs0KkA2n/i
+7BCfpM4wgVGOGm23wF0z5BzfJe6ZGj3hpzg0iBT/m3vg6MbZJqeFx4XzOTJ7fNS
NWsnKATSssK30VVYzB3H7DbTs/0DI1Z52FhGG+A17zSrPPFhuwvZ3oS39a8/2CRy
V9QBK8t86IWLKbiqmQqmiElaMi4PWXYCdlNDZrQsVI5837KVU19xayvpklgnnq/U
kpQIMB3Rh7KEewf0SGn50gHs8iHD0y0XO4WoZ0Y0a/zVYNv7QNY7siWX/1MZLRTD
Ga5DqAeV4+HGKyngq2PmHjHKwCtktKzgspBljaKCGG3bNl8NbheGuFcJG7hOtUxX
N5Qa87YHZoAuFPT7z/nFGHcmPb7D6L2Tm8EvsdI3/tNeJhP/AYRRODUVAKPIaOnN
lQYy9PdjF/Vpq7ZKsAQLZUM99j+Wim6Mb8ofkR3ouL19xIt6pZkT5pktwZ7/Bmpg
j71QnOHH+hvVexiu9XJrOodunmXvI+TooGNul1RF2yv2hMQWs+BHN0uJJHu+e6i4
UNhnUnWBUTkThUY9CD8e54z52ISF54zWBeZ30Vh96loV38w9DiGYavJbGhwIRXbC
J80k2mQw+DaWGMsLX6X1rv5F8vtzxSKIagPTR+1NHRpbMM1MKGrt2h1LzmhuR+4A
hUdSFitThJtH4VnoXgnkGFSxodjbBoiYgoAw/MqvVJKYObqWqvJXo9YJYDWY8VWd
ExNi8dhU4XMWD3mfY8TzZbI1Mm/T4bXuH8b8JnuQgylrqzfy30XejAXEvF1pmlWb
Rdb2fO68lxXPzDgwk+DmmYrtXzvkS7LgYu08zsgb/FAUuHdqm7Mk7L2kGjxHRlLG
LFv4GrUmHltEt2GDXvev/LgwrHWHB2NjLObUGmVa1cbrG8Ru9L6FlGGbXD+md9ze
eDetO9RqPQ59InWQkUOq/IzNtzds7F2mJKUQAdCRAR8m3LXqqjPVzOHvrlZA8KwO
xOBGp665lB6g1KCjw0TbgGtQvv0/wraClR8Ju8vZ9751njIf7W9MqJMbzmIqvxXF
Y9ppkJWHcZH7cpe/hnX5O9sazod2r8J4ROq4S1zF2ke7nqJnVruvI1kwo6u6+4A7
FwsDFzxtqgLGmWBSgWQQflRFZn693AowFYXMAwWFiUX+3XfdKL9XKHeY70yZm1Fy
0RLESYazDdsdOwXMUuZIkUwUgQwfRNvyWdH1fiyW2FKLGtWXGA6YjO7VGkcjmIjw
gmUQwUy71K5SQZcrH4GQsSP+cufbLVxTHgkiqMp4rIpc9Mt13myks33xaR56dwqq
xz1Q3Ty6Qenn1C2Ea7prEViP/mWLZu8Csj9f0DWyZKHeaPCZtPn2keJtUNT20nmO
qGq4uGWlmFvKx4/huwGFEk9p3YTuMyyMmaBjqhBXssCAb+3rx3ijlvAsmDSFSDkp
49x2hcetjqoo112W0qQ1E3YX+DDIuWq2d9UTWs3TfDRhC3ySs2B6dH3DOApVJUg2
iKUxkdBUpbkruq6cDljMcxeTfndULn65r/oz5iCY3BKLS6LZOvg8/MdV3U8qAt+z
p6dd15NT3Pcu3XOv35RDOVO7CkOqo+M2v07RPSzcZYa2AzhDaXPBICrNA4cvs8t/
WUmRaVeo5xJ6N8+KImIukjX0r4JjbdEoER2PNTZDH7nmNDTquJqSt9pEaZavkdZZ
0y7X80nJF0Tr1y6ChUe+rh1chhe4sOBAKxNQLer9CX3GhHGycl15VQKFTiEtF3a8
ByLDOcF8QB+X9ssL/eNoaNwwgHLuHfEdxhj/FhRJkb2fj7wbuTUQaUQuiN0HD88O
EwN1JA/FcOHiaW71Ze4cyt4c9oInVTjNvz6Sn7sNz+erRzQ/8YDKAmaNzK5CjgA3
+kN2w2aa4Z+JNa3A/RFydORczsmBpwJAo0Kn6Vz1vjJ3MUZXftLrIc2S7KYogvpo
rvDJxkTgbtaIbP4E+H+FB2jlm1y/CSvfrayHfzDVxd076CFNzTB3MtHchiov2qsC
2yhQG4oqAihwhV3gu76GSSOG8++H6VAqmcT4J7e/Sqb6Mbt74162jJ8jCgx3YdgO
CcdjSPGJLJG/hRo/5CD1MepR1Qf71N/mgU78+Mac7W8Vh/+lVzPyNUcHMxgbJw3U
sUDZQuwE3D7nWLEkGetM9UEmMQffUrSa+wnvOQNoq60YUzAJNeIW6U+ePHqrIQ3m
99KVr2+Vwb0+OI8lBZsX+KEro8vBXaVVXGlgqNZl/wnvecqZfSlyfLt5JwxvtO2G
x8snnAJDnmwch+4+271HwqWO/X3AT9H7PjGbRFxsEAq3zvvbOKdSmATHhuy7XQRa
MJMysKqhodwJB7czWsjgSYwuF091BnHrXg3ORcrn17hlVuDjMbTGY/+eHgWi3Fup
DGdfXNpGgC8gKB6HW+iga1FTlYpG+6k71R+JU6SHCC7yE8y4peZCTj5J0rLpvHoi
C2zBkX3J+EztW7WGem4bL9IkZNyaZMzFNBU5erDVMF8fndiiyhtJl8QchvJ6brZB
KUoaZQsYYMbArdM+b1n8aAeh0iUWCcscRTMH5SOJ1MTZs1eXdYgqIVbpOCyU5P2y
5df28CjiKkZXQY+WZWUdsKFFGjZ+sciztLXjxweO+nbo17LNXaRtgz9T5DxbrhEQ
RytWPrLoQBfC8PKXRPXzcpOgJTaBArh5fs2YTSw37x7IWifdDcesFnMgiAh/DtRt
VAhM81M4I+R/eoPhc2EWCckFKkCRlz2Rdg8Ty5xjP7n3w1vALBDT/yThKc79akrR
MH0f+gWq8togEzhojQ7P72NkXATgYO5DiAvIvwAk5ZAzTJ+pohbovssWotU65ox+
YL/CGd6CS4Ys49+4WVujI4A6vgsXQy//B9zkmVo/0CR6EyUTodS7LNGAe2M2A3Ml
oj77f+QbQursPSwXBct65fUma+AljCD++c+Hzv7rnXllkYmY3+SbvcG4CzizHcsW
5AMpi0rZl+37djK/qGBv4oYu+nZw3BtOzrBkVIKYCd+B7I4LOKNahl5WI9FjdGTN
D/iWPYbhw7/kUFzoLB1rUCVJbwgpIBGZTSJDoNs1r9P6E+MKYQAYFs3YZ/frDVV4
Ptinz0uACVD9FknASb/HB6J7V35KEcKMuUgPSjQzm9XZU+Pz6VgafJqUki+j6j1A
0fYBv6p4q9PT3JYFCoBNqhA8yoWX/D9i02e3RHfr5X1W5yRBEiWvgGxyOX0p0pW8
dcYgHbdkiQ5rRaOkNN8zeSsGrNlpWxMI11RN4uiNZb0OLlbRYknfdOG0rndxjz2O
YDryMGv58yDunL9dsDHPqXXx2wIzsppmglaZguNulRhPCyR6FCkyIf1/pcfYAMlA
rXJ7wqn2f8cFmrj3GRiV+RnCepmUeCMIxK8jpYCyr0J7zhQMyclib602WRRl6dRn
cHTgjIE1b1lOryQLKyw2l80rOk4CkL2O6lx2/wsQFEtnmRfeIMaSK21+1mcZ40xo
836mdq7mxWFZRoaPfN5/51S9rnDlCeRtZ33Ix33ktdGG/EdBNcRAk/cK6b/lYHcN
wI4qEsTHHclwod6gvvtC0xKH9uS6DWMpCdRbzl9qCMC11O2JTu6Q7MBa1a0glAFj
ZLT9a3HnAIsA0YciJ7I4hok/gUclnYS6pZ+rKqggX7fOy7Udv6Ld86XEV6UOntRp
DHt1XoBYiUo0yWXhx+l7Ze6iDk1WE0Xc3mqev+z/YNIcyynXOuWIoYuG4j6BYBSG
6jDsWk8fwlmAuvNyRjMMqFu7yACg5s2ApSextUdJXzWlZBYv1S5pdlDSJFwp8R7b
jMfwfJHvEJg78S08thSFPD9eEO8A7a+EFbVjv7B4cF6CsTOlMUiGSThghQAdlcdX
C6rNR+dL6qzOW3EvoxEzH4LRDZes8esmQMX6wrZOLTci3gl7RI/mUf0z99+hJ4iX
0PtRAGOScthHZRjinFiH51k0TApy7Q5CRQONCxmZQSqW9WdVMaY8IZKsGLpIZdPJ
TXXvHWsKeis1qMyF/qtTQ6FM8s6AiX/dX6EJJWzrDzxy+XRjl7UxX1d3vpT3WSl9
9LBJsrPY+sjoKfxbxj7p0lXqE8nAkEW4yMBoTORUVg8Et5Lxk5YqFn6cU8UmJh53
a2WlRa9FX8j239m5c0Vu9xH276UKBrIb/rfBBkP+CanqlVa18zqogHZetbfi/Aqp
plKddp7TfmtWL27RaiQjCHY7OzZED3PhYEcgDdpkBAm2KcBJ0cS+2QKW2F/4p7AX
bKsN4rKO3KqfdTH+Nls+DqvqHEUJthf2691umaukY7Ve1WWyVA5lAvFdjkdFPclE
Ht7iWRcJXfcU44Qge9UDjjLT25l9UxVDAWwNwnaExQSCd2I7gF7nQ3pp7+BJ+rN9
PeMNWMF4ZTTnOmc9fR+dzC/YgAfDnqaMro0SzghqeGZON06tL42VdDGSPlcys4Jr
lsWYRhWXvcZcxvvOfkFXY/gqY4/PA6w0Qs2dfhrugl/tkyY5NDn56bzCZQsGSp+C
xIgxXUEHpRkBBpvLqYWiVoXiVoWktC3mdmkUqBqDOzDisYO94LArjPMpveFoUbPi
diN3NwBTPIMxpIzvXDpfeNtP04n9EZ8RUQoYDZMzvea6Iyn+iCsCEU5JD4HLdmVd
QCfnXCYa7Ui8TSJ31MX1GvvD8DctlNXeLuB1gTVO2okTNAuKhvYxIeddpJ7mpP98
7lcyyPeqegnK7A3aVaIR25DWBGm/4sz5W9l1Z5mVtXfPkE/N9bRQjEqn/jX2/ciG
pfmEQ3B6Vk9mDi/4Tx3whEcUUBsAazJyns76YZ+/EKH6UP420g94cVTJlrXzGKtc
JKhfDxByghleD+my5oDbe/Gz8RmKf8SLzbSWRqyVfOaKgXw0qvsCMaYT+xE993wS
tE9vzID99UGtzt1SgmOWpM7ZDAn+pF2Hw1PAJZ8R6Uo2wEZTuD/pBkexDanw0WEu
JEWMhpV7CC3N7m+K9RWeF4N7n+++l7bi9nz/lL/Lv8Hf9TWZby1rxZM8a9qGY7mU
+mhqw4iTbAENcm00P5Eg0mYucllqHkw2+7KogMXgLoPspGUaWlIMl66acT+EA68n
XhmGB3GcPUB2zJTcxG4loZDoxRiV6pwHSXmgkfKPB1vLjO9ItR8pSM5p/YlCKqHa
anGfA6/JF6HUHgQj87B3DFCLr2fqRc853QSigmBnK/yM6ldnQ0xbDGvbJT13JeNq
oY/cwmw72VCqO5sKSnefRZa8xM8g9YC9fUo5Msv9nkiUP1Gpd84REHKrDN9swL7A
JD62k2enqy9ibHj+xzrD/r1BzempBcvF1Ss3KEqa+NCv8zD21c2wFisdT1z1oQ10
C0Wpyg3I2Lc2hDag28SccG/u9hJlpKdzyrHmEVRf/W1OfpVrLwubU95rAwR3Irjt
v4T5cLs/KovkzXVCfeEX/SwSM8QBagozP95dO0hEhMp159EurqOXBUK4qNGhP95f
ZunSwVlLB556CUASwn3jsjT9oLliq6zED4gDY7ehmyzlvNkx3I5XwtpXRkI+LYv/
yVyDa/Nw5FEnhfSstyU6ue3cp2b1nn4I+XVgeHCQFQAMN/TCKt4soScpyEhMhfsk
XValHs+aNifhLsBqjmGvLGJrZl59TiTOzGwToZjXQkHL535MuCxIrSmQaZr43C3o
6qA4D8imF8CWbWPAZwT4sAOOIEak15wrIq3ujmXGOvjLA2Gl5ZxQXsNUqW+30iaQ
6bIhNStUYEvJUmmQUVlaXUg+3ETaofmD4ApAiTQROvUf/WYhXPe5z48omdL8fO2h
CTtwcetbfNcU+hnrMxVl0tWB56XwUn4scqU8xDQR7NtE42mFU6U1F/afZBb1IO6b
sb3wxYxGAhuFY97A/kPPDrRZB/2Svm1OQ3rDtbZHgHKr4JBtpMC2dqwimlZ1C1Hv
/zGwO+GaXIDwvUPbmm/GrMWH6UwqndMxMuCYJPq/Rvs33DmtWrjQRz3MAoCxcgP1
H+DXqe/cyz+rZbCL/RHLtVJ06zAi1IXt2zCxjbKuJT5b9p5deWDAQ8bhdx/W6vHJ
yTEXQCvtZXZLp+azJnkrVStYfbO2yi0HGgCzt6/fXElTspKKqz9MnoOvoF/xym/4
7igw54TYsCL/kA9Yha63ISTvvlv+7VI8MGD/yofdTRgkeOX59uU7ZKc8FUwRCRsD
4ZjH/Xc14+Mc1SYxwtQv0HeWKtuTfIxHcEUwcAYI2eF0foNmCsfrVdfb0ZpH34QM
QjFkM7evebiUQV1Je257vEJ/Jz2RXtu2aoZ2v0KzXrlhY7D2CxlNBeZdppb0LEAd
C3owSA127vaSwrRutondDqBH1vifUIdPEtUOwmYO7Uy7eF594E6WA5lPtCeoc/J5
k/tVKnWlb1OwPDae5ZUyKaz7pTHd8UgTmOajgjx/3YfCzMga62Z22XAxfjJ2UTvG
5r+hn1Qp628GbMGaunCiQODYW2/R+MGuvML8Dkm6ULrIc6I/6UtlJoJr6QqSjENR
7igxAGg3wa1Com6iTURaE0mQBg72aZLcnhmaI2JGABpD9ZSDYn3l6D8uBTRwQAip
X0b2/olStmFC5VyZ6/sCRmsL5S0bAG8vbVopcFWw7YTeSXf4zJRXkmj9+xt/R9ET
ugSl7zt4cftIPxuHQrP1DlbRyEazanODzOnYtAC9z7PaGVbooj3mQDwBGkYhre2z
IGb4ZU/0hUo2C90QJpQL4jKyatNIjOtXsABUfTQyi1bc52faKegsqdhClRAVCfEP
ZpOJrJlzu8v6n/Tx/AacYzQS5IFfIiwgoC2Q30yDUlU4ciKGK5Hfb+MM6ZZqMZ6B
1fJqNdpiXILccCnSTxJv6HBz1O3p8ECXeb6IhFkDbga/CkwgC1pObVGJmecmjmRe
jn1uAzttr8yBBFq4Wu08J9+ONHvvPm02DpOzWbVPrkkyTu0R5oDbepH7PR4JUS5r
nX2N/WoOlsN/Ksu1rwqJKyWJGnCMjkMsYN9LI1QTaFEA4NGpatJuyHAQ4iuR2LBh
66NVy8DzyOBtDKY/xgE7vRZVXJbFcvOOGEWGwipC3c5QYhGGVDbH+dsMvFL1xHoh
uNJTpjKBh2ck/yqTzDFGrBZoBZnVBhogmI2GfRcQh2bHLn3zUF1kiIpQsJyf465V
pKTj9h9uyh3N8NehKdZrF19XGU2wYZ4vQ8TtaWzoe54eb8jLDsemzXFCrAdoGVKA
kAgci1t1IzUn+YXeNPuV3fI2NMr+frRFk+aXoijQ9L2OlV9HsLZgIPN3vQN5Vxu8
JnIUJl3oMQyGGSpxDGD3CG77f8CJLqBn5c46r6o2sA6a11kLW3THIDK+8j9HmSMg
phmrDK4JLk4+R0k/qzTJQhDgWZFQni2X10ow9HqgaIzUkZn+BalCKJROYNcSG4tF
NT6suvHDTEv6HVC6sZxQsEd7bAnydM1XPiaMJ8GKJqDpDQXaJ8XtDOg3kZTN6yF9
5UdXrArtTC00Bl/D1c1+eOvB6HWKPFhx9e+ZVBrL0JhjmyiUornpLRyj5iKtspqs
fRNH06V+8r49t7Kiho0EmuinRXsv0RLpt95pNpZkm60BllnEQxXa+laMEdSd1kUq
Rm4qE7aoBOwXBOSr+u7OjClJpWvvzyjqjJOCjwZcwXjC1VKQCUa/hgcCvNBKjQ+5
fLxbIfXPSChP5TJK7ruAfW1OSUVqT2O8leC8N4DTerfYmZxYHa+AHE95UbDw3QeH
6EXeGaP0bxZR9iiX1XndFurG74RR9CcYgckBY/SVataPpdw+si3wc4KRccNd7I+/
y4SZfeUt8uofndCjGBiv2xMHrTMFBg1PAbaABvIyigD7xrJI99Ont8ci/GV+3Wts
E1BahEw1SkzUVoppb0bbVzuTs8AII4CWaSyaoPitwMBTrcMWqyyudvVrzYh8Cchz
5XYoDiScX+GJp4qauS3ux4sVjyie2vzEiuQSUAgCixJLVBGpNKqy3CLp+K28SHSl
x4vQgZ7rvFHZyKLpLUWN2fDa5/ABc2UDabEG3btw981Ymooi+YxbR57/Tfy8c0eh
TfELYVfs0FCMVJ0LBOQ9VwidOspoDRtgWAybxClFmehcyHhV8JLkiOQioGZ16H3o
CqtN9yb04O2bas/nohDr223n7a4u3rVPsAzw2OM5NxFXSJFSRR+i+hnz+hZEdNmc
o+DHMFifDCQ8n0F/J6jPicZczhK8cG4xRJcdrq5ogWjEN5Dzc/eiX8ghICx3SuDv
AQFZSxluK7lHZPE1jKR/2oxNcjHm5DUiSYYXp1e1CHdl75BziDTASs11AaJiAxs8
4O5AM3Dn5D3LA+Ng/cpsW2PvKgW6pl4QAZDa+0PhFUHNAb1pjK/HIaLtDy0xWHP+
Y/NuycfpdJj9OunxkloVcIsSDaIFN9fNqNUUjr7i3PSZmNS8ZODxGxPxCJEcNhLa
fhucyX1l76v0vCYq9EAQrA==
`pragma protect end_protected
