`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AIMj5fHH9N4MTtqwjwO5CxnWBoMwHThIaiUY++21bcz0k/hIHtsoJalZiMXx3DfG
9F2/u1GAGmC6ax1e8Vi9LhUdfWszr3wtiJpulIRaA2QtQuXlfoVlcI/KZRqkwBjO
JQESi/0C1INtjSDwmPfze5Joz/2CRErzLWA+comG26s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5648)
OhdD4HpRBxL3M5Jeo6+gRL3lEUujMIkv5epLEX0nuOEVNWT2nFCpEvKqFsqLv9z5
BIa68kVTI/iFwZteP+Ka32kZTtFBwXEJv1O+E8Cft/7U9kPdee7U6UlUQXltqx+o
nyx4naBqHDtbeQXIkQYJfiqRy/SE/fGt3Tvsun4z2sXVkQOqTErlcrN27n0TgiYv
JilxQFybq7eNsLV7DFtjsyPgQJoB5bZD84gMA3cx38OVBj0JO2IyG/OkC+gmLLuY
Um2BB2iAip2FXbm5OzPhe3qsnopyPuWVTObeT/qpPxx8ZPB013ncc7K5zpdQuUeJ
02vDGW8ILyNB9s9u0tkauPP+e1l0aKh6zUiNwOLL4N8r6k3qi/IkICO7K5X4qit5
ATra2fv3p/FrXfL7fMrSkJs/MCe6m+HfAx00dx+rPORrACLV/0gg9V6jJWW2Gn7y
hif1c8t9D5WeKrfddyf8okTFiw/zTLKwtFahSkE7RgyITxdCkdx4cJEMocKApleq
x2VlV9XQMZQw9RCAWPr7ctDpWn1WiD+5fqrcO3KvfgTYCCPqTd6iJkUI3VXREU4j
nKPOEGetehLTN4bnY4CX0vugRlCwgMBnWd6JcKPTXwfSCVsBDxZm160pR5/wps6k
+U+lVPC4OLbABkuu5+iNYYEmARGV1wdSe7qyP3DKEP+/aPnV3UvDV9cqu8YcwDiO
lH6S9BlszNdzr8hqsFannumw6SMRrUE/WjIYwmMDA2FIkf0gEH+jBftNKBQ/EdOd
KE3eOmGejCECkKrHDEVt7XfDfcdnRHjV5USKyW8FYZlTklTbqCbxlIW14ilBZKoo
qLhL/guur99oSm37qGLvEZ/7B6MGpNEzF9cat53Ta1x7GgHR2I4EvlHjYeWrLCAG
XUh/CfAQgSYAb5bArcDsJMfy8K+vf8HoQRUjWNWicoPYb2PyDvkWAPkrR2+iw8Kk
q0002htdl3ghHiorsPMusW7yRJGJOSkO2dsDlj7mU70YAlRG6a3GPfPhX0+ktG2A
WxnYOZxpSMJWgbNHP6k14ao/XEnNcMLLclbgpGb+rkbajbgqMID2t8ER7WnOL2Jy
cFYZrAGDfhQ0+rmcLxPfw0bc49s3L1u/0ogCa29AnoW2v8SBlN/RLQSqnp2Fq2p0
LOeWbyihH4qXxysALTpRvx2Bk1vpmSPQUTg/7Ty67LWfDEznGlsRFIFN+TLI5XCY
8LVIA+5IUEZVtJlo3k6yyUGn07wGcGLX/mEwESziPHBkuxSIx7zwMyqHypA9x+CC
9jQDhAm040mjYzOWvLXWDRmIWBglOTslHbr8bI4X/PiepPwEtJtmPjYVZxE1UF6+
BucUhqyCgmiZG+P8lioKQkCyKi4PGngaPiPAC/AxbvSSdlxYCMI/wzYKO6mr0MjB
Q4TLjnJOLnxvuT9lqTbeOE4yqc97OC22Aqhvg2g7WdkNx6/IjvBz5UkqZ7uIaKpd
h1717it9PvSppIMpBIU1mmw0nyXHCXNTUYqJcB9D+Yrc5nP8YnHFS/2u9nryh9X0
7Te3nhpWuTBnVItZW9F96zGzUT89aCx5VmaNtjxlMbBxkyJsyHpeym0TP69wPsnM
wQ3hpQ/mUDRBOu3epSFAttUmZfwZ4mcWYG2E8T25waktBECfoeoukziCjUO3Jmng
MWAYShQLGVDDuu7CCKB4fcPWDVbWpHZpEPR6vATiJRloVniz7kZn5yVih4g8KCU6
L/8lm31TSI7wfIasEG8QZI174tbQAD61/mah2j1gVW30m1JMKnT6SrQEFF5E03KS
+wUqOeJa9TGVtGD2NsDiGm49QnlzkbxvJjlvCuTQIsQJfAPpcqz035WIH2yQTcV7
RbyiicZp2cyqw8Q8l1vW+Gv/PsRGY341F5C8uMGHbDCsxYrYtBYfcdOnVk9w8GOi
kHxau5LoKzu1/gDrF8TB772StO80kxdzzdbp/F7eg+cFWhzz5XNFemThWaCOxg/A
CFFEgrjuR/T43ygvFfEzdZ1K8FdgLrXZLuP8u8XG+r/DQqBoxOG+E3mUe1ytvKyX
5T4Dh+1Zkh4zG9ahVp4qWUU5uv5PnHT/FrrGFknjpumWpa1zfNmwHoiHM+J3eWHP
9+6E58qJ1nBtODIhZWEMsq08VpipRRP5fzUQzLSo/4X6mEz+zgm91qCcvgE3Zibh
mPxEkz79b0O8s0xbJA4w3N7Fg0kObiwL5JrUIEsq3leiQf2rt5Icyz0MiwJRABzN
FoeGj+WmCPrQxnhEGiu+jA1rpkh1f8nW+tblBCNbFqo4ysw2E15p24b53pewgmMb
xKL2GwIUI4lnAstwU7VXCOb2SmiPdzr6Y+uxia/blwv8f22P5H5EDpM/FiWkQ7ZR
9k2GEFg0emnDJh1eNBNd+fwoKDefwcHHPK23BmEB3lEejuIDOA9hrMrj5fA6/F1n
fkg3HfgUmaedyO8RbN18JPIwXXe3v20mCTjTe7oDEeqGah7DU5Tf08T6wTQgeskl
pgeJG6/4qd7gEdjwRs5kqRtkXPiOfZ90DFjUOWO66ylBMkJTwiWK0g5uBgeC2LiT
TthNwFFJoZx2FT8ENqebXXUW8/rBW2t7BFs+NRojJa7t5DxApknrg6ElNlRfUrSK
VO8xujHK80tyFe9M443nSQxUNAZSr56wxujEcm6TibKdmkRU8D874/EnwS33F1y9
/0PhVOQpkMBL0ibBJIng+jol16+mfPBLsWEAzr9o1HtZEx5jhrncWAhE1SdWrRke
JAfD1aS3Bq/hOA3uLPnOG6AUA37zxAIvmvzoqVD7eAiE2L2ZpGI42JmVIc/AORTw
zbekvgdVMEh/NoUr0KV4FCZCEjBuN0zgz06TND3mP6i5P6lcmsdUuAU0diOz0IOK
dxJQyW4oAu/g7ZqH4eBFQfLG4WRP6gwAuN/2xwBC0z5/JFOxz/+r9KdOfSC+2ZFR
NO3oY9GvOp8MYSocCw8/qjtU+W93inssqLh7Q4CnRPRFEX8NBOmYeNCAiGswhseo
agAdZodY6GIASG/rP1QUlJcDWSYXyeLmz4HQKAffRg4NbuDVGexrpaxPqviDrui4
bwghn1F1cFVCrqqRC4qEZ3whvj0iJHCH8YmD5OrKgDuQm5zxxpBtTtbR2DGG7IDL
2c7Rzx+OzrDZZFM75i9Sz96bP+zrcOvORh3mKE3pLbgnhxHjhgYsnT0yv9a3tRtA
gfRNgQf6ZbK5diab52VrVXzsH+ZSOtWIlStLlDQvtZoLOrxjIPtSjxtvkUlkt/yH
spOnoGmhXgqjc7vqRQjHu4P2mluNFUNEFkHduHznzITD74J+eqRR81p+tLeBeqre
4xHuWxckCnZ+JurgpZMgxwp0ZzGrUkUZGxR5JqQudP09prYKxpU5y+qPorPMzvm8
LqB5yLPXwiUnAgd/RBpw6Jaey+0z1LvNVqWF31aaJe8pWrRZwdie0lUdniltkSu5
3QDCxb3x2rYQKhStk6RqeWSf+t0Nn4Qqb1aVRPs2tUE3A23+TF7J1Xl3HXyXS01d
aTditP7dIzlOWaFozl4MdXS7YOChvXp72MxAOycBb+3sMYRn0EeaigW/6OTl/gCq
FWnYd4BkvdqJLFykR8OJVPrOItv6ntJgQMqL+zW/glel+WFtO2rcR7NwEgW4K5F/
dxVvp9cONnJIpxpWc61DqW3Vt4VadNrYf4IYLala0aZYNoCym2NIannh6ylnfjeb
Yv4eP5XG6QhMeHGUp7dXaaQWGLMCbuB4G6AE3muQ/dcD2vjiuTz4TD0/1s2yOHmf
8UPksZIA8Kca85o4kOXzy+F1UiGtTOx1UWd3XX9I2afljWmWb40hRansRcn+ryLB
z8RYjE25Pl2U0wBZXYbXIb2LZZRIPqpEHOtLJIjmTSnvB+iV0xrnViSP+FO/704V
LEEOlvJV9nKk+DxSxHkPgUSZ+x1Mh6Yi341w4N3lo6PBh9ZtgMP/Inuw5dhArIxp
RABzngxDnmz/ghHC19nQpdWc8XxgnlkKj39Wb/KXD+IlyV0nQi+yz7AMieGVH6Vr
BbsHJx3LJ4goaE3JV91qQknPzHAsUuOZNxmh0Dw5QpT4uNwUrAWv2Ab0V4O6bNjk
tT4TzEgfk8qqFZ46gCdhecMSfizsnBl56UfbHgizg2dN6rR9/nZ3cFrHkKcUxh9d
Ojjzck1SrPDvtfPQAiKAAORsyXOO6QQS/t9H9sxFXtYlXc2biV1Jg7OOziEhulci
kiskCS7wp/7q3M5Vos41bHsjGCPZczzVnOy4xwKkO4er0a3jZdMk18jH5yGzs0Y9
JpfAmO8r648ouytuN66Bw9/eLDIeE4bl99tX4zZG7C7rLRLlYlMIezGUfglRFqHA
G4W1DJb004+aqqX5bOMfn3KJBuEjeeyvIjCeKIXNC/FH07GXHnhDjuyXN5G9pD1x
75Gu28ySFwBeP2YmSWpNBoHP8qU+JfVxZgoomj+pm3V4fktZu4VEo/yNRe206E+M
XOyJnKAgsvDDg9I9pXN6R7sl0zkEymdQxBpzPRVIddecBgw1kXP/VWNpXOSPysiK
znWjtaqGk4VwqTXRxL2y6dlhigjZ4VKFkX7rVCnt3zRq1URcAqcxbmilVpRPc9LX
3I7Ia6WCtBDTnxqocTsEnckjNN0Fwy8KClT39OMXRBvQIpNJfqk3JUFV0ATf+cPx
c6HAFsuX0kTR3bh5oI8QG9tpWAZG0XldH6Fh1do8fccMmmzPMam84no+A3kMNLBW
EqvBayiHwf2pn65/STGuzy0NftHXAxfE9w/cm2raSF954bVtPiilTz245dPvFtLm
sUjKD4U4yrJVDwfTVuujs3Cs/Cv0GumDwnwv4wC2L1PMrUtb87sy1FAdjNZl014X
XL0gfWK933HHOXHBg3emLPn0+3X4drkFwOFgMjqF9nSvMogfgcdJ+WWwfmPQcpy5
v+USI4Ys55VYCHUTsG7wj40yAx9CT8HmcsXgdLRX/5+Gm5rQBEQwMGditwcal7rO
LkljE+jwKx/kn0Hd1mOE9C/Cl5GGs37BRpK0Ve+NotqdU1GA36i6O9A0lztxekvS
X8SxgEtWN5axIjU9CtiPSluR7/9SADzdgxcqNqgOsKwgNzhP+4j1dt0qLISFaKI0
vYXSNvZ2eks9+vPFlyULiAkKrLjp12wsjlz7NNvUoeDHMPCefGncmcq28KUzebwz
kPeISW71AQzRFoh415GpMSvQjUJRGPSIMGNXOU1myQbwCurJl2D2YvsUmihaHdSk
8Yrt0qYtirWdGE7jzgfxmX9xQGeTe75/YUu4/QhxC2HWlfKX009uWHVtrc2FvlLo
4ALzys/LTwBewsyURSFDIr5vw3Zj89oXv4yd6MOfneci3UtEzkK5u/96kthWkMZN
+zIGmpD5YYYDKsWLuan2AmBNSRYdUpxcUQdA7TkbC0O66Ofe/w2ZRul2scAo+IEE
y+mj0nusDERuDIA4SpLUqu3n1VLRkDFoI3M4KzX7zgVEPvx6oDK5eRAL/mBRCB/g
NOVaVG99upLdSgJFg7fKsrpe2yCGpLowRZglJzwhwhAq1eXNrb3QhavZbsmFRXRL
Lqrtv180chdUE0xHUiAcIbjAN6FHmYP3fu5n0FJZ69SXrv1s0IZK1QoyrfqJDb5s
O0REYlZCw1p0/bG2w62f8voAXnARlgXrmg7LhS4p41eWf7Q3cVhgOJzWfT0Na9cy
QI9jgmhD7tSi0kABQxlwy71UXUtrYXllWAAnpF1NuaNx/aksZbXy0AOzWb74Wlir
99Vsa8hqqX7QvqiOOuGjHwnYsq7SsP512ddDEFYXPXwoQwqxyabi+cSXp6pLngO1
PQN0R8L9UxswjadAMlSE8IzkN91Q3AuhZ7odnv2liYQYlOb8pqrBCsECQsDXNEW6
LDHg6OCj3bxSXU4cK+sqsKhalj0xBe26mC3IUQMPKOrSPOcVfopPe73IsupsQL+Z
cNAL0N0u8DS4lSkE7clwOzksz+BnAPGmy+TOvbA1rHpE5K0kL0Cdr+Z2wZHq2WDU
NVVekrZxYHh0g6z1zx2yZTHDYV0b4X2kxnZp9uWc3SDwHBUukZ+oD2Ge/xOovBtb
Xu0Kv1rPsFZ6SQYYYHvqcKxBXAP03itEJCBn/Q9dT6O0dj2YfybXmWOPTm3eL+xF
Hw8V2Lqs3Z9ehz1vDQhJxtM6W5fPb5Y3EmW0ExCYzuLBHElAsgBO1/N8gDJATHX+
X5HtL2oDJ015bbScH9rKAK+nfgVf2j2Ir+VvCd8vo27mWXV4X+ihYCrxPt+fTlNd
ZH66MzUkkiBTbu7XGhULVGg0rEUKQAn/522IBzLEM7hzBTuus2J2ARJ3TKYXT5Ud
04EmRD0c2sHVlxWcqhJMrTDsAZitRpgL8g8sChGxbmE5TPSE1hfQ+uaUpg41qWYq
qu8ENiB3wtYGzXjSOcPj9a0its/exr7ZrA2tvTFUQjBj6UovlEpk7GW2Jw29Ii8T
rl6gglRcTMJDk4zj6ZBHbqy9lTKnVSJeU0VoCFT5Lr/lZADm/Casrr9O6b9J5DZh
s8Fm9UTdH2j8smUXpsyN5TAFx1yuECJdzu/I60krbWXT+bG0JC2KBxbfDsm3pGO7
BMF3nbzZVC50cbCP9P0ucQLy9A6UPWuHby+nhJ9yr0xaWr5fFJh3IzCX6V1oYJIQ
kaB1hSnSB/Tg/DASr6iXSYCtgOK5y+bdfSvgmhJ3kfRFuynMH2jiwVp9bEBogtSc
bprzu15WDUa4Y/47AfmqRh9biBBvXoL8aF3xG3m0ubAMEDFpU0onvaLXJGZ3o3jL
/3JbUnZGZlLjDnDdxZLUYM17NEz8W1n18zhUF81BEZfra7I3FiAACJ+24xhiB5br
llIKyeS9KuZcWCNwSoALQGOZdoYdh4fvdD/DDSmF87BOqXS40fNWaj+MhBnW7z2K
Pgkf02f4bIjLB1ISu6Moo/Zk9AWaTFHdog2jN6Plv7eesRoH4EsiadYF4AknZ00t
JD7QDhsrNTv7QMjn/dzuuqOv0aofEkUTVFqr+EJy1YxOAIgqxnhwgJB4My7xsJ4q
NJ+Uw8Rkw2K3BobSJE1zZLMW0nYcaL7JY6/sjIdGoj6uV41MuWCmuzt5+ZJrDgj2
s44eRp5EROkAGU349FCnqZo6oDkP6m0Qq2vs3hCKy0GjHz+8Jjm1sLG0xiEBFfLB
L5Vf4GJGBwP8iqFSGMzj6bMypFG2RCsPDC6ef3M6TWN48kI4eNq2iIgI+jUcC7Ur
gTZBG0FoOU6YtK4v8hCzacwTc30B96IlMQcKt/doqkO+ZX8Hqm96VDlWqRGvhgXF
m04gd35gSx4pc8S+Vtgrmkwj8b47I6VBgbg4nOZF6wR1hiHGnQskwBSOi3Y31uGY
PzI+nx+ZQuQ0xi/+D6E8XdAeBAaDYny1jyz5b6hR1t3cfgM4Hp+H0CLxW3un7nQK
o9DcSVCGGWP3a/WwRQc7iAwZEBA1nGhpGRtrzrmHvWqTu7ac9bI0S3/yIatCfRVw
SlyXIZmzSztqCNAVS3Ey+UuYtoGzlQpWiDyfHPlzI1g=
`pragma protect end_protected
