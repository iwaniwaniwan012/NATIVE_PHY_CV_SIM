`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IbJN8ZoE3QXz2Ip635sNX31P5Bnxo2YdC6dnDzRHDPMfgi4F49GdFxC2yLn8Wajz
X7wk1KMvY9BKc7ZOhFcKUn9ctjeP88I42CrWvGKayqtXQ3i+qdj/YrM+r4P99Fyw
PtdQZkXgbmdRD3CqWyE8HWWP95kp8CaeORfE3Oj3w0c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 57008)
8soBqPBWA8a+QAxaWkqdEicBRIYLVUuXKdfnsmUoZd0gptDuqy0CXBRWriSUsO2J
e8K6bRYDP0aJpC+GuxJQ3offlG5ewLCetce68tqTnxWSiIiN4jkh3MHgZ7Hc9V0q
9hrrzbudzfXWhoCK7SeuApe3f7DZUo2gbuH5R7J/DJ/h/NirFouJ0LmESrCShpHE
61orTcwJdl56CJPJb8eTDhpGaeoI6/9pkEQJzQm1OXk97FbVqO3mxSR5rClW7d2u
RZuAaHPrXlVOwthOz+ujSxNhHMlbkFu++wK6t9/kheouAkTg0InQUPPmUneoEN0j
ksfRM6OsM7o/8N1HEXXh4ObbKrkQEWadjIjLL2t3AyLAbkhdR7g1P1xXBBHgVZAf
lw0qo2wF5ShkbJssV0P80wdm66jgYH61NVeTRLEdtrkvRU/V321COvzQi2Yr2QYa
z3V+veYftYpXqqaVbG/RZhj/RWaQ1buzHcidTmOnXEeJ2BqBDjmNZk1CePj6foHM
Bsb3DF7EdALlJma8awCuUKUmvYUJKqMZCPT1Gh8ufztPV8EYljCT+mcPIeDD6Xpm
8zUC1GmbvtIe1UfnqQA/Rop8e5wsv10lcruPx7BrkCpotN4YzjIsYj+uh2H8dYlm
7A+iad9jcSvhSfQFNmOA4y6uoHX8pe2naMXNNh1Wbw+ZoB5TLIijMGG2ZmTGtnFn
MgBFY0ptrEtJNO4OtG/DzcVrNhAgUpeSB+g/qL1VKT1BDRvf5k5EPb2bWCZwawt1
EII3T76vjlN25z7v/YQ9rTn9tUNIIfS/Uy0W0G0BZTnF+zsEREZxgwbu4mhxDWLR
gb/86TWbcFCUDynXlJoOFrv0dznABi4hTN5ZqSF7gVN0n0NjL1trVI3A08irVOn+
8d/7lz7SRxW1ptofQTWJTU9b4fuQJD+VizO3LJ6Qix5vLm8QGHZD8Y7KiJ8lINoq
l0BUjG5ap2Fe51M3F98H06jvChR/tJg6ePfXUlOKioAz8dwUozoFR1u6YrFSwBSm
tYxvU52L87vBL0iOhqoYNRnpb2S2x3xZSonICRC5OvYwBRCgIMiw+FIy9Gh/dwm3
5cqsBiaQtBt3GD7Zh+TKXdORDRWLMe2wdLb421MU9/RYYKIvEiBzguV6gr2v2kol
D5zpQJqi31RNpNf6fSf4di3zQdsHJExaq+pfeBn6Km7gefhnbkbMHJyTvbhD7Jt+
H/lTQgajkFdBwuTNy0nGOgFLEoozE2U+M6KsSbPy/urzb25V+vbk1qsJFjvZ9d1s
swsz8Oipzj6XVyY6nIO6r5xRqqbE6tYlmdiZYAKdDZ2fZcpi/LjB3c1LJw9MxH42
sLhm54/TW4JRYzD4ksCIBHS+DMhOQN+GyvL5Pb3UtPuEwtV7YF1G72MzSPOXkCLm
uDE0Dez9lJ1NEZLtb/pwWYd13ZkzN8ux9tsFefJlXdBsImToKgc1vnLcQKqhgPG8
p1fskroxUNtC17eGfZMd8bnGUT1U9ZgkEM1zK6Nk5jgrhUg5qHOmOo4P0jgqzmJi
uF9BLrsBqHXBKNdNXjDXxfmgl7ODjpI2W21zWoJfYVD8IFDGjTFBhUF9pvAbXJZH
ad0bqwQX7xh3qokL5Q1gnWxMCPkvx2BWTin6937KKFyApLsLVtw7nG7UOMTCjPaY
OEae/hDFjVaUHNto2yyU3iDeZ7SPSFGn2AXVDYRKGZuev/5A1RTl9TirTEKCvKCf
x46Suo0X4ssL/Eg/ME2xYdo7YBo34MwyT4v1tN1P8ANbQNVodKPzr4yNGwOjQRkC
byeaJkxAi+eGf1MztLaGWH8CuD4SeonFtIMNgTM2N9KYK8PXdL1HxQyIDb7A8RFI
n83U30Vm+/ou1m9xzTarY4glMrmCvqP4/1P0nmZ380A2pMP8qMHUr7jei9Qtc2e2
koOYo25RU6QnD7XRpxhCEoTcarFFrQ1M2HJY8N4cwaw/FfCC/Lcvt4a/KS8XshUc
Hnk6qV3X1h1Zw+RsQv7HsbTCDgds4iHjFuIETvwTmadOCX9iFPsab8WjTt3HHh3b
oiL8EBZJ6K96XyAUB/3EJdunt6vnPrJ8s8ulkjqEF9YeQ7kOXVkWdwUQbqXBbNTW
0mUCHYKLb+B7SM8wjbtwaUfvmQ/N5X9ryLUjbiGFEENVzKZQ4IxJiMCFbMsICQqA
Ip5UPny5xEBLvD9nlLtxnrtH/DsfbCPZnxZAI/sxTkJscx0qn191LVFuRPmLoi+f
4hKI8KHf+blhMqH3Ur3gQOiI/4kGsJm6BL5j1YD73YiodaeetE6IJJobthlcA3Rs
pKjAoGW+5lbi0JAwpxxC+poEUf2YzZBhRUJzrcULzhniVN2v65giqqKzkZC6qaH5
EzhT/Ug3/GpnZt9MJnfX3YSWiJWSdKVZ5iFVb9Y3yEmc9ReWnBfmVs867Jv1tdh5
8MHS54RPefsSAm8j3a+MUHfPo/rasfGFIOrJWQgGB78lorEvY0yD/Du562Vsku9N
vheszuHsi8bnQK23SlJ8Eia9IrgwEDQE4b2Uwh0nlIuhNdFjohG7zGDCUsWXdgTc
wEdgTXwTfJ0p6LY2cqAPMkpZ9jlGSn+Ri022z2HBSJUgsm/igeQWNj6EIbyHhRhl
EcdYrqin4fSEaXD/9k0mKzrgOE6tm1sXTxhmyH9rqaniDP2dw4TAEVvIgLCUKIew
P8DkR9IVWH9DSibqYJLzXyAZo/9gU+eUkI7358H8I0TNj5StHBOskeAiJiRzidph
e8tUp574SPKv9S5KvgXJGNc1aOFv2IT/cq78OuvoUyoVb25ONswmJVZz0iZKhUFj
5FWnhCV9r6nHXAFn2IHqZhnCremDaMYNUn7n+wLSRYcz1NSMljBVhtrFsRlicjb0
NihOXxHXt2HRWu0AmrbZ8cgka3CO0+areT3O6DsV5YiwUP3HVbCo1YWqSDVwLAaE
hTvhLe8X7Hxs+uLvMZrQyhCvgkGq0n+Q+zKVJ73EkO3xSDPxIflLSptXslqRmuHq
UBLfFkJUmYy5MYkO4Av+y0+0UlaTo86czWlLLZFKbohz+QIDK3ZC4rw+CEKNN9W3
WUUdHshbapd/k95FoZsr3nq/dUlmy9XOYMw93LjB5jgvy+X8lErENDsqNtvobkUW
LgwfogmrbVH6Z9jeh8ViOazdyQ1KuSuZkHeS6yzUtak4ezL7l1L7aLSFrEuTQ1QX
56B3q+rL7Olkymo8GB0dJTMALbmXA9gO2iUc7gZ/uPF3qFRPwI+Gx23kB06dsMD5
vs3V3I7BKyvK09F71SwArqFTJL6K7W/n+froxvTPjGt9SmqZB04/G4buip3q5E2n
yx/SFlJXgnEiBAIEmk3R8klf+skErhSzy7xV2Giol3rJqOOWF69cP1VmMY+MSLpG
zVbKjpnSr/LiGNpLdQLeUFSCy9HM6qjsUvOse0/tVp+eIoWWI63rfeWV9+GsRr5B
wbu+tgTkvFuJenpbkibHqeYiK+jHCY9T/ovfhWmz4GDyCigF5tlXu6mWvKjEi8CP
RuYcePFP++Jmx3oMIHDTgIL0YBglBpy3LOJTaPWmAR7ZzQ7CXdGZOic6+cotv65v
FvPBy1huHupKnojbltu07V/a52k7+KrNQjI0HRIbvh8Ff9QJzWem/FdEgV1fvET6
6YJeL8RA0E5Gao7MjBqSpkbx9zaLou+2A9d+NLRr5+R+Tl16ob9R2RYhtZ6UpYVD
7X+fpw2czAntyapLhKGc01UZkYJFtehAeRoi2M9PraGC0CF3nqMuM9hbJ6eJa1Vb
6gfaygrM+5DRe6/hGnBHw6+HrOLlv7IaA41TKyeznxPs5RXzRskzNGB9LQKtvSi+
64AD6M3UXl+NoworFvM8w7DfRgHxG2kcF2TFXwZJ6VgkLPA6WdWx8V59c+heX3Yj
hVyp34z9A+yOpKG7ApESr6HuvAuxdNLT+01ZVjMQo38kc8lOqGFTiF+GHRHhBHZQ
mxLe4PIDW7upp6Qf7ySGcLDRxCn4SCuYcffcsHTcKnoW3ceY0NS1GGsWj2tFCglk
EmJk0Qa2PRZaZhQXoEsazEgadxgBtS5iPMcYdgIk4tXnGp2u00MzYWRMRfrXb0Ny
7OoxyrNIEpipA86mOFM7PJ0sSe3y2QqGgZSZIPtKkqsNuOIxVV59Uzu/bXS7QqVG
kDmCUX1VFjMyI8dOm1i2HZ15R2UQgVJ+KeFaH8v42ObELoHO+KFsXvH5HeMgSMEw
+TkMmJtdw6VIYr6PPVRQpauVPaVJJuapr6CTdWg14rKq7w4UYngCm/gbooryJJLX
bMoUh86ky4JBBYnMUq16T5/MBvjLPoVgG8kG64CrpfPL8IPuOQopaCy2Qy5MHmUD
7ZSWHnnawL++o5kQ0MQRXEut0nRdKcRADE6a7dz3P+BAzEVnVB9NLLJhWw31Fi5C
k8GscJ4/F0HSc4SRtEYq9v20VtLAF3Dol6SQoA9FJBiwanwRQiQZGb0NVy3MWW44
SU0/MacZi+aOr98UcY95aeOEWk3JzvmhDqRyH58R17ToKafrGkw41VHl9PDoDKGS
USLJxTzI77pUaVX4voBhK29z4Bgij2aUKENfraOSiqP+6tnNWxewQ7vgxmx3EGBO
rZY6wVB5jfKN7IOgho/6XUKKwZ7YcDzFbhbvwT6G2Jm9ypuOV7Mc2KEnNCohUoih
lmiF3b2nghKf87qeeT9Z7QFJTOF8+dzHE3bvmZ8C56hlkrSQZkCW0mE4ip6Xzy6y
l87qeE5vyg7yp97Ea1sjWuAQ152Ix978x7SlOigXmhqirXYXlTicICwi3vZfdna7
1PXtRR3De1Y//8jRGWNUaeS2jTYGgdX4r1dTZ6AA0NPxfrQa0/d56DH/xKkdNFlX
eCQQ7EHrW8J4c/fjfg+zds9YEx2W5+HAhQ3KnDGZedlCcvqEZ6i43VrZZ89YlYik
SySSul4oVoO57jV/oJ66BCZsomJ0nD71FabWPaslWrhMiq5R19sxokvhCJio3fDK
lh806/Y/Rjr7Q3fcLaDMY0LowYd9m9dTZj06hVWPNXPppaEWSfxqw7bGsJPYVn8u
PN2o4PavPDEUrfTZDX0q2e7CNFiTVjh6I/PwuPKwqpLFx3b5VJemkcPlB33axhhg
DdIHYAuL5knpBikqIv485hiL0VRNplUnFiaEswUf7ygcB3qvm6nOjO3kzgrUpke4
DeWnxmIU2+hMb8ZX2E1FoBlRfTgAufsUt9xIVkoHYuUdnNI2aNoSveKsZ693opGQ
r2CCrGRAeWBhoUV6pr/8SplU16cOtz7cAmlfaTD0rYt+bbNT5LYKLMP6nEfXNXE6
Zb8LLbhWiZoZissLGJOxyx7dwRJWWy7u/C82+oDo2+p040I+wM7gqIawsYpMkJvl
iCpWHAh2YAa55RE3Ae64BIwhuMGgeAQbZ9h/s93dLiaU5mGLkecPBi2R0GwNKkTp
Nb9AZx+emSOk8SnFuGZpWwZajQyTzZWc3xFYq4jkkqg9fOv3QWWfCUiSqIfIR1uq
97hgklEFX/1jq73P0HotD3TxZKpI6jChDezccyC0efSLJDnglJ63EbjWL2eeqsI+
RHZgX7gpgfkkmEhviNw9kra2JpkkxWG1PWIKSzOc43cBgz+rWbWwElY9bDAl48Hn
ta7Rduxc1QyL/vJWKiGlNFI6SWegnuMDm5+i1XJ+lwWCGpGoKjfFwxhb22uPeg9w
6nKvSHSjMaAbNr5hRxgHedsLoBWZlO2EWkrabBwkV6LTBMILpCILuUT7qD8kziab
8p7WIOUUuGDHFfUtUiayFz8J20eRSJZBffzW8tesjgwSC1gtuHcwdriz7TETzRKf
dYdCA3icA1nGZzqhC/crJK0grso8Sm01T4UHs1gOQTA/RluwsR08ismL3InHMV7U
u3zRjrR/GcGXsH7SAB1w7DmUVUu5Knk39jAHeRBbI+TIDzfx5fYVPiUqlGGIOhWN
rv9vd1ehtvW6bRDZLJ5LXhb4DMztF/At4iLxWglfzUBUIX4rryF9JNBPiMi3bvdT
V+scuTouNHwtgihGb9l6LwynAOlPJBupTQjjlXX0XrdaeScQD6/MMT8cPpfjF8jw
2Umz+wcs4Rztm7CBZl9z70BEslQQvIWy/DPd/WNJ9Tt1S57DKFsraIAB4QZ91lOe
4I7NWgk/foqPJZz5PG4aenYB10kWTSwwC7uoxkoOqtKMV2K4CdIyMGryqMWgwINT
ZJxGVzSNp4dbpC2gsYHeJH31NceO4Zmta4BpwghMp/rIhSA6QasUoUd23tsNyvUo
xjxu94phwLP/75O5Rvf7ru3OJi1WgSp3Ym0vcotkiPWI4QbVSb/hbMymqFo3EK6V
SIDShrMrUffv7WrFHRMW31qduqGWl1qXkhpijHl4xcef4e6IUqTRCDNFOntFM94V
dh7D3MZESy6OzvcMTlcWUefK9Hs/yl0cDIDZozBhFYkxK4NRy+3fKKJeEyoi3QYi
VBvW5ImXd4idsqC9+YfMS5Pg7I++N4ldPa1lTDyzfqxHsuSlfaHb9TCN5M7jCTME
gH4Oaa9ktUHD7Yzh3OzNRweKuS1VnihOjNXDn++llguCkuwiXchMov11YcZvbND0
4bLJdIC4uOsz9pbsgkLrY5sBfaAWKvGGQ2D1EAPxWl+c9bhMWcH3REuECLF4S1V1
4CaKv7tb/+YlOd9FQkkS59bKLW5XjE6z/wrKuQLbrbQb8pWClhe3rJhl8exreXPa
lU1YE06tL7/1xrYNjkKD4f42Mo1Qnlrpfs+JvklvbIWLrk6j7b1BE5AnV2WKd5+f
F56tZTYwmAIq828PXmtqMsCSp8QoBnY6S9L+Q1/eSlGE6Cvgn45WDwlTWQ0JPc0e
XnVZGE/SjIMtp/C78uUieoONRxwpdmQyqKtQBd8jTjb/Iqk6SrtovOijjJ6IiWQF
OAi3xlhfr0hhvbVf5UYPr0ftS1yQzSF7xlf0GKIw7nwMjctWVzy/PLxpcMnwstpG
IoUEhZ1GiLxS4RZsGEt9vT6NpmnLhz+C++emVE2yCY2QvrL1mxT/HLyVAsek6SaR
uHeo49z/bs7xxzQVEHcYBw80loH/1i89smJdQKx4DLza2yUVqsXjVDm8pd7JmX0w
GgKLgTl+IxSO7PSkH+43Laz9EgASdESGHRWwfSHb2WvJ0zpDcUc16p85Mj475bBs
9KbSoWwWVd+olE/bN4KGri3UYXuQGZjLVVBK6ZXP+t6NtVHzoj8Rpd+CjkV2JJBV
jNqBP6bzZWtHLav2MTdNysCP6+rYtoZp0W/+su4ENoZHqrWtjC6BCzqPnROXIpHz
7IO8GWStoPe5ZAeSeH3xD3cwnYZjRZK0tEXuUOA3yVy/ZNEDj038vhnI6mMrIe1r
UsABPlYz0b01wP4lxDdxIfF/Ax/L3FLBBBHgn0RPxhuBfac6E50vYDoM7uc2kYjn
oAWSTlDUarZ3ddmngqfsXLlPl9aeZBuGY7/QmPGonGezDgLZoN+d6n6XZrTv3x3d
Yk/S0OuXtiD/8rx8YhpBsrIEZBYOFdN+seVESAxwydO/bByH+Ti1tVXDZ4KxER5u
KCvCA27u+zqCiTogSmWWHTGknUT/xH74u7rckN9aFW3Oh3eg3BrnqSsoIxa7rxgS
uyOxstDS1T9Tb3uXcf1hiPJtez9DrGHXr9xcCPWcIaHcY9us2T7mIHgJT6lbThFq
c4rEMbOWDf9LDyU9zZCPBBFeppHUqZp932oYaSpQ9W2xoXmt/qYSF6ZZFzv/DSEX
uHMIdMnabKY51uvmqKdtcysdcVnwlRPl3iwuFA68vIr63pzhduonpv5SADgp8Fe7
8MiySr9JICTO+no0vWDj66UYSNrdcWa3LmVu4zlnngI+k2ULy2/TzTh1qNJxP/Kg
RB+CWedmGbfZSFFXgn9GOif4I60tx9xDf8XpKTuEsn4WpGhcb/kLpVmGvcrKxgp6
9/HMhoXKkfMKUyKIVuooXrDJ5ePnuPM2WxtF1Q3wvQ6R29+igWkqIfaU8550wTMs
w9KMbnYlmz3AwDNS8McLZD7jigWvRpbLJ28zl1wNjiUhLudBlgszfL1RR8Bo1QZA
cgkVYQBQIaQmc44dDhq4DIFCKOGzwUrEjDjaZoqn05GrOmSXY78n6Hc+6e8OkNQu
bbc8d+OWIFOgxQrmJUstKkKXLqksj/bQ906AyZY8nM1CTv+fofx3G4aJXFLCwQVX
F8gNSWJy92ktzPZO6GYQxKK8CV1zTGG7QZlnhG1tQsHbGNk5ruxGvrtuxZajSWJv
eJo7pNHEslA+GNHZ3NfQxWh65ZkjVNlv8Aiq/Gw2tNV6fLjJB7lnbMYe1Csp4QZ5
B91Q0TrhTdblsRmYDTgUHlbxN+t204XbFEMt21bD0TgzmKyfNXGD0lFIch9qmSNS
2EIFMOyqU/Qv4MLJLczj/vz1AOwGJcLf8GhDkSP9AwFVPnZPajEeI0MifwTtUxKH
6zxXvos6xWErT/tdxZNgdlRnbLnu4jYtZYNAEF0kPgAy9wKNQwfy7Zp3C6wCMLaR
m+Jvb+/BT+3W3HiKBQsl7dFS8pUItec7MCTxQbkkXAjyHazEpt12PHG03/XKUF7B
ccMhqRKAZ0VGNQDo730JaO/7NnHBZIfWAvSD0hHJ4hejGyH40WEWWgzfLlROF0C4
xq5zraqwsWdg8LN7FyVfDlKTrDQAfs6DcsRooMv1GNaX+tTBCvyvpDALZH3tan3V
XlQzMshTCSd19FxEKhe0f8VYaNFijoDDaF9/NTl5bSfDlM0KnbYAVxc/CwJrT1Pz
JbV351qe19O5OZBeVfzIDd5bFRE1gwMcOJlIKqN+Jsi/a1C0bI+n1ZHpioGAHlZo
PK0c1UDjhDW6m6PP21bh3mScw6VEfoyPcZsRPHQoCipngD0cnu9XX7CBlKasNQYB
FIF9OpGTCQBHYVGpHVCwwCy2LmPuQYm90ig9DbHWSLcZ4AS7FczqCwmaH5C9Nbjq
91L2ccrubimU70CvDP60eM/8U+Uyco9Q+FkamiMQEuV45o2lFBA6noRXGniSX6pJ
f0E1JAwFPKUEe1JzN4M/MdulJ2qNfTOWwAGCzlG6kd07iogFFcSm6YVs5kDIvgWY
E7N//n5z5zCcgw+ArN0+tm2V2eVZzSiBz3rm24g5BCwXxP2S1pIN8UyUWkzWLaDp
mtxPL2QHiIT9jTC6COz1QKFWCyvLJZNuHygt2gz6hlv88CGYEuHjj7cArwvTpWwr
EJJ9aLTZlodhaPs6vWNFdoFLbGheXNp2lkg4X8PKWcgi2lOOFWcUWbLKMf/DVbR+
OIaAfw+VYXowNJnZgkP6njS6E16Kij/zv/0OjuUOd76wJlGlYnTXlzIW+9IScZ8n
ZNvHtQPmizE3lfDv6ERmDTNKBx7pBW7RI+sJI2MLaaEz4QacrtcMbe24ciQuvMpX
nrf3RQeIW8+WMgfh5GY0ERtKO0CJCTrN9NjJD3DPS9LVD76zFq1TcKoRWFg0BjfQ
KJpmQsFrQ5ho6ImnkmnsLlCeFE9tlYUQDCiTb1JwhqDxnB1gLJ1omJ5+Xf3PvRGD
l9YPwLzMe0LFZlDf0CG7xdtJJFH2cCsML9kB5KqfKASOBfuVL7dSCrEUhXl3q+p/
/0QTgdy6hmisSUhcIsP4mqA4/ZKBMZIzTondHFmGBfCUYI8UcClVr2UEFVPFmvbh
QYjxJPmqEKCIcc8d//O8ATJ6uiiUTDzZp0PS6iS2FEOFUxM4efaXrGGFoI100NJY
gerzCNrOP6fL7gV96CBmMJ7MTGwoVqS/pLjkd1gMZ1tuCOpTXLl5m2iOfsqLJwod
4tNxCpb6FSiCkvBkildAHPizRqztdo7OSfkHR7x+8VQ9q0y+N0ZbwHaMBOaQsaGm
AbXHRWRIKDenGNJfMk6wbKdW0vovz2Qw32lDEVNTvfIa/KgmKheR3XhYwF83w0g0
6eI/1p9OcL3XLQZF8o8RI4d2wQXGSpFUhqkj9FIck/cHMKoorj2yQWjAChPUzWM5
toDvRbMyo4ksW+yfVtA74eg0vEHmvzTr6wM/TvomT+j36UYk8H7FdEcrrHUaqTjJ
STh8a5UmqmT5gehfga4HC8WTqTb6XnCaSIhDVAVAaNAgMAojs3r8GjijylzVyuaY
IhcFUE6hpJd6EPqbvWh0mYF6lfg4isuXiqUUBn4sUO0+DI92xCU+mXBl9mhRLxSS
M8XNYQZldDozM9Lmmg3Rbyt7MpKe7/2s5CghChpNlxYjBx1TNleu6c9MCxuG4eUo
F0UyaIXNInCNxxVpd1UuRLxdnVYHVMygya7ys16a9Ki4Cznlsh3u3KVL+5XGA3dF
2UcWPe7aiurGnVwpngDuGflKJQPmKcPxaGTZWlE5PEEWu3sk0oGfb+YOjtMxmRnR
jAYyEK4+Ewge2B5XuvrtdcMRRRqfXmjquQfjDxOUqfmxay6q6iw8BaBkyRSeKZXX
B7BmebkekXuXUs4/eRsKtnsNljc9eCQST/PNsnKawZi0FMpu9r8ByGnxuqLXEXYn
+DTQvEjchCWbNSS1eSoS/9AUugX/ixLgK3tr0TUbk4poc8eGZEGVzVjq0IiYUPuh
Tt0wp82H/U4VAugGlaZvSgT5sK+H1VvULkGbjIpTa3U/qJB5IxzwnhSp3UV8RHsU
oOtA9DSmMr126VOt2vABlMlS8QKkMaHdQ3M1KI5vguIhP5a8c6/fHryJoEWsJpbw
siIgI4sHbHhecsC2Hl4RogoCvOUcdr/WlJ773QTmYmJ3+9NiC3gILs0SCjZm+hgR
6EUbX6Ms1FNMLmyQ0B2bZ+MrBc5xg0yAfyXYnTP7JBJ69J8Qa2hC83ZQmW4Pl9Xu
eevrQLSlvvgHEY2qlNbOCVkHfFmYhy5Xc1AmlnwAijr5itCzPZxThztU8nJvfiU7
Az3zXx4OV4zT76gieeF+nrRjeElo/IkTymCdmGgwZiHmgSr+UfWan5EXkknv4xi+
bq2qBpknNx1TMYDdNTzZqvio4HzfC7M3j9WMWp12RoNKwDhQNqlY9swXPv7UJ5Jm
1vuQ2VC6pyLJuneXNyyTubLVGqdjgsG/LihVSx+JRAazvqAUOGd3QSiwFNPnQvWI
iczFIyiYoOmOh3qcJEShY8W6eDeCeJz62NgyAVNZhU4+CLYDsqhgMo83R4fQcYbI
GKtu7FrKplWk1uJEuaX5f4tVDDabKq9b6UNDa6tsASZvPYmkdUspfrxwOqHULM7V
aOqxUJfKf5p/TGT4e0eSczhbVqRzCakFWP+sWFIRnH4TxZt2NTId2IXN9pEmuF4j
MehLzmR5y+feHRbeY8hi8UuQVS3hop0dtrz315bQziFPauiEtrAxR78Dw8v+0QH2
oB4duItxtw9mbNYzyls5CRRMSY0ncaGKB+7azpWFyOQ1G7NtTzgUed2R1uQtexj9
9n8G6N0N0P2iZxJ0lmgKXqgHFfgjD0PbxqrfSbvlMDT4AWLQ8rZ4VYM4mzRQjv8/
mmOwKZu89rtLfQpvjovK4PofHlcVe+Ipd801qBjDCOyB9FHc4K+wuXwlHua5hLHQ
Jmh2RcrKkRDlPzO0dGbRpW293OeZ3Tjn+hXApRcAkEPZE+E62RLIOnsNRtBp7gWo
VZ/YCBPAz2D0+CEWibqZ2Vf2W4uRGzyp2PSKonSkGPzFvWYLdmiGevRyWj+mJZic
7TUD2t8lBObZrPjuNVrF/XivTqfYbAj8Sga+D1yA3Rz7cNUey1UFw+2Most0TUzR
XtvUBd1VRxzXbfqpkoDVdnBu8qdsxW4hWNll6PBAL/YcTAAakJuZTG30pvAyKPxt
YQnk2EUFCiskuMjP/7y3fgc6QK2O30GuKG5jVULLer8424x5neyX+d2kQGjAStc6
/KcvySFNxTxJsmGfx+1fpWYF1751ubqJaUiBWMwWM3t4Y0b1UyqKXEC8CiWLZqz9
hTxRKQitvK/5NJ81tee09w4B02uOPrWpypcihUoS81DaRiJkAq5YDeLRslTpXAS5
HuuMvLfM8Ip6NDP9t8Q6Fq0SaeZmKVrGWiLkT9aOcSCBEt0gKXG7sQTtGQG+N+9s
4m6CznStXUc5eSuGd1wysfSwomoUmdm3p/8F7qbry5qOOWWiPVFhf/3lbt5IgL0o
SGy9MgchdADl1m7d/y0WcrkF5kZ/9e3KACtsz3iRx52GTuQMUq2Xi4NpUZ0H8wXw
UWmg1UeSbLVDIv9FwMsgntgqD942VzfGydhGkjrT/TJyZE7Ym/jt8c1v20zTkuHn
Y6qr9IStEZBDtryD38xXG1L/BR49YIflMjMfPXJ685dJ0Cc8+moiSYZRwyl9orC2
CS3BeUbwZdcRJA+6XB6ELiGwv2JIObSXJ6tNK69K2D5bl+SjenRMHAxPMwrcnMqr
mWlduAjPoH92z2gUodFC6fxE9RkMbe0z2sG3ottaEOp03EBzkxmhJZmQDAyd8PnF
roLDu6xXbIgIaq2IfSEqw8B/Lq2MkN6azBVbi2EEXCHmo+xxpXQz7NWtq24Wn4XV
CSuwhoFEUJm1CwVSFrz3/DzS1h5B92AGaaKeeLXs8ErBtH7SzdvcSsHEEQKKasyb
fvNZRZJGnveARsedDf90x7uznbmbGSkZBbUIhMueRLV8kYtx4oBIV7YrKCVYzzaY
ekLKwYY+ld56Xxa7shcpsSbd/zdhkGxEBUOFlHZDDIi7G7HSSn0Kh/FXE5mc1iEo
fSr14i5UW7MV6Dx4mx53yRhAt5nQ8lL95EvX6D3ALiQDhfbXaV6IeaIDI/Svxuzo
iPB5hwLKMK7mRL3ToLH0Hew45xpldBDCJ0owHXuuF1dvrgGxZB0Az5qNMJcUYJ3p
9icxRAZahll3UZyOUAiKRF624fHNP7B1OESDzpYFR/hrdeDLthCJLohJ1bWIOe7T
NB8WZWWieKm8gxKhod2q3U0f52M6UJQL32wcRrTNDu0tDCOjQec9soxr6utfCyaV
fdiDzhVRbzgOAL4OlqeQpi8B2pfWDLMeHPKWxXH5wZE8hwW4yhqSRHGXOYlxHWk1
G7pvY41lAsQg2PC+tf9+B4KxDp1QhojtgDbHgDP+YPRcGOyO/UfmCypenhLzyGPb
/haf34JYArggt8+YFRr7W262BW3wjRc9g69WTvuVZ8WiqkZDI66PJmJkrcyhKSTP
lrZJ6YfxzcJhxpF+Gvd8s/6gdwJl+zLRNyMgKhlNlHO4s82BCOBN52DgQd2DV6vb
LuBeeTIAF0DsObVd4qLEiM7EZ4O6yWofVgEi6SVuzuWrwBq1A+AZO5nneKCwlEiy
LtD27FBecLEtTNYHBk4GVl72pW14Oi9naScSDLuTN+ornWbAUVbsDDn3aQ066/oP
kk9nI89bt3s5HpH6AfRQrxLhKornLywwhfEQR1i6RzV5iIz9P5NUhr/GyGw5o07N
ylGxnZB82OW/uY5O1LkGKUp0l8ERereAfg9V2X8t7zhJqRHmchwlVKfulMSto5F9
S2xZ6s5DOfuCEj1232/Cqo+X0Ppa+Q4yJNR0wTbubVO+xjp8us+ftYchYZs7mGQI
XsH/921GVoP0zrpLzCVPOI9j6J42MQFSwJ+41IgM2CbCnn3V60ZRc6MeDDO04CxC
IXFTRGMBi1u3hzxxhzy6BHIECRhOjehauyt5DxRm3RNIqEZ4emvh8b565d2y1XJP
Vos+14jK/pp56QyoX91K7OACyCuykRKGZeWQwNbQWBelzJwK5p+ecLVPWMb24QC1
GvaZ++nRL/g1VUMTzkWw+OucLSmnIhvakjzJmRTPJKNoqtWa8zmXqJXmz5i8OiPP
3nR8SbILqbQr7mtQdncVFLYjT2vsLqIsItp34KST2IGBVyHqRarTNG5LtJU+VrS4
lP/VXwmgfHo8KQdbgEf+okHW/Euz+uwPH5LFNE+DCYVRYh4lsCAormRO62Syrtg3
R4xmWz6hoZoaWRACxubcEKajZGVE8GbCjHtPaEq0qleCoQRi8NPjZINQYCGMCAMa
lUArfcTGEjYLy/EZuASrsGXDj74Hrgsa8CFYoH53spe6HfLtQTNrS1nPoeB7Jzce
97SrVjrXh+sEE4oPVejzNVA61vmGlJoXiTt0Rme3DlbPyfg2x3FP2v0wogEb6Xar
BWVBZgAiaojiV2OJnxPh7nqUVwP0G4MwJwsnCcZz/NK0amjm+y3kTCM19HE846ji
qjPxD/eSHwoQ0i0ZuEqh+oJfGuuYeirjp7gfQJo3z18jSu/I2aUdJCoxSR2OHLTd
ZlNhdt4axvQhs/qxeY5V7cGzHAh07Sd+Aeriks6z3TsB36/oxh+v9/7skkBbFtyT
fBxP7b3c2DkSah9d+KshP0io58iCeorQ4/vzwJbfT1z+G9vm1V8Lw4kiSuw/Dq0I
NVn3w1+z7x3u9ZnFRIvdsrCxTiTslw7O9kQd3YAVVddEd+sN8DWwSkvyXyvhzRe7
3l56Nx5ck9lOCGpQlcsbtZngL14hC47d34tIY32cH34h0ortzMJAhdjzTMvkPvZ2
4wzuOdh6f6RAf9PDgA8vC7UyRC2tO3StLa//2ZK0Wm838lX6j9GuP5PgC5p6Xfw5
nPsKRCQ3Iaiscnkx5cJcb2YiOIYU4ncAEMuAhzGlckJXp7cX4f5xES3iEeE+vf5s
YyCtsbn/oFyxGT9AIsb+OEqcdN2PnAuTQwBT1AFo4gML0sE6wUuA/qszEZFms4O0
b1lUaGX7IyYL+90ELx4Wd94SehJmhfR1b8O0QCAvxdbAkw7j7ExJuoNqFDe10Pb4
9C94vvTx2bAX8u7wpBE0aSXPQEt3ovDmNQleA4EBPEcJTt+3674XmC2uoqZX8/78
2jPZV/dNLgu7+7cfsy9EBaUeoxKaST3ccCMJ9kH3G2K80FQ203dTT5VYjvREB62B
IL0wSeTgATBeUCh1EeZVY4zguG6xF87KH01ORrxMN1aJM66S2IN9vizwICy3MExQ
x2tuWk43OoWx/GT5/bn2ifvUOz1AnylgXzXI7x6HfQ+A8uh/2PwpBiixWC7h2BjA
MpSPthJFCI5jk0h6hdR0vL8LN7Igd6my/aWVYc1ASlPnjQG/kQSRdv3SpLzXCLnO
8/CwLZvlza/IaG3v1b1CFKTzqrRqgiwYTy4QlfDTbbKC8dSnWhmO6jJ4C1sAzYwi
vALSYiAUJN9Id/73qPP2CmDz9GnWebBSFgJeADVlBhgyKYoZpU6EwbExW6L4CIKC
hmdeZs1v9Bk+njxCkjJytU0nEdzEQdkJrg1zda90DZa/SHkRZS8iIoxeJjNnvrsz
54hoLYy+DF+d9wJbOMoTikI1bqu07OWUKYO6p1hrYH9y5SwovXytFUxbDRdL7Fp5
nZh6m0ea9qPUkddF82d9o2joj8eDAEdIC/9Skvr7AVQfqjdX7Hm0q3B6Y0KNRKnO
6BmnGtsZtl0RtZMPk8oyyn8CgoUju1JroR4ZhFV8LakMg2hjwyoMU6wM0/Gv6UdT
8toPq4ICT7Ob1/9SpHBULbynnI/c2QBJmlupICHHuhAw8rH2NRPso/sBbGGxYoev
YTZ4KJUEWYNYBeu8LG/dCr6R20Ewt+EPLUFvVYmKA8CrZtUZ9P/HtPqDOAmYjhm0
eIpmst3kjD3TYFLgWELQgL/T1zg7bsldh0GU1gdG/EhUDjD4MwOgtYDLWbAGVLb+
Z1HS5ukibi3eFhu2QKFXiFSYe1aRoiV6xEHr1fDeF+d5fY4CLjRDuy1oUiadLuyo
voQie1IML/sj5pjUlTFlnTeYKIq5JnOqdNtuxXIDNxVULhwsEh/1LGsibOWGLRSr
55FhAzj9qAyQsNl0F4bjfcRcj1n4Y086Gcv7M5ppxdaYfQZkIluNN7wrHRPwemRU
LlsNB2k4xEHHRYHhi8eAlQf6X1+2wlIbWDYBFMT0JhctwruahLJo8PwUFtQzJi4F
lU8+N9/C45flACsvACGDS74tKTb+7t6BVFi8SvMIIkDhpQ9l9oPNXxBDc3hnfS/9
toYyTvtfnkTKFpTOSoGTCDT2GBYFuzWbotgBbowzZRxk7NrX9i6Hc2nEFE28M3JY
o1ZmiPISmtm3+2YI1i+Oq2J5OSEdQv3KYSKc2xQ26TavJQBvl4WGFO1HUF0c9XCC
JtZbTCDdzNNITLPdvD1TB8O6wQUP3tDknEYum29WDw2hsVOAKWzB6JSgHRpLiqzS
ZotU+4aPR/9/9NDN77vozlaFOIBGx011OX7Hsz+qnx2l5FXkgDTNBHb0u5f8oBGo
pc+ipL8FMnuab5aDeLIKlrvRyOXtmdWixCA1Wl3nQyAdj7TH79AgypOPhq/WUcmb
kIqkI2NVRukPI7QtJRXTpn54Yjb02lor+GCdOCaTk8r7Z+OrzOeO4Z/4DLK903bs
iYRlvCJ+DEz86iyVfOPxvptY/ju1LoDS5vHf12NCkfKCX7TqWUfX8sb+HBAIHzP1
V6Y7s5WYdURj1i2Rbq6tEeZz7lHk7P6ww18I+9J3OCZ6Bcv/le1bwrIr3qZWa/IY
sKsGe7hZnhcWoJvvxoT/gds6XWP8rIpQAjB7kppdmHov7o7gWAaz5Sv3bPSwjMFp
uVT/PWGta7qyjRjpd73w+tWhpRdRKUEXf37K8FX3x3l+bBOcyxGl31Lka25O9jcr
dEdBITJVFN3G+3Y0sHjs0yhxPavvN6f5wuFSIOLemtSynR1p38hNMNuxNSJMyPTs
o3yHch63LkGUzntkfyJ6jaG44+YQupTUWYp5ZcA30+Ru8kkiarGh0ALiqAq2I7VV
rndIUsnD5/mCFxyyVREhgIAc6k8/q2p4j/3azqd+0K6U3ECxHtd3YwzAOinzARsE
hYFBVc+nkCPg2jGzSTWcPB8hOFX7s8cAMx1f0BvrlHZk586neSG4nDYEG65YIh7r
w1CMCL+2llHn+ZvJMlOead/kIo9hmu363prsbfPj7FesliH8BEqQGUYmQijAqR2o
6DZvKAq92xPAiDX7DoTApipbFn0/cSaO7QQ54DmYr4s/Cb4yJd76GvXO6SWC6+Im
9mGawqQPIfbhwxXZfWD3Dy3YMVSxo78PaB76RHls+oBZgJN/GFmdLDNioxwUK5VX
nfp0B54GPCDAvUjWZSGiuI+TOZ6wonNEssf0RnjOIhkKdsDWL2FWViQR8gQAlnVe
GacP/LfygKwK6d+LpYE76jsLnGKqE7QUaLe8a0bNrJ2Pi8kE3qhjsjz/sx+B338C
Q78mnvcwvyM+Rt7k63gBhdIVUE8SsogQtvS+5L2rg7a8CJElqDItozuM8CBVxleV
JCpAdwghZBRxyxCF7UDOOkDDcqqRCw0HqbAj4BWChu3CQ3ISL8GPk/TAjY8WGc0y
2pvUJ5smSFgikaFyxfQwXGdx4KnkwWeu/lImUP86nURW8m2OCQjjXSSuzqUdc7fD
OhrcOUyt5wQte2zgxEAdTsvwU933egg9E2tPFGTZfcarOkwKu8si/1s/ggwMXtTz
eGui09h9a4FuVZc2x469gt+aMdtLXmdB6Q6QxXoDlB4eMHYJfhhtpa8elBxgRa9R
KxUWDtYPu3e4qRw00rEAMBGR8eI3RA3K8YFoUndZe09JoJBX1WeADjVh2AtOoHzS
cVbi+EU10QJuw0RnD84TdVgtp6+psGMnRlHdtEy2ht5E0fKsT+nWiRECo58sAOlP
wDfTOY12lofpDs+vN/ev8bNeA5UPes2Z4dXNP5sqxXPnxhJiGHcwJwk1npKV01zE
fp2iLrVisUGl9FrSF5+QVEIyWc/GE7RMf3y1Aa1mdb1RLsUINbxqx45HPcB8WMW/
e0ef3Bp6Ld2dHqHu4Cfzven/L9NfGSBZ3dwqZD4SlhoyCDPUxbleA0MT18srhmnW
AOEMtnjoUeIffYGnEErwjSyp47Fnt6jvYGHuGOYNchlaWOn7MVHxxShy3Q1LEtGY
VslvJmRdxZxLyamwhMZwfixvfXYMCTQ0legt3nz1r6BdzYqNEdMD3g/11Hs2hGP9
EdyBxN7W8HxGjpB91SBqZ9LDxJ+NKuCAUjtscPZB0FJOd6FfvC9FyYddUQmjWJRR
dNoRALzHTdouPMlKpun95tlNBaz0LKVbJs7H25WcEH4x1Ex+ousx8w0ylpz2BoGj
Pd2lKgX8QJXFK96SdSidzqOhO1iNL/jh7ZnqAwFjg8jpsDvTr22aapRLvtEyeBIK
lKEiacN9Tgc/2y6Q6C2z0yQhLCJ6VuNpRZTqAvZk1W0WYrsW4DOY2jch3u1kVjjc
L0PP7lE1SnJW0sOpmLyz9n1k8FIAxWoEwi+FkXKpUbnjnKspQOdhO8atup6O5a4f
79eOO0oWBnYPaQpVM6GKCuKWmBCWmCkVQ/XjKt8ro5jX0xmJpIeDZZ4XS1L5NpHg
jbX5aRTG3NDnTj8R85XpAfjst10jbJskR0E8X5Poi/gXL3Sh5jW8YP3TWgefyqG7
T+gRC5igqdWIn+LKF3MyeUD57cqiGPbPs8nI5gPPVe0BKdJOtu9fBYjJoZLbtxIt
tCP/tQFyZyHkHsge5DEX6Q1MSlBYqxGZdnIArKHz8P3IbtkW2yDVi/xZrB/1WC9Y
0uM5It8fQ1Bct8HBimXqygppFgqVohCIFI9alKjLWzLy+MjRgWG6boN2L88dF813
d5BsNiusKE3SgUKWGdL3VczCQXzRVagkNg/uzqFfHFFHYqGOX4wLd0UCgJmVgJlX
+KDRitYRnGFQCCM+6PT2bauZhlp/nVNf++PxhE+nEoYpnHXfjXb4smGYvC8bvvMl
V31n7j+gt4fWI5zlwI00MeNfUgnehWVy2jfQ1MFgLiaF9Pa9OrYzo7QN+CYlhg1/
qez4P0dwL35ADedTRt7uJ+RwDFFazlRNsYjLgE2axV5czIKCxRHsfb2ke+q5+LxT
tN3X0TK3nhuRqehK0PB4RfGQ8lcWEGd2jjFEJQ74HgmCISuZFLnBmi1jdo/BdRa5
Ob5bSubC9XD3c5Cqe9MP6NpDxy4xsSxt3Gt97sR04cNIP4Ajme54ZXOiRxmaLJ4Q
IiFUJKJ1V6rHngofRV5X23yAl3zSuejwZbHRoWq7i5PG9+2vQSt7DHlFMBqF8g5z
ICJF3Mcej96dfQgJ68BMSKM2eI1o5ozgBeTfjexb0fuHz5j/nsbuyHl62cJaBiT1
SNS82fUi5XC4HcYf5TNjpiFdf3j1jPCbw06BnfJ/kdeZeGi01Ne/Zw6jseazwjaA
HJjmndE4mwKU54y9cjYaLBLMVHvgDrUPxoVM7m6N7vGhzRVC/vrUkjPJl+1xxABI
RXpwQNrJHW4jmruucG0IL+yq5iqWu7bANSPCTHTXmtvoSFN9O3BMHBBW5ozPekt4
GA0qVHvnupI16FK33hjOkRUNsgSUYa3uRcz5XCJLDn9w+m/VfznMSU+1Ne2qsrWE
kZFoIqzIvdFxDtYQJIqZUGIMhWrkBdh/VhxMiLEd5rGrAbRPwaHeAVucnRdvuie7
SBFdfOztYU/4o9Mpcf7U568GgNXS/XRjFJ1qHGKM5BbvDpUcBmLwCjBqOgOwV+89
BbyYHS5erYAlz8Ptg39v1HBNv76GBSrYVC2ZdXmhDygYsG/i8krZJEHmx8hlQYg/
MOX+S+jTZk0UzumFPcCPx5l9RcPgSGAyQDW7wvnwc4Y3xgeJcEJPTOgNrPzTq7nt
tjqhTUI4crWAcYolYj6PVCOjWDept70RgvCvseikZ5IluJ6VTWxu/T0ReAicStIx
uxfIXzIt9uNM93+4/qKGIScTUdR1QzyZAEr2sKfEP+2t2iIF/CE8zrHV6k+bVxHp
QLNzdBXA9hlbLYEKNTtu3LFRbz5BZq/pjaN9N0OQ+7TCS/8d5kWHRcC5ITFMJyzA
8MBanq7HNw9SdHkWNrexY8PgPyUbbNzfwUzMc172kSyZobuxDZ574Oy3CvRrIO2Q
TFMBNYz3lbuzM4n8o9+TCQ6DJyArqZMuHEY9PQBadu5VX+LFF+BDNmDuQ+VcYc7B
6O7im7eseWW2PVdDnxDo2rHrcJ00h4X8JUPt7NbY6YrfaEfuXk33eR/E7tAdmzY0
hcX/v9+gMNUL3jIvgEykmAfcuENWwk8B3cYnhcHWkQX9Xg4EocdpKWO5S5IVM4gA
HQ5RSrIH3Vfq2vXVYeKg6pV+ob9PHCQSv8x7eraHd2ylahrYnP2rYy/NprvRyxPe
Q6ntIr8v2/XyPKhsQW7ygx/yRiqtHaenHi8oEHWV+RbOpq/ugVWTUKXO3k5x8DCm
qaPzFrq/UTlsJL2vRdxjcU50DK1WJYWZ+r+CmoFzqjcraJnA0XY0qvk9c5E3oZju
EswSVjayGQTpnt6jLZf6kqv3jp/v6zjgMWeQCQlYh13Tty4uRIW68nup0S1FE3uJ
6zDugM/OAIeOwXKc1qxexit0QzS8CsneKk82NB53zy6UiWC8jeypDGG0L5z7yNkB
cDuGjfPkaSfpKpSNJIC/UBdry57BfZptH6vjWAf/SROsutHKzvKd/C+IkLifHSrm
+9pXdNGczjyFuFZUaJNcwek305TZtEv9hLNKtAqxAtgoCBcUwMB3kXCTSOx/ghxK
s2SvdOWp1OFBBNQSPC40Lqb3fBmXU78PvdkQo8YzN6rjd4Ug0YBoV4jqiwSuH5yh
/4pJHFWhSVOlQ/zcctcUaABarr7SQ5B9EMjQ81ALO01C5Cblejox8jh+6Kwet7nS
BfNtlN01DKPNadKhEP1rCOwnT4kjSjV7oL1+8UtjuL8Q3RxS5Iaqlls43fM/wXTz
VNWfUBBiE0DLpED1jPvx73fWYiEM7SbbaWewsqMNWEF220xGaQ3kUftnl4M82e2S
iCS1BZqo8NpU7yE9kEu5qdz0DeXC0w47+Y9ML5NfyCf1DY4BFGjMti6C+/Uigg/v
mZ1HVl1UKzXimBYEATyd6RzsYb+Ys1G+m1Nye7bCDdXJzktpM4RgY9Mryeh0PVp0
lHEvUZyq4sBwe4S1EndJ8z96dJjh5zPECGPPw8oO66ZKTJGAT1ODF81xNM7841oD
tLCKzIyv7pKrJM+9Biol5PBmEKaOdxhA1CHMfnUUPBpCUCSb11NJ3DAflwWAsfoJ
HmtRwVy7dQ04y9Sl9PCO0ufKhRuCcEtY0DsjjHKcrmNLFGkqnM/qaGS3IkQcMZLZ
b3XR7mip/Hry5KnTRWknVeEDsmp6nMSQKPdNkXITuj1A26u8lNNLZSbOl19d2pnE
SqF2lgM+dE0VT3XMh4qL6a54bsyL14Yc9ok6ybWaixu8zzQF7z04uXjfttlq8fwG
jXodjiF1F3Ek+JivVQpKRypGT94vSxdJ+zdgqEGePf6JOxwngN0GIvxrcReWzRNN
1rZnHzapc92wXgwketOY7mJPy+IMbDW2Z/sNOV+Cs5tvPktBAC/aTG3ggfEJZ9LV
9woiR5OXz5SYcLiKNirgg/gMXxnmnweq4V3UraCIBUQVVzyjeDLo+VP5GA2DFscf
FGaGpqxFz8/AFHoStBDU9CyZ9rPA5sREYzVh36Vzbajg2Su8dl9niLuZZ7E04eic
HZ/rtNwTVvFAuH2+ncW59T4uW0McahIA69BbcpdHbly1qK76PkESEyBq2frLK6YH
wAWsVQwWEYAmPRPRSRGNjrx3my8TQUct9mVE6n2F1wFFXEjPYbJLcorJ8EaWb0ZB
UhV4aw2BSooWtWcusY07PX4+VLF1lGj1pWldZOLU3X6ynKJjQUopKPPnmH5koceI
NYzsAPbNMfSVljBhMzIRF54iB2l2CK3gJFwioESyZLMmrLl7wrfe/LZQ0gR7gbj8
9sGl2F93ozP8U1OaxqwABglFyYzMp4MDJjlGwm277AE5uCwvWsuaqXWwQldoBiI9
BpDT+mmSPL38vfCgxWdXwzJ7ZWh6P7j4vJ73MLb9Xnnqe/G8ULXPqAGlUM/mF0vq
zK8bYgydz6diR8ZjzkyMMT+gXG3EZXig1h4TeL+1Ho/6zCDzifOjx9nXCubfPvLr
KDrcgb8kU2gpjgRfQBMZ18umgAhIi8dxmz9V7UAFjq2PgyjSV4Vc3UHgQfiIUMzd
544KIfcrp9drT/p2doItR8+jyjh2Te/dK6cQMlCVuMvxEeE38YJ9XWxJ144r6l+G
AntQVum8TjfA8Le4BQY3r7k5hTRrXyQFpV/w15FvoJI1l8PaHRuknnK0MiYPCHVy
HEPKJEITX3SVZllGwq83N7PaEjTDFIUy/KDGV9IQX37iYtgFltXTtEtIURLZRleG
mXti5lpbE4BODv5a+VX5SAl1U6yb9LAt/Zc7FRfuXt6+aAEG0SNQYVZPnV1arqLU
oMhEuV1+a/Opu6yN+R2jcLnP7jzbZI+hCtOG6/4R+lICzekWrFVnQpRxsSThlFvN
BCmxGjrTH7p+C6eQucoHGG51aTVpC+oQr3egE+PbYQNCR/Ie0nDT9DW946tYdTmR
p4frFsvohEVcnmjnPYdzoTEwzhXTKE7gNOy1J5C9jdaz+5ApsHiGDoXe10Ul/hYz
EVbsRZZSi/lw544CDW2Nt9/tky53Q8tyErUIvJQbD37XryjPdYoom534KTsUA5If
KYPNNXw8SiDcI72AnvldOW2uumAQRwcja9TXun8P6FjnpRI9g3jTmM2d+D1k9+bw
wK+Ib8uliHJtQnyHjc8+4dSZFgJgON9TgCjgruOViVA462rhHTjrOTuzLwtRFCz9
eMlCwMcZI0sZx3RC3f83lRhNwH/wDEKTyTHcnMA3qHmkUsobAZRu+H3OyiDeLi7H
mHKs+Q9UNYlf/xBXcifSMpIJf5o6H01LaxbvBvxvZVfSLTphw3j1r1cqiU4JbJUh
l3yVeCTd09rpF46ol9FI4k8nUWof6LJukP609aCzwkEXuYnBy07r7vH8JiDLhRkh
Qrbo6eJhGKgBao/v3f1wbLCeDmzgSby63utdKxCSP22YW2qP1TpppV4S0Mq1wBt8
2cGp4rK1y1zxKlxQ8+87YBGw7oeZWIklxwL6cVrkccPWRzw20dneSTJpsakBELXG
y7rFEmVQZXKB38SLPT6HqUOW+1SVQeGGzmzlYg45eeh16m/m++wiv80n4JpN2ZiY
2DMZqX3xKCEKr/pn6BsNcOXPXE2ERtT7cqTHbiUUbELUPCSYJSIFOjvqZEsyLPyp
qeDCUmBqIxJZ1fivkxxvPcfe2Cluyh2ImqufdffFCo5gQOl0Mlo6W7ECggelFI/R
OJUpDY0+csnf08VZt6uzxo/oH8HPRYyKK723dFSuevj/PtaSRKXXG5769E12lN0O
TI2Oh9K+h7UYX+sEW3xsBwg6lR2eQu6lsDKL/lLpFX7p3xtC/1sU32Vuc8Wy0Fjk
tu3cM+BOi3ThPJruw3QhTI1X8bBdXrMXDlz94OwDhMpMSmGgoZu6ExbftkSxwm9t
GHumBloiMqB6557Z+/wkGLb4xa6vanppuUhbhITX0OVthAdLr3GGtTB+qkb62phS
iS+CfY+Eja5oQbtlbQAeFDAqtvgl/dE4xdL8L21BY0ZKzKyuXXy3QLkMQ9geNr7e
2TTweaFLLZx3vWtPMpMKlQJBPWlaFLZ6sxYu/lwqBM06GISLbXYmFnQEYSoDBw77
GyGdRn3Fgx4pEdu8THv1K8/1S+sWMRmdgI9uaC+dagE8iUdt3zTdc87jY3t20KaR
GSIaSWaSWPgxwGp/3zLOoWcTqZRx/+KZm2t1LbQb79grPhF+HgvoIYW18BfxywMg
+n7li+BgRrxrMB7reutyHvjzuOUHbV+TMqlVsElV7eVciuu/1am65aiTApwD9Gyw
PvgPNit2y030VcqJxf22ph+1SPP/Q6DjKYDTO1Gat607WSiY3Q+7cnOSTEqtIUfv
HbXXGDMy2lBEmjUPya1uHPiWNsOQqWHXiDVdpQ6NjcrS0zYMl3b0Gr1RKt5d8aci
nkcEI44r/paZunC++Qdx1rXpQ+7oo2BdpDqVnWQfXcdSbfhq6JAhCpPdhN7opc/q
5EZi47ja4gNy7rd95sTVQfFXStijskrtJJE1LMhBNIWuWhdInSkoE8utb10QWqjl
nIoYdMjr1L/XG1P9dyXDVzlAetjpFTd01egYufzwKplbtX50ctcLnXft+H7ywR1H
MsSveayhn4AtN6eo14SRueyzT11/hVll9isahZL/Ht1frNag8e58N7P3oAE+QsH2
ut4VqK2hRU94t0nR7Nj7uHQKVgS1zLCiOCoh+GKUdTQ49GxMRscUfvNCU6WnXT0Z
k+HRuMMQTtToK9Qmm6+j4F+Gwc5nmws9BgoSqDgQ9+h64+Kats8qC11r6bi0JzlU
ejs/a7MGytmqfLtkP8Z+snBUdms00wzSFmIWg6PqdPAdGHRIVsPM14wOzZcjO4uz
HVPQ3sN01hWOv2oESOcFz4+juyZXKQ+7UwPWJ9wm2FaGhLpk42DovrzTKAxhRWaG
/5qyQJ2w7XlbuQXb+YqMOYUf8v6/3oEPPT8fj/kq3wO8SFQIGqAwkZ2FPByksvFY
qWWYBZlvT6VR0/x2qhK/RJOPX/9KARFMLtIiCL/d1NygjUR6Gv02awcIBe3gUFty
djlXtDLguZAbq5fc5Ictp9/S9Sv4CHTv+LnTkt5Sqd6cPDzdKEV+jov8RmxMXy8t
etbLwrEl3g29rnodd5VAdac66MTPjpRL2W6GOEyKAWGQsuR7GKUcv5YcUVyggnku
/njJvJ+XDSN9sYTWNSXVu/m3ULrztppu0getVU/t2H6iIpJ8Bvpp90USbF3xDq82
iwVwuf0GzByKSzSM+YbjzbK9vVSjQiIjYOBGE3bnZ44p0Gq0O2xofMxcdMhowEyg
PPjU04L6ydGesqu3dWCncnSg9IZlJgQ2g5opvTlx/jGT4iUYjElpNrBtxA2c1w46
PhtTXKj1NX+HunKuwAC2gHMpsPeIdEYtCJaYNHFePsEXIy+/VsYCbzqRgIjb3Ml1
TLosZxuKIYt+7+SPBsSOG4KT5q3Hq3Bn3t0LX+26Xe6dOdH0/5174WKevBi4lw5Y
hqa7ojkbNtR9hBN0KH6MkQOwz6iLZtMQZq55I/J31WJm08a8nDsCBc0Rw/JwVZ2W
CdeTa8kKx52K8XqQw8bYOxFKVgEjVYdl8TYUH9VpK5gjGeBdtUoWQm2O9EJEtNZo
f7VlbLIoo1O/+ZKoYbAKY0BmnwuHNin39gODiFXRvLQkk4LIB475pYygTdDSrvyj
ZhFedw/+Kkqw2CUeYiQQRwNGoTaGoKFk0fGJwiWpXIhZhKxD1n1ICidhtEB2MDij
U0uzqaGw0ZIvHK+OEVEe8nZ7NsDw4JO6q9iAJbVQzU/dVORZhO3LW6FNKScchRNC
Qtx0P1IdRnjzK+7O90Oqk7Kdxsx0U7fTRwwmVXX4jlVFYZ97fxbWO6sxGVZeq5CW
8qHKtyWIJF6fdYH0fesCYLwgq+enhn/3ml3CSkXBPC3P89f/QYFRU80deAB3kxlm
8unXKnlIos/DpKNdlu4V0DW1AK2p2rhh5WDwliLt2CL6sdn1GCkK4EPzeT7zQAHY
N7XAgb+G+3Hv1Fp79OpPN4hOGUxiaXI64jsgU9OCkLnpYU1kO1C2yxdwJfKq4Wxn
Y7OcKHUOMp+BCbYe9Q8IIISAKsLUHAVEywb01e8LVhqPvJns2GQRPaSrT52bc0cR
k2PfAPxS7yy111IrkyjLqL/tFvHP/TxbYxUXWF8Z2ifdlo9SM8h0K2h5UMTIJvPg
6/b3Y7Te4a1A8c65Ezc5qDrxDVyBJN8uuKJEcuhqgeqlMeDVLqpXAG/azCLviMEx
4NxLco16QoA0RKatDjvJS8ihGnM4v7Y6pfZuN9kLSryKaGelXUvlJ2yEpKvbCrJI
6PnxNEoVATSjVN+1Zd/4TdxT0FJx0KhzRYRdxUJ6uJnK8VWQJfY7DGFtaF6X+Ows
VJmvZeC2wzvKeWF8VxvUusjhEVSnf8EizJNi8j2JkoEoGRY3mmzS2yhekkNgnkT3
OXdYXstFN5pzNGQVCs7HleW1FEVidqbKb7H1vbU54s3k2E1RagpdiSP5H/I2CO7Z
RsbKmPzEwvPpPZIg0C91pajaZC/jLW8E64OmodfuyTuVEYCnGYJ7vBnbAsMBt6wm
F++D4X6k+gVxWBOnZ+vikKhbcNU7imR2acoy8TzYHlHhqPceKA5tWQFcDve7oKiZ
f5qXpOtwraUI0uBsqYpPmrm4LRH7Yeu47fenVnPUJi4kNFbCXE6EgMXzKMBjpO74
owqvKpEef3sleWlNafcxaIjqfc67fuojrqYO/FFbUYrWCq5lyG9nqJfAwD3gxD0T
W7CZj3mpvJufddxCzYlMR0F1lv7IehKxWe5y95DfGRavyIXImWEp2iUIPn+tndPd
7p+Wm0hb3PKrVEImxSrAKJGwFU91Os07Aww1GzRhVHjXwsNLOcup5ADf2IdQN3Ze
e0mcrB75B3cH/Mor2Uke9q6bCnEG93GBaH4AyuDsmClQlRqQqSi+hRY8eKTxsHCL
YSwCd8uL0FtuElzGal+neoq8yFaLWfEyAm5cww9GoRUBrLXxkNMhVOP6o28b+7Wh
qxrdwnw8x4Qri+85n65NoQLKLGNLtVp5SeAl6pG9aN5+lJ/6Sr6HZ6cY+jv5WSbW
FoO2SvcK33bd1yZsdayrJBo7FBSrvfx/TeieGDiJclprkKTntE5+Fj9hX4q56GfZ
bh84czK9XIHA8AZvyzVEBAt4kVLnyxhVF5G0p68Un3Mo+tc6XgXjXlD+73xoJvLz
YlFevsW+tr78tpV54oJZcNjfePhnAJaj+hgZXPrRka7e8q0eu8cXHyY6HvE2DfP8
U3+eIW9UkjJIo8Xx5VXBIZ80t67AaSZ16LWrlpBeMBT6FTnk0Vp2UXB9HeD5nCHj
TO2cZLHBVVsvM4BRyuB7NLDPjimeCKVrLjezgAy9ODo4mnLvwCzmBN26UYooo+tx
FnDxMz3mOYYJicEDhKmD35H7UdJaV9fG9rYG4WbXQUDG47t2MO3E4bRoXeNxe+hv
TjpBEzmCU3ZUnnotthTBFeX3k/jBrgkcUog0qZXDsFiQMweAEHBeI5MfdMC4W5X9
5niOrF7jd8OqLeWk8U4buDl/zBDiA8S4TxxeDOpSoADqRO0LPICnf36Dhv1HulrH
s15WngeNU1gheJu6LZM8RWzpwAJmQtpdTp/zCnSX7ZvA8NRGNKy9NXVsN9ZgHMaJ
VOPOg14M84rXGvzuyLr9ZW0mm63y3vWFs1mPsvdRoLb3mkZQoICbDOLW73CI5KBq
hY5nASDQ6fZgAmjZwprZ2/lCQ2E+db1/3rmNKXaY9rujT5ATMOjFxrTBNvjC5Uf2
ixuax7D7wKIf4bV+WvDtmeWa+jF0jmYsnVsVJE7qjDwCaBsPWmzgFoXZbsT9PR+9
vqbC6nJgPhwE6J0FUngcFeLirAe6Bp6uZsnGqPUc5qxwLR9A4odiO2SNELnErGAg
UAD22S6lJqS8xkcZ4LHGKQvdd+FwuIT2CXaQNRBoKROspuy44bd/z3VU3on8A9jZ
POV39ITDM5/8MRipdlXcuHgOBeRu3RJ2k0tHwDSssVN0voF8+F1bXQyviurjRZrL
nO12IKCFe5yH7s8jpD8wpM7wyeLY7GCbdKBl0HkdCXpaRvjrtERL0vXiSUEdnI2K
2WHdaBBkiFkPuPWCZTXd6sp2BOZ2XJDYeLuSYR4jigPUp/2rimrcqW+hSDFQ4LT1
5hiXF/zTVfcvKU1jKvDe2jBZeqg7hZQjyWjrai6qrHHtW3F9tIxKEzB+TrZ0MrXY
1UoQBXm78MGcFTQwivFut6Fvyq4O9v3HhK6F8zNgdMYlOkCdAfmdwJPpEKUAMRJE
QxwXrk3ChTrB3j57u/3Tf9kCTlM0z2hx80qgeRbVJGFDjSQXc6XeMoAoFZnVf50w
JbMWKasQmxDpZPtsd344molA6T+Pt9Xn/5oQCmvPlar2wgaPa97H40xybgMp/mtj
zZljQkJScXCaOKFq4PWJv8xZW+SAOD9oblW/sQgAjDtr3h+Njy3agBqHvPfW6DMR
+LkJx7fxOVqAuAxn4FLTyxuiK0o24daFBqdKnCdBHWVu30vQ41kxoicCVcKd8hBM
2SuLHUXTP5lPr+vOtRx9UWAMtnUs51F9tODjFe0A08rg4q6QWKVIeMVWSs7c1EgB
W0ADsQnjSn54Obgwi25hUyceM/rpPkiZzxv+YS5nsMvg3pq6/opMlc/JMw5L7/Cm
rechmoumu8nLxhOXDA+KXdQ7qO92c/JlhfJIMEjgNmtsw1AwF2TCHsO/Y5ltgf9l
sqvQ0J4l1GiIEsKUEVPL8vhxAkXBMMQdZaVrV5YM37Zw5XpFaTaQNcDmKbYhP+xd
bk+H6v6xzMS5IZAec5mJPCLbPRInaxLtnMmEBUDpiS+MFfi7aFrpEG9F0TY/gtFo
UDZN1V2DVdWrToObbo4BcJU4C01vSWIivTKPAhucJ/Ee0IdQvP2vwXXXmNC7lq/l
ezHzoMLCEjeI0Sk5DlmHA+HDRxVE0LJ1KhINgoIBwIyC2ieJJlzhKqkHXggKwPMb
8oIYpNnHLHSKRQsMYwQgdPoRISuu4VYLNwB/eP6oa71Oi6oXMrD/2x9pfEouZfU0
gZ6Rcdr6Kq/ai7hGPjKDBYgXYceQR69+G3BhF395uUZw47b/BmvZNEKTOQyh6SYZ
dquUx86nmZoBgghGPRqhrdZnZNMFPnxyX0JwDj8cS2iiTDBhNoDT6kHHyvruWmFm
uBpKzr8Gua1o8yOsFg7Rd/9AAMLKG2Lpfr5ofWocmPAdo3yhjzGuGDHl9Rnlvxmb
4B0eav6SkcrPIlJ5yb15r4EhdpZWsM0ecZNsdQHePY1CUJ7LZJXc8KgcEUcw+JHh
R8uWNpdld1wr45N+vTt69Ek3ZAXWoaRictiMAmtNmUEBxBpN37IOYsvxvOFU4gzi
s78V/QaT2PnflGZ/zad60WaiNcjsOp65CCG+bKzd5CU+ZT3GxZ2nk/PYHr4qjNWC
Vad6dJMm5tlKJKsJWlz9G+jQub3uVRko7leHawNHzpILyYK1Mi0q0d/rfd6FuanA
3KdGyvRifITAFdVw08flQQifzTi+IKigxjwMVA4yYbH9uGqJC8w/zhNUZ3frIIfY
yYBgj0tVFBW0Tv0rG6WLlti9zj4csmGB1b16hLjhn9wsEgzXlkQ+WMmUDb/ZzK64
QDvpA0lMrNfftkHO0H5c+vrxrSQqHUZo0qebZ8O604DnxpRWAsrm6td5R6p73e4T
I7DuN4VZrvpMOzsx/Nj25bjyNOHMDLUXMCY5n8mvCCFQHnC1jSuBKsrrqGjr29Zm
3NIUwf4dRIfA8r4Q2EoKmMZL2YKb34U0ukB1acSeG2cLZ/YPTAaWIWmv1mIGdvz5
sc5F6jJnTq8XlAGvkjOXSd/grBo1Z+GBj9FjYJLjEQrj+bixVcPyD47e8rsmFkDL
QIESJ9msyywbYcfGHu3/Y2YLg4/Y3bnY6iQT8GZIRg3YZyTd9uzQpXnoJqu5l8Bt
FGNAqv2HCtm8y68G4Xlh4K6I6cctuD/VzuY1iT/KSFUoV22YFVdPSZYpRxLgAvTr
xDOvuK1EX4fY2NxLG8ut9kfeWYCMOt5vFLPxom+6bsizVfjkYEuxGmm/w3HWh5Ze
ubpToTdCvBllmXc+Jm0jgjHzj/d3tgl0ADpL5J5RgFGvF/Gbwrt95JceNwAMrG8e
zST10aOIGdWXO5K6BlZxNOAaaJT4/tO77iW/4Ccf8rdhsdRX7UJsy/klc4z0wRy8
VxM1zVf+hZ1xzPLgfUOw/suCmEJ5eymsGvzHuQdSycqBKaF/Pvl71bzyYDWaSyqN
BTMUhPJNOUExsXHJJZSxTPlm0KiSmiBB5KHUAE+GrXpL6DsvxcAU8rOn/V2jhBep
gvp8q9hsA5vRnz+HwPzvznCrEyVF0CXBuzK33Czd7kBksJVGtkI2+0pzIuPR1kH8
xh2jDThhMEX4BN0EBDKZPalu/ocdS7EA9iUEmX8iBhzO4N9PJ+5liONbPJn7EBNX
m5D1ePP1mphbo6rVdC3k/fjeUUuy5se0fIn8ynHIww+97by4BM3xkEJde8FFEIT1
OR8yBxZAlnKSGGAVHlOtJ3Gnd+qYdDmchN8Ov7EdJ9/v/A7b7htg0tDultgcbBEU
Um90C/aYTYQCNeNYa/D+PAjTRVpLrpnxDrE85K7X73PWc+YBB7iXSYwxVjCKIhMs
OY3qaqxHujY1yfctPoELfMJ5hKVtdP8uElGvt7MH3fIrjkVSFDo9WtSvle7vFrrD
DSbPBVaDl+9hatfyQ5sQmgg4d3RkubxWS9pxc9s6xOP6KCDVVHm7Gi7G4icVbV9O
KYv7t2k11Na20q+GrMBZRT8ByLTJGSFj7oLmNWFJm2eTfNdVhcZoxepBNsDCSjA1
2AcOCirtw9F8pQHvFhkW7o2QmJ4eDe8f78Fk394L5VfPe61csotlzvig/10xTRjj
bwZjPohKtfU4d+CKj1kn2X1pILovshGtSXH3klHM5dGAHAITeJVI5fOcDIzyUnMn
8EfZq5eJ+NE2c8tJZEwFN6u4NuA9i6+kRl+ji2nobM95wvSpUVAhQLwzqqjte9aA
n6pNg6cHKwyQ2o3ZQF84Y5MeeuWLQNeJxbbw9RmjXFt59qDFjM4mIwUOmSYPPpDA
NtrHbxA07R6jSGOgjiAbK/Vyt8tkGcz8TY09UP1rHcdv/v4KZ2SGOEglP8VlrZik
gL4g+P1elxsYLz7fAWbDt/Zx6O+CjjFng9dIQXvMeZXvvADKgCZlHTAU8aEKphzK
5kDy7bwbgaDHEoFzrBIZHXUhAzqZT6+4r3I2Bg8Ork3XiAbL2myeoAnhftnh8N/8
CYZlWjYy+3t/EjOVtwMmfggGhUBNQsnDcV1ssVSOKE5OUXE0J0qSIbQMrMG412ux
LCxXCw9Pe3IUdeKzlq/BGI3rnVZqe28yLNsv+9U7Ugesrps0uyHEdIqu+9cPc4Oj
EDvzC5IG9mWpodNAHFSgbKSJ06hs7ljnbOfkXCmUYZ/lg1Mi8fTwlzCPeYetfS6I
uZ2xs69aYROLvx/TBgptwuDBKz7B0ZTG60KZpHfMADus3lPoRPijWW0jLPfMuTFl
mIViLxgs8rUgSzqvhBtj+iwlp/qbyIJmPdH52YxavLZ2TluyINDMmJS6JBg2Q3Cb
shKolUjyIBy+1sA8ttU4jPBWLp8d4ZUF79WAbIbRmWUr76c9mZoQJ0zY5Iol9Adq
qaW+yBgMCzl5rn5An4kEwThZLk8kp/OCNBlMUXAJmNITIGdm80V1yh5j1YI5wMAY
xcItK/4Izos0M7arnbv5H7WULOE4TQOpVUVWWkzSiFx0WNThKk68dVIWiMwgEmLi
6aDjrrpLNO5m9OY8+RBhIzjlvDnI3Ee4pb6WhU5vq8ks5VpX2SUhh6UPEudSv/YD
KrJXqoHJw+auBqm7ObCnElmYb0e0WcTQxhra/q9H1xdoVmlyItF1iykY1IoloC61
Fqbpa8lv5+h4XtMqydGMcS48y6XEInwWzrgF4J4/Estcbseya1vR+IhpMNjpctVL
OlTgjTSx/8A4eilHiRITdijjOhwQo7o0DStH+mz9iSbRIZ0/rmtjy5FSM3HR4FUO
q8jquzb8sy9ub/JhCcbqTwh0hKdDCGMrPnEK3ulUSYuEpdG9yKw1ELg1UUBYHtQy
unJvFCptHZHOBNGM5rSdqMTHI/JFkmKewjJ0l8N+dGAxfUXhxB0Up9zueZOYNCAX
ta0mCN6+xMStIQBWNVNkxv1XOEQmVEoIBINU16a/4gmen40OnaERH6YODwSi2rjj
lb9RvKBZ3CIOhWByM5Oy6kV0VGDzxd+kr1WWKhOZXbmzDwGZWAz7qVfS5LOn8YAw
CW1F8gT8HimEcFBvvOmXBnWNB3HLhPEw/tv5AkwU3TGhlwGzpTYNHghVyNwvHFRV
ExNoi7OwOEyqcv3aUJW4E1eKmlHUilB1tfA55HROFCbuo2ZYXMAhxIr0Nzu4lwio
uQZxx9fPswp9yrdFP/+lGcic4pFLlh/vipVpjVt/pU2HtTuowZPinstG50PsSJOD
aRfDuDfLoT7rk2J99M3kBuSvXpMtwfbQyIxJJq7k93rBUscLOw8rfSacRhGMr1Cl
Nbz2YmSM7FMbEgJ75ZHaaZ2DxPFTUt5eLjtT7QR0cHKmYioNmjXVRBdo1PvKFUZL
Pn9PSa97GvZraS5mbcN+TKSU/vO02ewrVgDxpy7mTXcjPO6KY4fOux0oB5MC2mdm
88L606xCgO91qZCnJIYfsDUKJnxMe/824y84lZyKHKVR2wscTOHsz/iI8aLJwNuD
t6MVi2oXufEV17p/DgFurkvE9qUmKmGXdRh6v/hnHrThtHybI2VcCxMt0HiS6AYo
fq1GXi+1/JgaTbjtvnJiorclSF4GTXn14O3aCbftJaQm8br/xViBqQ2ikPTaIW/W
G73Gjp2cSnc2OuHv6uo6u0xIWhD2dcJsoD+bpZSTO+OmkBlk3ssVFb0yV/jE9sWL
x6mmxTia3FuE8Zi6gBcrar5UUjREPF+Hntoi7qy8KY+SjsCN/dNU3ktxFMy6tNnG
4vKw8eRHyZzLWJQHqVzjkz847XxkaYvhoX3ivJj5cFv7Tm4AbyjnxTHiRPOdqrnH
8Et1T+hOxr02WiFyOI11TNREwOrnPJ+uFwiIHkDlhDQfWBrKJrkWXNQBdLotuau2
F7kAq/FKkZL/3GggiWfJUZ/BovQD+jAnUJePUNhqnmWgiWa44V9AeM4O99itBKJl
oFszdrI2m//xWBPqIdzl1ehn+t/y0HTO0axSsXvq21joA/rpHpnOuMyS2PXHkf6+
H7yDRNUXCMEHsye6qb6KABJj/CTXaTQEdyjU28IpFj0itVNEGtqRUB265nlBAnUW
GfUBgqzKnjxXNMX57xIqVZrxmBnIkWE0yCK5XtSFcskMmzwWSBU3MLNN0AM8eAOs
dk3gxniMXaavq00JNV1mmBq+utYYY2MoXpaNSa+JZsgtRxjyr/GjdwRaPRLUpTZC
oGgvpT3IjRZP5p/YcSpGFLDy1tPU7sTR9QsYcj7PW8K/wy2Q/P4VULtaRRfSVIFd
UOxT/Zk5etV99fJGxGGzuZV2+279yu/T7RoXUZh2ZYirfdjeMR9GnpkqSCLzCRCc
JYe+6galcKSD7TzdGn5ADuvSYs/jGoDtT7xaZPvPKztOOIbVkMSQiiu3POh+uL0T
n8MLlFrkDZGmk273C+46hmMrmkLaWVp/GJ/aFRjpGhW+bO8u8w0slEFzOlycv9R6
qPN07/eoyQsnfV2DUWxq7fO/G6CA1SEASmNb0AL5iTv/qA5eg/mOoov0TDANcLgu
T2CFp6dwpZuWGnjkT6MWEnvkwmUxGsVk4HO6PW2SHAZ7FC6kI620dbhjdUt05ZOV
h1io3Jge49s1mNRCnbsQCvE7weReRq0VizSgSC6lFLz7Y8ECuryN0QBat7b0qHyg
GkIi6H15Kid1le1cJZph2fmR1SbINquaiUvWSQtM4DGgf4qgjwqRcMAr2nY94ksZ
nXtmz6VDSowW9bBOeNzdA/d3NHl4X6m2bWXXis+6d/gHpnR9mhQTFj+Q/cQ28YNj
J5rWvm3awtrfQD2aTueeTof+onjqmJSBfwEJNlysY6Prod1LEZ/IWeq9fkykHxP8
OvLrRZuZzPwJEWZITWgeXRen5yAY/jvXzefCiwMxoWf9XMYtTSkUJiZ4P6OB2GY9
/3fC+D0GGLhVX4FifYmlZNM6e44EB+xw3J9YJ6TsB68HrlYK4P4n3AvtKoYG7px0
UNIpdvU4L7TlCLjGt2h+ryndds+/hwFaMoJZWXxj3k2EWcn2S0xmt5RgbALZNS6I
1pqQKSX83jOmLBxLJYN2bUTFcuR/by87Z9rNyT7dt5vy0mdwiGGwMDEDQkM34J/l
JjM7rztyFkFc41iZTjz5GOsPaO/9b+TleyOvKGJWKbUzXGVl4+tLmJQzh+Ltr+7r
bkHyqDWE00AeW2MtM4uHdpGG3bLIssntKBXQ7NH3Nv13sq+0zGjawMdgfQHgyGdq
+/Mja7MU8H/hZ6kAaQsJZ4mzT8JXsTe5YhnVh9Cu55678mmAiek7h1nd0sqx4Qv+
QLSaMLm4i67JMB9G4R8QgX8vvEAwK1gYJ8ZKMkFQZ4Y3CNz+NE39Ro/QFBsc7dru
8UUKVr8B7jBLwr/KPO5GRDHcluZIOtsLFkkmpV7bbzyXkGZXdpU4LB7WvaYTA0Rs
1GbfkvpJS5hM0QPxSH4bU/c2N/vZwHSNuV2g89io1nT5TlMbCC9EpEozHoHnnixv
8Ydfsd6hnaSkYt5EUpVN7rjIkfionQtcbkynWC/ljqMNY73dBZ2vS79cnZ0Cra7n
aIdkR1eNbbBjKPAvTuTX6jN2IdlGGxuxDF2fAsJwMPJL1omRlnH10d4BLxDuhgK+
Aa/Vgjt/CB5oEb008d1JInBjLQ99v+LhqgGyIETMltH5Qn7n6oqdRXKIr+3uapTx
McpBZlaluP7O1e/yMW0SOnMV9bh8jf63HLxMByOQM7Vha0ZMPZcYWL1D+neNlJqW
QHbQGmNCqBjZNAxoEANgKj3QPBgS8p0H6puyrwvUNBdG0uxstf7+433gNIzqDJ5b
Rd1f9FlV8WlGSwe5NoAC31Ogee3HZFGkunaROcTYe6HmI+FS70B7Vo4+Ai+rSdbo
Bp6OL41+oye2NMZ4wbAom96laouMn1P8yfyjsdFpjqFKunmFnJ6RCUHPMPu+2xfD
f6vot+6yMI2nLm645NlVvP0TG0JQPAFkci5WLtYEDsTxppvjZjdrhyZmkTi5epOO
x+EytnlxL6cmeOfshIZ9xR4fbku8Wp2sVMNfrphoGZtMz5yPppAyHu8E1aEMx/h7
ihB/sS5i8NysQZaN5q3Xzx3ylxI+ZVOKKRwrrbqAhRcAP6JifwHW7uzd1bUTDDJk
ulUGbZrdgQgGvm1+9FeFVuG4oIRR33pirCpc+Uznmf3bUL+lV2XdWKnb79e1npru
dkZBT9oVfWIKsbhxjTN7IhELaP4aiS0okR+HbPQEsJgTd6nHmeVXq4stLQnfXLDd
D28GUojT8hwu0lG1FY9ZjXiBtDpM3cKYiZbOwU1uk6LdV9oK/osmCNgS5cxDoAhO
5qUIQVGM7Te8WWKDo+dEhNbIsAC9m/pm1TNygNHiHIkl99xIQj450UzurUg5Zxo1
ZqLUndocYFvU3L5ayHtC+7ex3oXPkVKFY/XxSQY4Ej/Dw+H/ynIHogLqY1tHjeI7
ofKb5PZyPE5WYj4rYlSM7ahtSpW7CrARYd+gONp69HgkClHCfnVjZ6XcR+Due4ky
COqHV5ugmrwEYrSysuB4FjvTlK4dI8O8h5EKYFikfugaWfg42IuG2+j7mF5BnXPB
jos7eELIqcKu7hGWhgUpQwHojoPWMP9E9+MPGDG/QTbFqOJ1M/z6lQYckKziUOcW
Bjlg9U8xPoGVUfHkMU8UVXT/ynvkllHdZdyz+KeBtjI/DAE3LsTssTjv0k9u9NHu
8DBd8nkcQxFpPMWbE91T6yymdXURJpnVhsVM84NUxHvlh76AndHB6xCZKGW9NHiz
YNCGRWoVOx/H0qcE6gGneikj4dI0wsL19hEQRef/dILyXJixpUrPcpXWeAfgt+hm
1mo3Mt0nwZ3O6Ft06IqKlvZPhMBlJM0b75HwOyZaarmJl1uqgivcrMjRRHvDk++H
vo1BN2125s0xT2ZMuYc2nJ8VbVudM/phmsQIHDO+B9crZrC71GTeb4IvrekFc+QD
54xNIu0i5ifWu1pk6icXkLKyJB4shj6gbPMih2KelOP7FcvgLOoD9C2sCO3MZwcn
CJokKoCNC1tSKSBBuDoV/sabQ1cGu3Uu/6I3k9S9kRyde7OiVOXDWH0zEx4MOPSh
GoOw0cwleSoD0xljxo7n6IOpyrGom2xjjdGteSF/b3JgrihoYvVhB9omIfhTSCrR
FdSiXDw/uOP3UVe1CVVklYrB1Ro5JEISdokyDLHK1136Spc4xibExtFElfJQeU40
C7AMCgWVfdhpoGMmb8TshPcS4piFi4mbFZ6CKeokSSKNedXxW4RAY7l8/rp2wlkC
4YKMp3l+0n/kgHC1wFRLRZmQ1Zs5klI8Jm+RJMPdVfRBqgF7Zx8lZUsfaPjxJgK9
YSy2VR/L9G6IrdwBue0Fr6HxB9zJlYh626m/0SACKeVntCYD9Z1AyH22LhphsStO
q6aXRtVClb0nfGP/PnX/j8mNEqpznaop7nQvxXYtDtXGeEy6nHWxkPnUagnJOfhQ
dVD/dlzdCQ52WzbkZGNXQd1fA7pCs37Y1eiD9OU3NAg3VaBciyM/xa6QtPdwcOad
5b/bfny0ZaUjM72oKS0aHBOXxzzntgzMQOCVR/T5lNACCkY+pjajSYVOJv6OSXjr
E2Dc5ACDe2goxHqCZey6Qm+kPviyNQnJZ8R38r3ABaSEGHat5YNkWhk/G/EgQO07
DGTzlmyAEpWiaDnMsHgBgvapgda79hRwUaevRSIUJwJewJy83o+Js4JPl0CqUs5A
xx0RPwcb9p2SXmZYAw1iXDaHro9I/7ZL/AMdfAYbROvcS/hz8d2kcxuX69PTNTb9
AJ9xNQYTA0r01jeaMwWb2xX56ijOM3AKiLCIpYfkRLswjsuW4Tuw2BhqD5E+uSPZ
4p+zvw0Hbow9AolL3Abv3T9+zPloS80Bts5IzcClIq1oqNAhtF+cF3bvLpybjBZL
UWZZaprfl/pW3MrWnsna7qb8HOKQHqbzjZk/bdGVHzs6rIka1jlCQs8aYt9FlXU9
rvlBOeT8o2GYvbQF0UD8NcRR2leZixeye9KWoRr+KWDgzh+96xiR44fWkGky/UJR
s2r6qljIV2HiGYZFlzEGfgOTHc/SRmO3B43JZSwaMUx4bmr6a8ltmu8HXOBSYkRu
MyNkDBbyFOq7joe/hE2lAcft6GBB7MXtk09iSVfP3Fay1JXuyQmRycueTBKyUkO0
q0j+mJbl382isaXnUoVFSxHRI3pbnWP+adrVWzcLHDW8AKLrNiJZRxVen48/jPzB
UE8T4zPbpziIkSl+6EKOrqYHmFj95RY0g6HINB1O4cYN5Y3haHtfZe73e8bK5Gvp
ISJr/iBh6lTj9BsOqQjWS3dEfvgKcKOBvQHXoylKmigs0Cxgx16UHhIrGa4vNDD+
CRaS2AHD1mDDDycqL7SLSw/qlhORfG7YQU1PRqdZriPj+2cc9sdNUsmZ5QHxE9On
4vNN/ZvkA0YEN3RPuU4EcupXuiwlB7yNekDe/xXTvC3ef2pTfiKjJOi2Qs6t4EhK
F0vyaaF7p2+NHuENvZ30i+ygsQkoW0uAfc1GUoHKw1PCT5NpG3ivOwwZw3L7j1b4
O3G7V8YRY5EeOD4fPFbSfcgFznz1YDytBcP9zk+Przvg+SsTIJSXUn0RVrVSByZ3
NUwNX5eUBpOz4b9iHcPXLB5g2owd5DcFai5qtMlyg0yDl2hZ1HAweoFEjEwTfrG4
b5RVijEaS6ZwCBy6v3gBygawUbD1SHDFVO188YmTgxQParmNsQtlHl3WcM9rV82W
2yV9b0amQ4kRAlle4zpGZdsXx6W6lfHEmZmcEJzODaDJoE0SyjuX7gat8y4GzRgN
8HjjBfCnFL9XBJgwN1WpIT/fpgSDp1mABrEPgcHQ1XuYRshIaCEO+Run+bLLe8IW
ZSuYhcBwylGDawXTArh6XUGtH3IcY0H/YmYL/PbrPgKlG0yTFpJCIynA8Kz+1SMU
HJbersEeMZeV5Ahwqq6U/MHnIg3QTcD7vgm4l6ViLhz/VnwXqdcuhyEbx5xgr762
YbYeW4DvCJy/VxMk4Zh7EYmicPy9naEAGOpMSRDOzXAt5cwd878WKW6in5EuviiM
1atC7MNjZQ5Yi9a2KYAlD9dWFTM1M1Jc8Nx3/8QU8Qn1hk1G04r8dyBKUu294pVo
ILVzi/5VpYhpGmrnbHoNJTmwU2vjHHnZBFeznCr0HtcIl7YTaR9d2uswL00AXU5a
9qO/J1sII7X5TgpfOdxLfAzTuGJQZzN5UGhfSYOX39MO6Q17C3TxhB93yrxBWIqC
v7FYWvW6zNWeRcksGQwN5ZrQDK1+cAKczEebASDmojhRhjvFu1QcIGpS9Bn+N2xP
XMFnJ97RjcytuqRqizRF4BkcM5yBFXbDABLuEE0ZrQsr6Zhhwc9PTPrR+JewoPdl
z3OuvxTLr5elKhDEK2jsbDunEUdHeARhDdKa0+NN8fdHtd2mHY+HRJUYO9F9qfqV
oe9v9guroZCOYSIHjdrGECYg1qq6uCagBuS88FaM/fIFwfZR4lb6g5PI1dj32o08
hiJ3YE+jCkWKh4/bjz71H0u/2d9dXexKPox8w5/LbZfaQM00FZzzqHduuqh0xszg
mCEJ5lSQeFEFRFYecZB4QDC3lOvYqOu6q6/HzdSNN0DjntwHx91QeXiRGYdv7Jfb
h7sY0HUq0Zq5u6mI3fVjEMuL73LRe2PxX3/MAOktiptp7bsrQozcLXRqaag+EkBb
iuuPp0UiYUh6dOaXaEsf3aLgEREKjZ3205AAtQ0bTzhtXh+uhvPCTa9kpzbWx2xU
SOc652xXnqDJ0aPhGE2byMsAG4WGKbeNVKRJ3o9jns2jYqta2ga9gK0FXSgMNCP3
Tldss+69B/OFXOpZvBUjRuMXpge5yJSJ5kJdlwgDiAmNWXBSXYIP9R1CEvd/pv5A
RxTMcR5rCZdHk5RvF0STnrv1XnYq1gz86F++DKywJkSqNTU714mBUEIi1W1AmgmW
921mDuRsob+fg72dMDADrZvwLHO5Vvk0a/c7oM4ixL88/HwWLkKk0jV+Ob4ys0cO
XcOg21FW81TLOH+NWvMLWetyIPJvPGD4MY3FsTCqRLdjxnYtlZFhYYbsuKS7GG0+
HfOnM6wOWct2CEcBu2EuEDvMR1hc60T57krATpikjBuMws6gFof5dqzK2bTs486Z
Wkb15SzGfQYa80CjW3aZTbACzNjkviAWBDw7hKLq2ZQLxSDEs+l+zozgGiOyJOpu
HNHR4EcUeQbGxNvaBjFHvs0k6b2/rcPq2tB52nDezk1/zuOcX+UO2bdRX/P4C5t2
33k+jBxL1SdSbfd5uBrvnyuhFvyM0UJ2JGsIjK2r4f8qfeyog7ZytAgKlLdljnS7
MBsoWFKfTHzs83TD2NlkWwFXO0SiiVgwAxTDgeoOjUYXjznZCNYEI/VPJn22xBmr
qOg+sfKv3AdF+4FoMDj7f62pZUOZ2Hx8kStx4JDDfo+m0RGU1vnk3M0j2mDZME8e
YnYqhgfadMwojnF7k7MKKeme6rpUvyZc/SIh0ICim1VgzqexnX89e+kspPt3Ogab
44Qi+PD4YThhF1pV3AsXMEByaxy0G1R74j/2YFvp3friP173l3NIEmuseiPFtaT7
0A9KaMTnQS7D6qcp8DJp6Kv15E03qJW1rUtS3aHXgvObwcYTWw1tC2+4Wzxyd//f
+FuIsFMd1UlAnFAQZKhoXGgIuzMv2ZzQeUJFdLppy18G2BqQjSId5Q3Z29gASEDl
lt5+JlTsP6D4rDIBci1Z5sPbOF8360PGZGU6q/zO+ye6vAmAEh9uAR7b4pI8lig+
I4dNYI+YGu3BzZGRDpoNAcbOOIembbr/QjMyXVmxDZelrMO3M/u3oMM+Pwm3N8M3
ZjBMyNuXPwSFWs8n8N86gxNPa9gUtAT/bBk9R57D700AHvDiBDYfx/Zohl8O1zuz
EpjLdJBFYwDmKURWMwwYh4cNRtCc6QBSBvPNZ3KgWfjDDtmZK8bJ3RVFYcwYOWyl
/+YhjYhRu4+IxcXh6BJGp7yNjEXcfSngzPJhyb+uw8W2HTSJprc5nRJtcggLHTwd
4kViedJijuVd7WHSXJYQ5Ik8cK1vq11mbyAMTPTd3YaR5QYnxtKU9m+Ojz71Z3PL
UkaBgOQ77WhMJAitpPvcDw+I6ilC3Dq0rX/q+tzahWa0KfOwQLRDqZGv6E8LDaIX
fc6kczVmbSm0Nuv3hFTXruiYOBEybKr2oiCJqhELXRz3LAem44k0eBAuosbZTv8e
w370nstESZtpYZcQf30t+kLcw/g6ECb6jYfcpckXruI3PIZTMh2f0vM7kR/yTOt+
H5l5MACaNRH/S3H9Zy6TKjzak9rkxnEeMuFTFE2B7ypdqVJyeRSnChHEc5aE3+wQ
DFU5sh35+lHhituyctc4s4Cg688LrUXTlBeBzMePa7uiLmrRc2uQ+rmaINzJIyNo
RPhhRZzRMkFxTKn+7m/LkArregaCN/KKuglXPTft4drGkS3WAQ1APlBwtndsq99h
01yXZuufsp3X/RyMIrPQSrNglq87SetkNUnQI4XjzJ66jg+5EAWFEeDL88VjA0Ml
pGhsxmL1rtMg1Z2Ay+iW6UlpWcsCSGfAKWTR4/Fg4XYqRkzijbWrU2IWmQim/ccv
1V6+ooXO7z2oLIfw8leVsjwpVehpAMusQ62Z5TUHH1at1XbCfab2ZWEpVdY3eABU
kfGGqSVkMjDQzTjXkn/OJ8JGjgLFjPm5yquHFwI/Gnt1z8Tj0yVcK0ZJLmsX3KrO
ADYITWbC0Efjw5ZKWsjvrgNTLsuZJBtNM7HG2vHdNDOZiRG+Ym9baRJ2sLJ6wpqd
7gyaSROHULXqfBsaJUU6R54j6ZXP0+UPtsIRKxP+Uk8gW3oQIX6wwJLrxqMXz8qc
uoq6AJagqPM03ymCrIhq48FSwpoKBm+CH1KoEmEWGGy47nLgb1NrmR12/PRJUJap
HdqUbl24PJMQPgDYDBKcMLBUuaYx8K5hkRlyanwiK+jH27jpjbpU4+8iIAO+X81q
P9K9aqLnmsDVI0ofWVn+fnHAedKjdvGp7qWzUyU8NCFD8zrmf6UOaiX1ZrssljTv
pXBFecxhx21H/G5F27ymw93RSo70v1St708dUMx6FK0xnPrbYuhHRPyeisVKmV66
+ao/0FV4qbbFJXQLTWDjpm6poY9lqmVOrzLFkpClwY0nhrMWSYBS7bVLF1pwsOQB
0Zn89AoQXiI4lBnfmW6Tsgs8Kbreo8haTfo1KlTn1ZPQTh00+/um6UipoQb1iimO
85ERZHxDBtdQN8y3EWIXf4CAz4QNzWe86CwzaLL5AvxML+XZybE4LgVSmeFmkwPL
USjZYsyWyX0/kJPJ+GqZFHSBtyFzUYUxY5Ghi1p8GUVqjlsNDvZ9NPDgqcIdmbd0
ny8P1qhC9EO8WKgV13/3hcg7097ZQcj+L+LitIxnyTdwY94Cg9XNpw8Ssq2l8Kmj
1cxG9T4/Sr0iSMR73wMEWv/ao7XCJWNgIYV0RBvxGYrNdu2c3DzEvcmQHZhtVc6U
9a/EoGFuDV67cnQRlSsHX8Oy++I15Pxtg0GGnfpTyOlcG753NRVLXA5xEj80rPTQ
qAcUWvQGYpxlGFuFzbiZE+26ooDsWF/aXHI5Utd7+I4lFXx4jx8msN7qwOEfiugu
p4Ak7gpUJU/hXu3HfJQL3m4iBaRwPR2rLBWo3y6J4tF54WFQDwf+lh/WqystxKiy
T3Bn4SgckLT6iWEqiTm4i4I5R62zEMu6qmDcej1/DOKIOC7cwc/rlkDGUBzwQzbm
CAPkSwpoib6s05Y87ca5deeV/xLHYZV73quH5OsZf6k8tondiikp6t0an+IoKeUb
Dv5pJBcCfUzt0mg8PAn1CelK9bJSgbImIdD6SgzTjRLbpSWe1WSwit9fXGzJOqD5
f7wS9Apjp6imzAZ/d7LtIuC6Mm4ef0MOwTFm15y+G3LLcyv06nDRrMkL4FNzBWes
waBYfwzTDAjMXsJqTrxIn2KK6m6+D9iBiqEUhP1V6iBl8UFFatjEafFI7LnF/39Y
VkFh37xl3NYo86t+mx3g/4h6RNw+Z2lznu/s/Ter4tPGDeH8Vi31K00Jm/YkEBmV
InXdkQq2RLRP3YJ3p7Tc3YMNb/uvSQ/d607t6kUr1Gu7GJ8OtNw7FW9qnQoq8tLu
7db+IA5qBO7tUa4vBK9qTw5U5Qohfnfb5hRrHudLP/aB7jSuSCZSQQ+t6wUxz4MJ
YghJRyiRn0C8bR5STRVi4K8pBGZuSClATB9UDSMAyPoIfQ25jHZftmtpm/lBmQC5
EkMTSH2aynv6ULcrLqweFvF0zAaOAcNH2WYFO41K+SYj6KZkE2rkrPb3UNMfWMf4
m6Dql7dBZEmETHVj975vxmfdrVeoTIoN9LYGm2JLmdu5xT7W6Jr1Xu5N4KA2Cvzg
GiXXBIuu0EGL2LpiX+yMCjsrDNeS7Db14Fy/GIjYriYjX/f6moTrq4P1oJ4v2FLS
PfYmwr5QARvu2jtnrmfkArbv7A+qryaQ2zqpZq+FZsId5JLe/XtE4RweSvFUrNpk
Y4EWQ4iAWhw1e3Rdl1RWNF2VZmKuCrIFOpdJwcvzoRGQ3ecJIzbU/cRJGdDDI3Ii
ttGYQopEYQ57VDWjZpqO16hToOY8Y+XzeTL0odDpLWBA0ym3Z9S23SVA1xC4av8F
LNW4jx0lykVYAM9rqCwQhgEfAHflgSf076onKelY+Cb3DTzBVYLarazwfXsLjdIR
bffjM12Jdi/ZwXN//ftqVF4yG0qQBOxmnkqywcWgML68CMl4fMMnAc5OhcUE9dvi
s6qiokL7Kkc/6/0bmOZyrvLbVcv2cZPd3dNaWYHmioudYC4h3jSVLja68rx42HSu
KxoX3G/Apn0V5yaqKgbACv7cgwTQYpeMakjINeQGqz2zMpwuySIJOUtjNpcNetpR
bNgdUvzaOM+wlmRu0hvM11Ra43k16C+AtGM9zZPpfmcwQddEvW+GvGSnvDKRjKQV
x9yjICWMIJQ4X2X/f4NuaJNbrZY/jLiWm3Jaf8rtpDJli9fvEVkKlLCtm78Qv+Gq
PA/nPlZOfzjwqycfX9zkQBt0Xtj+8RgYZIylqxWi0klxPO9B1mXWPp70/YCfoJmC
noXPP9vYMuDuEVEsGYpYgTDgpfQhAWtnqZIxgBArNjJqams959qBNbTtY8MiLgau
W5lPPVVpCDx6KeaHVDEkWGqXtbQJxdG9Uhxi8TiUxhyHemo/h+SQs79r34+c+Mir
TwArztkb807q8liEyytXnpRIjy5L/unrvVaTTaasePoVBMZaTxEqUxFj22GXJimz
kBIXL0PV0U18k2QZKwCnzSbtv+7D47CeRamIWq5J/DqiAoHztvFlTny0bLFDUDg1
xVqdfvd28O1Kw4req0YjXu4utZOXXnHHXB4NbqTCbP6ASwjybkHWTt/QTvrSgyq4
h53UDPEpWN8/2QNFGJ2eRxjP3ScISoEuf/HqQAPj1ueRPKVf7yj6ggddQ2pnFnsP
F+UyCgvx8lFKDWB6EaWKnPBSwe/zUCX/wuOHd9gEkeqQThEYxiFOmZ9f3LKwYQpr
v//Ht6+sVNbY8G7exkgUqB3ymYI0V/vN07iLm5XQHyPjOxxeedi4a/cpd8OmCdQI
mUU0f5CsKCRGWWbMvPV2jJXtUyqMB3ibtUN7t8SBcAuMhWJnomglJzNQBL46vVSO
HOwrfBSbtQTpEejRvVyV44BcLEEsjDiNbbCTVtegJPd+WPjWBUE+FNVUc/y59iZv
G5TEFA5Z1UMz1/hCeSkw+dxqKFYJ475ETmZFeXGujWRDZbkawexhY7MXnx0rnDTo
cWA838R/INrH3qeQTj9G4DpCeY236XhUYP9J1SNgZVYRAVnfhbdLMjDlWaBJ7bgc
V18b3sSkUdajU/EcDuBJa1RXaU9VNplMxsejiyUzn8kTZohdZiS4hHmwi0wjnfmc
TSZSu8F50h9xWuf9tSLq171FYs57DJNZ0TCWYTOZvhvDxJmjbDwd6P7UOiuoQw2r
pk4u2LMztRYVjUNg1d+fFfCrlRAyMC1fo21IrhrhO57tNzBK49golp1/ESViQ3N5
uF9Z2OjZRqPDHKLXWTSYUFJmWlXQzLRJLMXu4yurtlfsz043euC0Eda+LOp+HMSf
z+/05HZKdHZbhADSdgqBluyi8drD4I+xO6pII34+4n9Bm4g/FZsUwNRMTdZ+n6F9
kTn4paBz1PCm9VF7VBNLhCogEicd4jzOrOprbvL/c1prxbsZOJwo1q5d0FFL8RxM
0YJpzP1k78ShKSnFHOsJ+uJoE2S7TfdstV+xI5rQX7NmNbIhANtgF8j5+Z37j+8I
ZU3NH3ZF3oWkwRTdvduroglFYOdOhuOWjnOsX/KQfdmVK6VCuZ8M+thUV09QTwc3
Fo+Y6cOZ6KYHxlZPDUxfeiJbEfX2Em6KB8LoBD0bRijaq2IvkS+QwZ+/Ocwirc05
QCnwsgv7OnKe0misHn0lq2Vo27C3uo+VHV4o7m+XwksBZPy9fji1+iuu2UplZSR2
wwYmdwsyb12SVQVf/9jtsL7Dl4hnYVXGFgzGJbxA+LVt0GpDLp4HP4z3K41b1kd8
R5sQkefzpJ+mo+EGUgiXujl5UWeg3LSHu/cyEL2pcuttEECySGw+iRYr8F+dA2Vw
tjcykmMzRCZaUxcbviFNlN4DuHuU1OuPwyKYCGvIcrl80b5Vwbgsb7SVfkBPzb50
35zCTo89pg1lOvyTAjYFus82OU79pyr36mcU6mxFEBBMwRjv9heNJ9NGZk+eU0pX
Fu3Nu/k+yv02bTlTHCOWGAWuyUTj9xnb3Z3g3qcACF1RE950n8U15gRv3cT4OoaJ
H+63bfSRw6b5nG1d4Kdv6xqgpQsn5/gGD7NLbmTC0l9RJJs5YxfLcXeepZwMRwKY
nqtjE9xWiLvqIc5LHD56PHvh2GUfvs8FgYqwV93SBSPNvOi4eWb3mU/YBSijKcsI
p3GufaRTj9/D7ipOXov74Yvw60QMtHCJDSvdoNoQYydvFAAbidKl7I1XuCoCmq+Z
oGkQ5uEhPKewdDWG+cMVktBg+Tp58k/4KQMWAdecLWVuc8u0JbAshe2ECvfxGZar
VYVDnNJV91Rc3EyPQu57IcYUqIU+gpElLZzhZQQYbiUehnM6VCzDgxxrZZJboGU+
EdsoSwGaIg9oYIbrrKM1S+H1fiHewKE2QwpBsu5k9IyJ2lKW3FCsyxk5Z+DNJ7YC
NhqXmIciwiCY7VFrnKQ7vCCcE2QKMhDy4zSBIGUyaVpbc/NiY8eEzUxP4RaLeZuX
wVEpqTj0Ou5KN159EHKE+SQoaI91sqoLuQ9agBDPW/TktJijRB1ZM0FZzoUnAckI
O6lksJS0d2AkA5ghbIH+I08xm9zT27ikObRlw2xvcnhcL2W4IUR65Dw1LcV9ZFoW
A0JVgXaOXSDv3k9IN34QK+8fnHZx4IoACisZEAIIsub9hL8MCDT/Y33ZWJod/s7H
9qeGI0N6TahiZhmISC4Odb+K8DivlukPpwwxDY6dWh1ri7pLTIj51eVSDyS6U0Uu
kNfBhvZd+Guq6nrIsV9MZsFcs++DiqQBM7vtf7P+OACdK/+kyoamMxwDYMWiE/hh
AfdVAa1t5YLg3v2cG98DHCplWIR5czoVlJ0f5wS7aJixKNPfMs9jxem073Z+jaXx
tiQd4XSNQ3hHTA/DH8ogUkex+TUu8agXG4IlCQFsYKX1HnCM4B3wbg2+aqC/TCpM
emUtxEo/ZSP9GNoFrczlrCOWp+cb66ri8u/6oIG3ykJF6ozp8KnxLy4UlXVt7VqG
pUrLstm/1ZkgnicmhQUMTyQ5RWU8z3RzeWi0IgsRKpy5uhS+Gnfr/q+cTpYzPjG3
ntvsC5pf4LcLwL9Dn0X0OBTathe9dgRdAkuKCUnQL5FDQkxIqmniPwLCmKcDzrR4
yIsfoeAR9Qe1We7wvQPH2SxMqaEiHPWIRXQpg8II9yQ9xcHWsQws61LzLnUXwOW0
vona1FGLUtxvw2NZh0stiWLRGi8gNWSobojoAxP/zuT9U0YUYgqUygSFmuq4YM5J
2erydxXwA0wmZ14Jn17jvkUBw9DwvyH60t90JsA5pVwdrcQ6u1ipUOrVWEgawV/Q
zx2c6/tdRhFl0OfqgRLWqH04RNfWlsa4T32SCLND2defmgXmqiOzeCkG0M3DPdz9
0Dg0Yo1i0BVN8Ok2+GeqthxbkddZ5O7nvbPw8r15huJNVyFO1xop8ZoHDau4QrU0
p1EhwYpFK898ezMtyZaFgd1bFsxOPvITq9Zec9DdCqCELhD40ddy3Jiiw0BTRl7W
S6h3MZ8v6DS8HpgsAQNoERhGVlE0xEeBYRsP7lnloX3Ef/wSKyIkVf2zxkwoWnrB
hnDDRbG9oE6FoYiRYfOYOjQ/r6sz3tkOf/0EZOgi4E1flSVvqUoqPn0Ucn5632Rc
51QYhHGGDg1OuCpTEzLkNCy2/6GnlEy6QqTROVNIwpvqPkFMg5L+EvChbtxdS1ON
VFFh9tf+MdkjRNvYsVWOo1v6y1o+cgrfgKZH8DtRMujeNzW87onDMpf0YP2ccWQ1
7IABnP2rMrpS7A3c37G9ZHCKZV8zVud+AaKqNhVdcUKM9uEO6L6LQ3jcNkZ2D8tH
PvQ1TaFoBg/nS9tWEM64jjym3HblfywhSCFbsWPbzlwJEGU4fCLcq3NcMXGJZlmf
bVqcS6XyAQ2PI3AzYSkK+afi+8BaZZ9MsqQo2OIO/j404yKUk8m1tR0XNKotrDWJ
iS66ipetYUfyw4L191a0mHmRiTEEwqieki6n0M2kJ2w+PvyyF/DOAbGEF45qYSlk
FnrbOFfjUpZEapy6E2r98F5pjHkt69F0Rd0QCu9u1bVTk0/ZI73ASd75PJ6mCkSV
l61JLYTw03ECDBoVw9jhcOPwmC0geQikIWllNB8PtNQBpzofbm84h+sLu4r/WKje
rOqVMn5gQuFKvsX3n082xheWJHiEwzRlf5EwbeUy7XR49m6gK5Qio/6i5+OFGySt
oM9jiPVeE3krqOwuO9UUOJzqCDNIh1gaF/fD7YyJeL0UhGDXHFdodpwPnX5+51V9
uBJx6BNxa2WjlxQgxp8iocrEv781C2ksvL+3kIhdu9xoLbNMHvGSf9tUWmW2qjtL
yaXOEYtCuaDUIv9UJlIYYBvHrqB2bbcKQAgdDayWzvMhoas8B2FMglxYKNLylsux
omDjrOORzMTW1CezkhIFMkzekiqp6jX/7Zs8O4gc9tYWgRm78Oa1C0pUiRmS8RYU
WGOZ2uMlJKxJToQ9GZZXGRrclVauaBnPc94XuV5DrusEKmVtNaphQ+hrep50RJjl
PI9Xrc3VwoJ2P14rIkEAx279yuoB0jeasZgwzLF36OceaT9p2vMR/B4FAFK+sL9r
t0jdkwcDRmX2Oa4qq1521AgUD+1aQXWevNsCVBQe5g4stAS4/DVYRDuHiyB0PQtC
Bdqk6wEpKUhyqvEdfQcWUcNC69SDJJ7yiyuzVgR6Mkejf0P6NYFgWdR/BcHcLXEw
R7ySlflS3glYA8QY87SrGicua1FNTl+BBYQ1w1ElVSQS1fJJrGCQUH2E7AKKNvLE
XUJiUwBtDrK0pwIVmjsJG6eCddgH/sDfg+P5CH9jOlvuqMe+DNaf/jEdi3GbMdXM
ihTKDhSPDBGhCxlXCV0NOs69ruBsMrxi+Wd7WTuHOJVeR+82f6LFb5nFCZAP4hzg
Spyeg4cTUcTf61FnKFskrLARvd3TJ3VHypZjhN7pk42uDVhYukZeVtWm9kr7ona6
ykTUgohCqDsoZQTIXGZyv80JC+CBC9Lpf7j09kDCtU5kJxF41Gh9zAY27T0SxOwh
KmKl8Ji1ZRAO3is/qaICGDkwtDjZjXxN7XYlbFgCmHb+ZsM7cCF5P1d5eo3zxWjY
gi44wsn7f4dt+rhOtTNrtkSvBOgsLAh1JVE0MlprP6VhqW29n7bHjchdW/CZqfYV
X4q8JvUiX/j1W4bpxfjGPWFtZYo4vbZd0JPTbCNiroy2ccIrUNPW5HexMKyn2q1B
EYKsQJzcRpiOPWgugW6724IeK18Ko0+RId9+DXZvlXrICcHy7RD9o0WdOOPJc1Gd
5tiisPgbbqBmLKba2DFe19ngK/hIL2tHDVvU9MoLsSGB0F//qyIxdthHRLkp2h+z
rFHgXlk1lr6mKPYMK3WOlCxxSAag0W2FpM3Ht0VXOn4TUJrlm2puqvZ/Y5dJ+sPR
8N/2FOIkL7EC9JcawuIhTcZU6rRAsYK7mnTMbdAMkgvnDpRBBibaNpjeD3T11t2d
Dpiux+Cq1ZKVoq4tCUA8MYAxbg/rNRbL3rEHk9Bl4pn+JCEn76WC1hAyxOcP8i4l
oeshwQoyRD0CUrIpDrwJD291RCQKp0kgN35dtl3s4JYxcT7kxlgg9zTiiO6IfCM1
tDYn4qv1OWVR/2F3i5UAavu8NphEugylFoMMaEuqeg3GEpZ0QuzeYFXFRxb++T8v
XH9i7YS9EcuDA4azzMSNgoklTSE0nGI2Q2ONdp18y6fUklGe1i6ucG7F7r4InrrF
yML8f9geA9dUWM9zUs/duPw9C+qcpUcgTmZwjLcj8xCEQ86PpfAMCJz1IMYqH828
RTvWL6OMFQ4E7uTPYukcjncX1H1YMRbTrEBmQMN/IrY9kVLuqOAkMIASrYjnGCM8
LBVm07gMDUDnWDDrYWMeMrLkW9l4QYH6b8VhRjj0+uIMmLhqDBC0cBqlI5YICgOK
8W7M+CUcR4PfvOuf3Iy9RbpEF6VVAT3ceyhoCqdAHjs+6vs2a5SSc2L97hKNTlS1
ayChLma4azghCoSJ6aPsuLS7YTES5Q8ibihyLjFubVGgeNUTC7/111JAcfrFteFv
LgGll/yGoZY2/5R+dkQ8sZv6cvnxLP/+yfH99JayGrjun0TxT1ZMiLIkmfHwTubv
OmTBLwm7/scz+x1gOTDb+o/bKJ3L2r3aMB1gjiIK67JilEp2ig4hYWeEeD7jOqMF
cu38X2H6xj/l1er7dohEC+ehQuJhQ8jkY6m03t4GGEFblQwzcCgm5ZupTIH8PmNd
pL/PHSNlCjw2otq0Y43DUXFbKsFBSe2MT3Yd/+l5os8TQUaYW5EHdj41wKAsLZeN
Rn5Qtdt5bpCaLolaiZQjZzy7L2Wk3oumx/T9xSVWNJ1gQMVc4JOA/H5Sj0l4kGZ9
kIjTFZTFIIdf40Wh+2DPT8Zn3wCxkserkiQBmaDb+uFRmpeBXwUfGFIXT1Lw2OH3
twkXr7aYj2SzX3vlMwWEZktlPlqeq76ccwmBOe17xJnKZu/VP8iRIeXZh5XembT2
yOolGf+kB2WjEtAtHZ1GqLqPjYqA8f/Qi/nHJfE2eSF2vugmSxs5WnYtGZpsPLbY
5E5yNizqMOnv7ArOD/YbijKfbRa3puqGwDjooh4o6w/lifkKRkH7IG5BHYHzkbax
tjiuEq473iTZMnXbvPyobxAUnpmOyD5LzWKyg6e3oxi5t2ksGJ0rhtb6daMePmkQ
nUw+ZF8Er+neNX2I7/nJ0gK5laHTNC0qWBZjmBQljcSVZ7WkgwTAJqiNH+BGnuGZ
3+ku9YbiuqxvFr73SiVUNoDOFcpmfvT95bXbdXANuTJOPU3+IQlZQve/NdT5KmVF
J03aMZQuDG6VZc5fS8UYS2vszOTS75wdFNgtUz701ruoRbdcnnqkj2oWOZwR3tHW
pbsDaWlTh8HOjjZqa+9QSd6fvhhnWZraEoBlLSJ7y7FonF8qljI/CGKBZvPwA5Zs
J8BHbTS6zlk7G34iWz0y+cXm3jmv4wqDkHD7nHWzli0hI5P8su97c4y7uMos1EHm
mzlVWcvMhbKk1WO75PctJvyPwptf5k/Ii3b5Ua2AUgxniwKnpv77sPXFzSyRqnXW
8Pkoh2xsTYlnfq+JCsDdP0Z2mBaWxI8meOW4EGf55QgSzjuxWXh+p6cbCcqRauz9
UM1SeBNaWnNgivpe62SQJkWjowxaKuqSWesB8YdB1RaDDb4pZ4jc5FiH4ss0zKy5
+EM8YWmUauxEPsZbHCBVVP9kRY+oXKnVWnkujC5s4wf+UK9KlEJHWxN+NjBqDhlF
dSIuXu0eDrjDqK0T/ewh5F20ZM2zH5Lz9N69D4ge4gsIA7RpktLhimL5lUELW5KP
RYK9NZ9snRoprBlHX/Z4+yeUoecAQbMdO8ct17J7jcqjxG5RTvkRcQq+sGppa6gZ
5tkqL2cr5KX8sPuMWLKw5FWiNXaLJ0XQa/u41DXZR2Ubsw5/nnc4N1haTwOVsbqi
oErmCOAOWBR+Ybf1UgkIXstIsLJRoi/vIFqGsUAF2cNrUz1xC+ByaT1sxYSprPhC
95vilEzVdDwqRu5PtS+95hkjY8ltPKKwdcsGb0BBufNUe1E0P9JdgRWu7f+dW+aM
KPe47QJI1344d64FAqdB94FNbTseEZ+uLK4MOZBSpSQ7Jgnd8bMbqT9RY30Ehk8H
kwOhuYA2gBEYSnPHxJbqFNlCR83o5+mvq2N9lT/Mlbi7kZ+edEutSPSgGDwVlG2J
xitcxqNeWjXLmo4IhsqUZw48DUh2El3Es2AZpkaJYQUmXoW90EprBrbEHv9M8snO
p7BrpBG02MhkX54YIjMyLVolorgvm3TdsbZlxuC6jfhb7BxJBZpbmxEyLmpGOIJi
dBjXrr8jTEFdZ9TQ1j+0kuaDXGwiMlSZP7yFWnWvfTi100rT507Ckt7uakOFNoKj
QdEPEMe+zUWcgxGKfcYvr4v4LfidFbDD4Q8KWZYAv8PuGiuQorVQBpCxUEZx+Pw9
ie4/SEmwsvv1bSIf5yID+aeb0Q4JN9kzDHTSWthyWIxNLwW4C7Mx5qDUxn7uglk+
UROL2yW/OOMZWQjc5lU+tHd63ZISvBSfnKFEopBRMeW233wLjyVzHiNpwqNM/G7a
oFZ4gJOEP74RiSG7mG6S9Yvm7kbOshf5HhW3fx1IoO2qVfEjVMsOaeipRAIW4heH
6eRy0mV2CDjQHoLf+QywaNmYWrXK4F8A1Z6Fr4aqVgRK2JfOoa9j6/GHoBRD9DaT
wVi4j5Kj97ia2zrJajr6wt4pyrRWQfV+B2PuWXsHN6cCHVAP2jK8vR/u35WNU5I1
fofkzR8ymfjXGKXERdkyCKg4aGqA8qn25KcCsn4vwZs4K9ZPO7VszGjDh4g+EPAw
YG80uaWaikCDvXrnXDw9OG08rsuysLO9aVXyfHbpVi7LONz8WfvGPSkPNaxmjjJb
OzNYRdwhhbDfpOLZ84fYyt0Jnz6O4rMlhS5ee0aaDCzkKqKG9pnCovs6nw9ueSsW
WERPGObnfUAdO13Td3R8sOIPV6Luw6hJY1N1M5C4/GLduuFnLYVhQ/mKDT4nGuwR
5iXmbwejDrpoe5Z8Ax0kkLl55vg1vHr5d9tmyXEvaHEh0MpUltZRRKr6J4XQOfDK
oX+noXZCqqbM5omOAW94OQOknbz0RQG3FS14yc0svHbGL3Qs8i0TKUTQb+9JyCYL
X1IizzMhgH2dyKuUYnq23+dJyixSOetI3C1772/Ucca3WEXYYzduOlkyMTAmLjAg
csUfNXWQgqlq9kyw+6IbkwR1C4fhhScGLTRyax+lj1wU5FMI3sjIoE/fAVaS0Lfk
m5Mxs4omEesyyndXppfGdW1X6yP2HVOjX7dhCkDHKRW/GHsstde2m5EnvVAVTfT1
yYjGRP3kx+SABedvqSCQKQbNfV0rsYQHtQ4lzH4VP/tASJbKa9dBFiCaXEGn65Yf
QE8GJum9HGy4J3tyhRa5NeCbuLhfI//ZSp1ce19QVrU/ouSmRPVDJ3Oa5q9CWPt3
4jcV/y9oPKR/BXALJOaEWABaAzyYtmqFYB0MupcGDFuy9hnyDb71htu1lzvM6qZA
Y9OWA8bkV8lf7ojCsUEUV2Uf0AmLAWLx+mRPTtVylN19YHa9SgPn5LrzNGVp+NNP
1bgi3H/XS657mtsGY1A+RjSWnvEB8bXFCm4/fuecYyejNPNdrKpFNbrYcyg6zqGe
olOu4adud3gDicaFUO33NXcmZGhtfTjIlWSiiBiSmINEzTtKuLo9qkej+AMvZ/48
60mFAe3SXxPECPAWuLJM6IfwkgO56RRxuTrtFsGfZk9C0Jg4HQVRgh3rcc3d6uhG
QcJcrFg94gMRVETsXX73uOQQwcrHuuguvDiEYRNH4Kd1ucxjrBXwqwGMHSiW+sXV
tlZf28yvZfBp18V1h2hulVjqc+mMki+Lq0/tWTxk4HALayqvq4Dg6WffnVi1RDwU
k+IXqbLwrqfWbQFw+JdQyJ8/qYhlGEQh/5XS5dNxqNvbaNR/9Y9j8EOjHR8UTf4V
xYdROe8/g3MgIJqADg9yoytETQ+pxbwo5KO1g8ewhG1FVI4H3PgZcOtai9a/CboG
XJKI/HI9UAULh2xftF1VxhiVGYQWVNs66L936CfR5sIDRm0p02Iuuxdm0qPHvBaA
7OCwlbVZ8K8PIStN7zVvZE8CrMTglBN/GJJ0vvczOJfqNZ4quKlKg+bZZcpSAL50
IRGXrYs0QqtRLpqKwX4WQwsurkfVXXhl+h/NOyW5UzQlc/0RnRaQQfh/fyHoXMxb
qdtzdvSeO2nx5EvBhXV7a/C9KeMnNeIKS0INcCdd+kkjc4/zthf5FD8DKv3PXXjH
tHPMe9AJmfohBAb149aXdceYiQmHWCiK1sMdJIvQxAn8csIhQtOiIMOXBmVCgtOu
EOvkoboYWqKXrQgG1eP5crp3QbAhn4OHljnCeTnAeu3ghF72xpko736g5zgVGbSa
cRTjnIZ69aard5H9iZSIpFxQ52MNio6Xx1gEdb0xkw3UI+BXdUjr5hqEWb0GDFKc
rtnBpus2z76vtF3omNlBZb2OI97Tl4nXZD6OQf80UKa9NZuaRz396TR3majB+T/G
lELPr0iXEiEniYq2Srk4tpXXoc+1d957n2cXotOa7Q4xP6peb2vZP00vA91iBP+3
gY+qgOM/aOW+Ug6+Xiq2/RvEqLr5aAaj3UBGgy1inEE3tq2nZFD22hSNUQ1j3Wwy
RvTWMb41P0veic8YS8NKBVnE9f2i3Uqoib49cfBWqXTtVgUmHilXoOgojrgeoT6s
C8BF8h0rWVMWCMvJqZkSziT8UN8RVT93iEhnRN5d2jUrCWtqu2Xbfv9VuIWfkL0O
QrETzmxRsvBjMPitWT+EogeZ07QF6w/OMUOQKjSkXTkCWYUmfPyIOU3oKIIb98uK
6OPLYN9MiIJTGU36XVX/bQvl1LSiqcS+2l9kKvtHeBhEUFqlCWS9rqJ4QInh1Qk1
YFIG1BJMtuZ1JXC2l4jGoIe2aA6esYr5viQf3vTjJwWSjZbVmQMUejPSZXctJiOT
3BUEMrj6LkkRcSKXeLfqzo/3jJoei1rn4O++cfhWuE02LymLBhi7b55EHm2oA8TM
fCVlZZVxnIdlg5WjTUvIpnlUYmj23Th931jWOCWBHZhMj/bt475NFmGFXvw8TPfi
vi7KZrrGboO0bYTadhItP7KpvGFETB9Bf9P62CZlMxcTckO690/TR/Ni4qvf/QId
KysL5JdRle5WiFLavR93n/C6oW3HWECLEItWQ0uo3ZBPAbCVQpNxtf0CqPMGmBqN
J5tKYuuNdgQBGnyFLESRur5od0ido/KvgVE0Z8pkRrIZziI5DzlXNUG5Lbnv4/AR
jcIjZhtMfZ0OV2ahwbF9CpqefWrPDRidj4K5F4LrC1cbfu95eeAILQ9pebg+jqtV
UFCBcYa+WKbdZHldUvqRLQYWw9F5QC9cxF2Vv01BsY5+X04n3onQ75NxCjjvw6yq
Hq+/6w0FR28JT+7CkUicQI9SquD9UIpXqLqYi6Yt8yYca5YEnDDS04RHUQmNqZ/I
wWghw1vycW4CBYj3FboFF/MBNUWZ8Qh4YeNRBl7is5SO7BrbNrshZ0uNm+pY+vdo
M/lOaj74SfhgoXRwjI6QHrGbF8hNJDK4UF2VkLdAlh0aFrioq8qs5IeL5cQBucIW
oOUEWTAuoExMXJNCts8xCAR6+940IZ3UfypaVH/mSdcKqWeyMwibyitikDgD0Wmu
WKndBZdcWLoure6LpzByqyjhMno7iiyXbepeLSrIuz45sFoi8cfM53jupDy9BrPf
w55EGap4bGLDvi/mTYN3q3kYNtReHkBL4+IM6noMQ8nIvVnAp5lNFA5tY/6nraD4
1+tSN3wMlSxhgrESYe6WwZBJiOfHKw4CBk60Gq9vXqDlywIdYkFlXSMvWbcxfo0G
tA8OuGQboT9tz5jfgB9uOWnRoO5UHjRPDVfzJ40W8eGl0YyG6XY4czfvXYs0wcgK
OozBODGFhxfSg5RlNDEGynTocfvM+1iFLoEijISdgP4IU2Qm1O/TJ8ySwG6GqtBc
0piHk4JXKtGvK2XOe/jSBsD9LLrKaKE2zwKdHCkbpjQnyxtfsd3aI6tanpW2o8EI
+TNZIQ/DakEZsCTGkNQ/fuTV2q/ja9GjbSnyzUBg5+JGMY2HV1V30/XskSkUe5Tq
6CAuk8n/PKz88gQxoLyXL9EAIuNnxsahfOedKJuA2uc7LK19++Fv0bk5YqQEnC2y
RFrc1XMecZbzoQ8O5TnLKKMGf0mdN3bwT/0c6BFcV16Iy1ykIogKJASVbWp7wBzy
jP2lc68X9xtbqs+YCMVvVakcXLsSRVvf6Oi83THDc+Gw9yYn8QWz/RdvLweupvo3
S9MlKCl3zM+vRKsFyN4GS7ZCoWbia8N0FNHm8Rvb9W7vFM4yIQQjv4KM7j9pZcOl
YFO8NJI2yx0yyxRWombUa09D0m+wgN8rDaiqqz/pojZa///9waH9mHKMJnHcq2/W
sO7QqklrT8MqrdPYJUwb7BlkFTRiavAT7bdwzHWYJEnRXJpJPOTvhUte07JSO7Wo
Z5sSkFEo54Bpje+BrVUblargbzhr7TU7yF+vmh9ZN2yaeZdwMOMUL8T8HIPdwgdP
ikMQACwhhsXVPsPygu+amOxxW5ofGbDk0qRvmuT8fpE9oqBk3yv5n2rrwJeoqSVZ
S9HslD6tPqsI62NU75nuuzK85omJq+BuGiaP941n2dZq4mcd98HXlw2BBlBiP+e1
m9kt7GH5z4P7FRB6+rp1XDqXCpvWAE2RAKiUZq6vUBAnudw8RpMl7VyARMyK07+J
EDAZvTP7stBfDXqeO3oBRTEA0PwpKo1kJHa/1m/s7EElcUkSar0l+hZEg/AxcqjB
BylC9d/KOPDJ6rQWqvDxLLwpiUYeMjs8XEs3R83Li1AnXVM8WUPXEx5h/Ml3WgUD
JAOIw6AR4nFanA9v6TAmXF0vhX5wzgsEgnSv1jc4CqAbA9JBRWOTtO6AdxawAU4k
sX9PbeaIHSAaDVTVvIxeEpCDN82NuxPL7gZcmje4LUoA7Tvyk4GKnfB1P5yZ9Owj
VJUhoPW/GH1oiuHfcQ6EiC6ATDKUe7AiZvW9/dwTyQ1uWFjjH/a6ZYTkZL4dPG4Q
boWR6/exWiszVO1bFTq2m6+vtIHxEnW+9N8XQc9E2Q5HCsKw/dp95BBkBqesPnwz
5CcUyxr9FOE9ipSS1KnBElfUy50Am3Gn5tiM3qgV0jG8Ede5d+OEmBn2ZtL4tQ7x
aLz08/CshVL/ZLY5hAxjvq96k/7KlYnqLc6zC/Ej/5mte290+KAOiwt5pj/i7iff
7w7jwB6s/chWk9hoeN8wVTO1GkXzXkPmd6hKnylep/Lf7jqdJEuQDVv6/qSF037f
tY8qQSJ2/j8q3ZLDoGp9ZxPcb8mCaTZzro5pqmaZLpQ/KQuc+FPd8km178LqME1p
Mc+ILXIrP9Yp72qjv034+2CRH1dLn89UJ47IeVKB/aZo8KqdOehHAgBujqA1HF/S
Kfgl51uOHYTomRaQxIZHLr8xbjeMW6i+sJxaA6ngIrC5h1Mlz/03xGTR7J3JO2jz
1oQUW45Am41UCZ+xETQEvK4dRWk4AMg09igD7TKW7JtKQhzdnt9sJP7rIXeYOTlQ
22ZcKnMvL3iOTkF5y2vtmuGwo5D1xZ0hUAMYcdkuueGDgv8BqEPzzlxjjgF97o9t
xobk7NJy04UFdbgxzhBfutqQY5x3oYTHxD//NmcwJY+QvPdFyNkgoI5sT1pRa8Ku
BnOn2O8tM0bJJxoW317yAEWc0Iau4qungQb2/iFcICGPj8vfl20Ql10kHdQlpt7m
k8hbuJIoA760kSMkHZGY8PM6NuLNa8GwJRO/qLHnNAGHTAAx495evcd1GNegxsGH
8+UGWMd9AGljeGCtI7tHA8BINp39FOeC5+7c/ySW0EiWvrCEkzKs459mjj33Fmzj
ECqdCaviffeLO2YSBJWZ8rYOmH7AQl4Ry9NwpPni9Qgb8763axrECX0YJA1mzsa9
yInqRPNpk20ySAOg7wbLF3odvIEfeONnKYTKQ53seiLmvO0MCqRZidwCe4EMR5/d
HVyYfcDqsen/5q++0suyqFb8TDpp9PI2Md44OQdoKqLjaur3QuNP7Wh4jUI+u9XY
CKe2dUxDmS2cdSDNWPfxpBMRL7oG7Nc+9aMVAFFt0g63ae4gzlUxV8z7hVH93aCw
a9eW75bkNgyFpsjc5ElPwHTo/xgbBWdU/w0UmBeSyOKOIbmtfhiLgX4eJMqWu8ON
tVgZC9FJG+wU146OY2uZBjHERRMAWWInp76J2b+V68+d3w+nZz4uP4zSDjNqCYNm
KmecWbGo8ieES3eoyeYEeMChhMnHLmpr/E1tCiy2Jhh3NblKQYDbxG9wql7aI12M
TD67kKRYby1kb2E3qZaWTy2jq5yaLatfEJRofLG15rWPMFsv+DJKFsyuaUje1rnP
KljF0PoC8vywAMDCcV2IqAlWxZ4dSRlwG2g6x3JIgErYN2WcZfzkWLnGqdrP943P
SrELJ+CX3Y5PONej8oFT2+VjmBj6juC7gqrXeze01591043PJb8Q581GmUwrkM06
HbB5ilI+fRSLmYsdrrIUYvLwuaK8hDwk9Ar8yQ30e12ajnUzoHBkFJp9F1agEodb
5NaOZiSiIkIsd17xUQcsI9VbChPv3uFD2zcPlpSTnlf8ceIVGIG1u1hZrLmC1FGZ
kx/O3j3h7Px4bbR3xfDbzgQmPzwt0/Vz5JlDMoYhhldxg9F63T+hpyR6N+GGgvV2
BdeCMu26reHAwFMWkoP2uF6fAhgqKXSvPqSnes7U+DXOzlfXBjM07l5IxzAQX/is
hx8PPEBn6ji3dKHpX78mN2OZAaGH3MHuIecd5DnFbenSUBSocmh0eGkg7CZccBsF
uOhgPA7rcoO9y6AKSAZKQHhLRH1R8aBV+6BkLpn3mGGz9fpn4taxZijVXD9QBA9b
1kZ87joqXoQ94aZfvKxLtCNuAOefwwwo/CJXm+w28RuaJUQ6d9cbOlJ7pnJ+iWe9
qzivvEOTJz1YnKYLkH9qaaqVhQeEen78gLS3JxY+j9+VfgRKz6uy3RmNwtqEyWQD
6LFHaFwS4CmOgNq6m5n90D6oL/JKHuyiGrwXHLYr9ljRIL/Gfc77y5Pnk9mrc3Lq
d43ozBpWFCHeVRz8JLdpH5G806vjveID5/FdawwWqb3BEt/+rgnzSxCAOQTX2+lr
EiFLmM3mIZc40LZ9Qq5xN5ryxfdr1IWsgh2TpDo/S5L0jMXxLszOsLdK8UQ1Z5jt
+1gVViBdmMv5WoZvKa1mr+sOYSdcG/hrTMXHOmiV3WaivZl+qiLGZyzJldMCaWcu
c4ipVlFNcyJDQZhdC5aaBDBcvPnWZ7i+xKvN2KgWwg6rXtlDgvAaDOtir1ebYlA9
ypFkVeXICb0Kls9dqWghy5lTbkFc6y4pNLIgpOXRu23c58jPEf9tGcJijNe3XVlT
RIjMU5NWFZY+K42cy+iRF10X31l9C2vETUwZC78vfQ4C1Mq9W1zbrAPXVGwRZHaw
FFCS8C348pkLFMss3zCYd+qPPVRlRwL2hoq9Eg7ZiK8NysrfTdM6fzUtCqmVU0Q1
nyW12SRAiRJnLILWyZrx6zSmVJm3c3VINnkGgKi11LqFC8HKafidDKQbbxBWhVRu
lBb0Jsi8AcR+wGL+wKJ3qhHq2N+xgEntPyFYZrHn6SzAoZVRTDsu+eS1v+yA/IVf
EwF7wTafYfUTns5/nzeKjRqF7hx92ZliR5ewEt5h7RDoLb1fet/V5gVkN/ydwLnu
HLahcW/jAYtTFOKRNFf4pgevexbvamPFKzvP4n8MLv+Ksh0xm+Fyv7ADPNw7BRJp
NT9dh/mTy3B3pQzhekorjecKMb2DbbA2S8SdqiPGu/BjGJjO039Z728UX+MgD2iG
55z5cMtV+HM8OoVAt3G897R/uUKEjWN++E1/ysfdo/2qIQiNKdHquLG6CGHaypMz
lHzIG0EqCuDjWuKWeW+G/TqtX6Y9uCznDZSCTrFs7Nd67Ue3xVChJbrPvoXZUZF0
nebuPXJx7Ca8VEvZ5WVUdWZ8CZfteMxyI3D3Pq2vmh9YKY2cIZ49kaMce0d4xyMo
iRmeznjJO7UGfczQF7lUwU8rTDG9l/ZQXfsvqQHNqwz76wpK3USRZHPFl67YunBS
P3EO57GndL8GkhBwaKO56QlNxT0ymxV656DOrSt8MUCJxWiludv0TcsbskcgPxwJ
3FM7P8VMvbHDyE8Elh0JXtbrY64Bzc3xHyab2lmrkCKA1L7pffBuZIVyHzTCx0qZ
2Z0PiM3wCYNZblVukGkhuZsOZgn50HzZ5xSdxcwq7RBEXZrS4OOJyqVkFwCBRTPZ
nvDSM1c1tWE6aRCy4AEtFFtOdx2Cw3hJlgv8dpDMq5VafvxGbZXtLscju+eOYaGx
n4AS+Xz0NZRirwws4Hv952TLs4MYF6S+Ngu14H+iB9+FrwzKKGZcRdxt3dMXIN6d
7zej5tszkh/0Ou6Zr6/F1FVnVix0Jst8VFIk0a002l2HLXev63HhzJk8Dsp2ch5f
IGMRV6Oaag8gXPZBlEU6kSmLSYEL7Z/IoRuXSrHcUzdE2HaLLJlIHPaMXTA1qyMR
fXWFR39F7gxu1Z4jj553YPGLaw62r4ej9bb/DCOmKkdngC7f9gMUsK94eD7GuIh7
p2DVcMJcTOCRcahJxg8edxNReq8R8pp3zKSJuvwr/WlbxATmKft/FKBPSuG1BfZs
FfLCCEpeG22xTn93s2VXzidoxkhOhT0Qg8xKgA46yIljw8chXNgap2ZwgIj614rX
AbTrnrLYmKFl7cfuySHfk5yPR4fpFRizdFXiX7n69f60GQkqd9IpkfPFJCtb+Wgj
ofTmhCQiHOmmlM6uOKhpq01+KoAMBplmGOw+PaDKBq3aUwrQTOChndx8SAFF5xI3
SE6XuabOEj8RIyiupujzG0YsHrQaBkRESqcZk2+WUh1f6XDjP19f6yavPXlwQgWF
rd41cJbFqWfcv7EmiY75dN3Egs7q/aUAVOEB/vtrq82FbyqKP4exORUi5ad11n3f
+CeaYsYhlRj2B1B121rEtWdoajtXCWTYQi3Hsd7YiKZTco3Mhq+jMixuEIpwyF4k
2xQP2PsF5AMpl/sF1ZxYXnuCQFkG1SFNtYOBQc5Lz2LSjZu23fyu1z9n8UHVSVIZ
KnAEcai3OhamQMvdNBqzxgC2tQq1fCyQNvbStA4LDjjLFmofgLzOf3wPwy0tzfH5
0YfxDiKTkZ9dWCFPBIvhnG2tDhvRLOSQwmOe7mNd1jnkBIv3aqKCxx4rjvbjBLsF
wtb6lu16V+9AtQ1fcg/+JS/0cDo7uywx98acQoi4jR3p32t4mWHddboI2fpPJYya
th4Ve9Ui3MLGE/1xt0nd0+oc4nR/F8klFERBtQmzeXBqqC6/ELlKIwzumOxQb4mn
ugyjS7sJLy2mAe7zednbLVqwq0BTyIdH2MrWukC3hshAyvr0RavDzxzqKd0rF6KL
Vw60V6aW4hbG4r3ZrgHloB/g4JTjFFjA3DaCYHG/JAZ9SQuretI6FMkbBTCo2AZa
ZJbaXWuHpintLBhhbc6HWTAiUlxy3HgXuHgvCL3GpnYUzIEm8p60KtXQjdsqLn3U
/2fIKgZ+GGNsoSVHkDduIxOSXuryLHbQbO+gXdTew/PaKjCZ7vTboNKXVr8Pz7Hp
6BOjLPYbPNbkpfm9XKXbQj4Few037HWP2ulzeChglRm3ZTARhzQZA3WdD4c6G46m
NFSg7TSrdvzL09yuc5weIdXlpySjQ0rksmaP29RTNBqQhDGScUGdOsiMLVg0GAMV
UuBu6bhk6QDOm1yRyhM1njOZHD4PpnDU26XlxpdBIP9ND8oMfDCTTAe+yDO9D2c7
RvFa9E8hVo4HXiLbFVUKcXRq2b7NMu/nBTAJsdmVRCOL7rUM6VeHjmx6G31v/bUK
+21S12ZjJ5jct7Iy2ysQa0Yl0zY2yk0MOzi8DHHfWvFuClxEKGuwZQAHN14i7FhJ
OEn7oMDMyY6h3ap9qAx4cdbYgFGzEYEI9a4TObRX3AQo4r8Xutxrx6CTrzxV7UVT
Y16k5imm2KKtvCRuDjQV7v4/UHzldL5cd8FAAuqSGuQ1fz7yHSycKiYEC5Imhj1O
OTxCUZt4AEntJrxs7SJPo3/wb8dCJM/YB117hdhu6AIjVVXsldSPyRQBWsPdBPG+
1CWl78LkUSD5fawI1SWH0PecG4e70j1NMYqLzLU7pVW5SAAWM6z/nIWl63IY7xyE
BwYrXhuKt2hGibPTB0WePU4VjVeFK1bjj8S+1h8IECmeHaXwBO3ZR1S7/QrFGGIx
ksQP1Dxgntpyvd8Y5eywePgMy18J+kbmJtnfZHMCKqTrWJeKf75yUZi4qgcJ9NEd
vUSTM99CmVlVbfeQHwF2n2EGIdewOCgyr19LKmWxNqaA+WWjPfUsacdngXX53II0
1STOf3QCv28oMFlVpLC/tcWbXC2KSiN2ncCNrEJ/O8ZDplxGAX82zsL7zUU4sJRz
UfwyjxyAChvenc/F/AHnCdFJA751u2co9qEdFGjPkVMV6TSpSt4nfuyEgDCAIazj
0FvV5Aj9WgIWmGz6mM33PomKv8oUZP2cy61ZF3BOviMT+UNDWslgWxzBwEVsLN78
pqJtiShWdu/aEl8kRMlreUSeZI3giMeJMp+4daN+RHSSopOCByoY3/zsShdK0614
M4jSQd9unefZxCOH44bvHiG8QG8x9OHimTmjj0kzcPCc/f6pImZiNLm1nmNo+WJh
PDm4WSWKd/nmqfEdMfVNKZ99Uy2jCowQufjJ1DERKPvsq20fBVRFIU62gIbMf8L6
CQmChbXvfNemUazgn1oCQlzSxrsmUbEDypZWCaW0Zz818ceQm7PdMS8iSZ3NYzEC
fNYHHGFzGaWXRMWNlnT8pCCD3DDSdvPk/xODqJeyTUQjNA+OLGY6A5RhoEZLE/lZ
YKnkcI0kqYPyBJzf0GUS8ZPAkvy9pAbT95IHApwPhfT5mLweNZTWtwaC3rlz/oeQ
wF7thdA4fkBlHeTtr5p6F0OFC2wOrYAnZ4bpY+Nh510IUMIpZAjpoRbNXdm0+gC4
8Kjli3U92gbPRgXKmJt0ol5I4VOAE+KenetkJu+2BqwhoCGmrenRI7L3GM82e1n4
NOyKH8ZcUqxZYG1klEzoNBQPsDIe7mVlUZAbdgNtyIi4p6c3GDHxTvma3ivdFSUx
ss0S7qym0BCwkpcfbn6tG92EUaZYOrrxKL9zZnK1xclq91aph78pzKHfCvrsamf4
fK5gDCMEFewHSsAVopsLBxl9lf3czmI3jSKlUkQMzH1sQIq5C72mmlU8RYSwyoKD
Z7JERdLnJCfUtqYrBS5/++bYv2TQLaCUmBdq2tlSamTockuk6Hy1nyHtsb8qxlNE
+sxiwb93qVVF+YErf0HLB2bps1fXKipTvd+bTwBK7osKSjImS1O1SQXhV7ndwuGN
wi9jwgvOkpljxUtKi9YK8nxEJak0H29kn+/DFvzBt40Sc96x2MkFZCetuyGXfOqZ
yfftx986CyXsx8E/00DOaDlbCcT+5iK7GpocpGDUgip7igFOhYEL1sVG+zqVPxu3
WB5MHcueRDUYDgQ3yBtVjtIn7kBX8ybeAoKj/KsGbaVj+bhysYWnQpub4X/j3/Ly
XvgWUktnIdNnMCFbaGe+Fhz31arzTspvRtMTJGa9nmtLgQp5DZV8YqKodPLTQrzZ
xntGGR8LNMzPcj7BoGMNbU2IhKUD39POVE1qZFh3YqgJgUFIv2Mt8BNwGBbd8Geo
baYdSImOp9NwCdtJ6RfXf0GTapji12D3P5JvNr55LPhMqvjxMVpljEM7760lw7Is
zB16U8UokQeBUABxCvys/3h0nRxmcE/1qzl/QWkkUXFbMWhIAT5Gco8rK8tGUlib
DBCC8Ki9KU0PN1di7PQBiL9hILwhbDjzCOrJjNFJ53dfynRuaailG7Ej4m5zkKTY
RyTcBDPVhgmJqAc88BYaEk0j9t8P1Umt8q38fMYiSITMVZ7RPYhFe68JSACJJszT
062/a+7e/5jisoeRiUYbctZgtZGwe/f3+A63FGU7tutm5KVye6x/4sEJ9Cef3mMR
Y8UuBwStwXeKHlXO/yyuIuPaYMfMlRSKdZkU4EeaPfaGonZPC3SxyckAZq/NyIuk
fs+9pmVKEb0b2l3g38D3GfisR9mP4LIl17uAibqaZ83Ijhm+bOp0ei04f0jWV4P4
qUNWJtqS++TQaxr8KcHMF5g96r7blc6Jdq93m9Iq0LGtvNF1qxLY11Ho2iRLm07K
RrF7iQLe4JEEiNXrAhksvKPY9A6hDpTD+hRImXGSFEQHkC8tz8aG+vfeGJeR21wN
EsTpAGvSk5T/VuO7wWhWAtvE5QodtP2Rn4SVU+zyJNhVSlONZhJqDl+sx2lqXBR7
Sz7y/g/N54LVdhNcAw/pfTePI5q7OLjqlfzMLksjMDI/2QTjaAwqijmJt5PqgiUT
mkJuZKRPHFfgpXg5CofdDNT+hbKr0dwBn46jaGsN5IIEhpqGftNi1VuHGcuWS9Gd
mTXZcTm9vZbPjIKNKIj4YoSIK+0Q5wzXLsdyyV8nZGDI9qMG/Qa+0OkrYSK4zHv9
GIht0HFtDB6kxOM9q1hSppWl7CAhrCZZgDSA9FFF8Li/cIEhh/bgypEboLE4CiDv
tnMay1m75YCoyvdAwRHKFLIH9gBYA0LY77Fsa3Gt3brp+4EhStzC4nCTsndlCz+k
VvjC8woGi5Ha3djuLzHLbvrqaEK3qVye9tjQJlrrqqHKDgQiQlSQ1FaPq7ldZOwy
titSZbC/agBeqsZ6v8LnHWD5sm7Mh0CYmyKg5GjeRYmp7u1afSppvPYKRmuEnDaZ
o5Qzk13cC9m0sq98niimLcyJll+piQNk/fJfmDbN03RnIdHBh48PAj6iPb3x+NTj
FTDML7Y10gZywqwaFWB8vHHDVQDdi9h5ZsOseKZBqwNERVxXUOA4GQhtos9bt0Nh
yjVZsrFWM4xyM53cscZN8e+FEKld+gp7MB0NMcxZsFy0Z7NZHQk7I4AM6nKEh1+5
kFe45+PZePfltBTxlkL8HnrgiujjVx1hlDiwj4O807wfvYInvGMvA3SHOQ0T6Jtk
1EFEHzxgc0Wbukds5ItMjiOb6d7J4po2UsFRLEv8+MOTkCQtXbjB0G9H51i76rae
SWTQO4DHItzB9wy65zQeiB+oB7+E8APX8LCyuu5giRd4cHVdfPBOq90/YOk5HtFX
GVuYJ3ra2PQ9J4LLdgUuD8QSVIqR4ESV0XBeS8rn3IEhhkHrFGsNn9T6fK7QpJ4J
uQaPwBJv6LBqaKjZdQLhrMD5ymtKW2w7+F9yHfRpcw3kJAfIbL7P3YPZiq2KIwGa
+iqu2IQ/KLnQXWCN05Jt6UkJgg3qFWNx/Ga0DuNd/hAyZKE9s2jniSoyKY5i7z3w
iaTFDsOyXR450c/epBh+dr7vOtDo2MDaCKmGTf0A9kemrEERz06dr9fNPaLFF27X
BkYAnqGecqVVZUmBV+FXOkPN0KXsi7qUaziucVL4B14puuuSAo6aqyKqXgAxZCPY
eE5V/pXiOclNVPAM1+KVXV/EMKeIIK9TGsyi4hQQv/4RUZfPLrZTvx+mOf89/gvt
toRqPLvj66czvSqkTsQRUs7rUlz6XcnJvlefQ8JCQ2oIOuwv6Sc7xQ8uXZZOZ1xx
nKbFrDjtmu83UEILrNEtdihtEOwETtk8Pr6O7cB+fJ+WjK3mdWJYcWKv/UwSnJ+V
34wf+qKbw0S+me8m2YrwqnhHohUp9ON/tEn464PfZmbyVcPIbBo/8YqLybgoa6Ue
yvS1mZS7Hs8DD+6C4HiptTKwsVoNtv0/dvDvnrzFH1HpKDSYttPrI1TIYYCKjRhK
0TMdrk85F0ieqomICd2qA5o3q2FfLSaM+9cuWMTUtm5tdbVJbkB6Y5Khg31BKxIk
YDcLx16jaWlKxHqTET4weJTAvOLASv09UEgA+xb7rqVQTBo3ZfidyCnkfAP7aNlf
bnpMtLN1qdwKr3zCrEBYVvCRK3s2DGhrthKmdS6iGt6lFvdFAl15Cof4c0lDEh2I
Sd/NIJ6eeW2PFnJElkVU/ZMLjZ7ric9sn6M8IkY7nCIn6AizCkoeDCbZypt6Ha5U
IfJddrF7uQsXLFTwOfaNXq00zWMNpub+EGRkVSiYIifOzxpNX/0M2zzXi0pKKrcN
sd9u03BEnLyO2oMTXwyRfM8yBK5jTJR3oTzuVp3nkdSK0GOK5O9GbYTHoZalwU4U
C2E6o/fFpF48wfZm/4zDiG2SLtzb+IL90hVrGpjkCGYo26aXNjINfZD/RxksHkrn
ZGn7fYuGKP5wUnLunWYZXfL/u7m4p2U7GrwfOE8kRO1pkJSZb930ZzT3HjBwBt3p
A36gIP3D6ZskX2glj9zKx0TTcnUvDwMyWhyCnzql+7fzPc3o5Ui8sTd34+fpKFY2
mr1Z9pMSJ12/0+sAJKLVEmbn3aeaCnN0lfq4J7Bivsn2x4CP+kzu/XrE2rD6SA9y
l9peXTpcb0FmH7lQ6U0SAGBlbp3m3Jq5AkmCh6qgnurfm3y5Q4DXq8MB/Kzut12w
0yx5LH5khgaS/pSnUeNcVpkTxj+0QeQYQauHeeeyQX/Q1u+g+plxZYTc03cmlqE6
lR+RKLeNvrj1lMnLPW19zcQ84BAfci5GIpj0E+sr6KHEdEpTzEn6tNNOc2DynzDx
eWx61SweIK4CNbKmSN94hrttdwo5KfCka7WO0sDZcY3ASSiZ5dmx+nfXBaRGnKLk
xGdUIme7lUidqWHhF+k4RoTac+8l7p0nSAtmGrwgmlkgjwXvxLU1s3gTtZN53Xfa
sF3frCEH3Mi7kjkc6oZJevlaJxUX+ZTto9mpwjpyeUtuNjTwKwp7nqkSG6m20BmB
YeUX2Hcl6BDc2CvS0LOAmeTJbZanBZtV+SF6IoqRGQmyZHjfJCHiwlct0WeZvujj
xuzMvN6aIPKm1lLvNGPtd2I1vO+NWCVgsirxexErB535uVWynmnXzTtLz8QyTB+j
/2gOBVJhzNFKlSJ+Ys8eDIgVj4M5jyslQ4tABBFgLPK+d0Pva+nQIoX6hUfuyjKA
UKynCO99PXl+TUoQyVG/mJ/xcQ7PMQJPItnwCVBxUdatwsakkORDP0vjCjL5k/nM
Qr+lworHpui2KxQCbd/W6yfiYt0SNugxWG2dJVq3OSIrabO8vRd7izNSJw7P4pt9
LkvdVBrpCjcipEn68GoWMOgFrp9DelQIRSe6n7RvtR2GsA9O+diWSGWVY+Qo18XB
MwJP1Y+8B8xRce3otDfX5jj/2vkjwMXMR9K8w0LUMI0bzf6LL92Jk8ZRSC8MQcDR
a7KE2Ks58hsa4XsFA8eXPQr9x6xET7JF3isKLgAG0emNGs2v1gihFCGupMvs34yq
tLvbhjT4HLjZJ/vOsEpWgM4JyD9QDKREagSkbwnJOFYCplBgP1/YEJ2TgrkE5bjn
DUzUD2YOtviKZgdAY+xl39ZCMlzghFOOpcRzHXXx2jBidlzV+MbdRIegcjRbQt1l
FItlwz/t361IjN68dgCi7hl6LCMZHSVcOS9gdJzw0WbPNnk5OKZpui96YLli3OMn
qNCvvoVoDsHggJHaAFIw1iZFqSWI2RuIoAhlBP6fwIqF2Q9nw65gmf8ceUtPCvtp
YqeUzhMmMlyVwXcxebd4cg0IueUc/faujRHwWB5HQWr0Vr0r+agiLkOcnXBU8VzD
eQUDX5NbRFoe7EzNOX0yddAFM4TIa8+JBAlF7OapPEJfyzKnPjLEIUKnWNTbUltr
RjohuFmRDghYE2yw3mvHppaomxoraF2G/VqqeeASIwSH6bC4wL9w8Itrlxmfp1tL
o9qA9LC1v8E0EvtsnOxfHeOgzivuilYWB6BeQ9CxT2Bt7F4nxO56G+7MfnrA85gT
EdKbJHjbF3wUABBBlrFujTSVhvCEzpxBR2O4nXn9I/4WpW4GzlwSpVQMl2yDGObc
0dFgPNVFdos2SEzt/CMojvmwcn8/8f8HPQQMiIcYuOGlhpmgduXTPN/Uy+qxuqWM
iY6uYBXkAWeR2Fj0C164dpenhi88IVb8K/MzFQOdiyrDMUl6RlVH6bt13CoFbrwy
Wphn0Qy5RrfbytFqemBVhQBQTiRhJ4fy39DZB4w5HO+b75t4mlz7FZxB1JIaLmq8
TP0X5zCar3Em1RLoWtreqLNKFTouI5Yho/3F7K7J0Umx2XO9Ii05W3Uh/Qrkpsbc
3PdTHbB3DMQithSD1bdL3rW1XOVNqO7iem8S+RF+Q7vIUe+IjXZBa0JGmwJC7ulz
iWTkUJPjijXI47kQTs7LJ8eWLKp/iyvlWVditx60jlLB4YNrqrtjJhcM/efOtU7V
MX+9Gqt6m2EBszEHhPRsBcsHgjDEY37NK1/rrIBHrmYmih51Ye346ljiOWVwiL3H
3OOzR/DtWk+RFb2eFOEm60eyM5rrGQ4mRi3bK/X7Mg1wNV6Q68kFLl+YzdMQAW12
hnF5lIxZuTu/hRJy7BGC7tyqoHjm2PXwpKs2fhRqxcaacCZgHqIR20Q+2AREeoGb
saeDEW/6eQ6O4AbesaRw0YSXaYnyhT9VrEHB2HWr8TtTJ8ITxNNnxzKcPiY5uh9J
/XkYI+4Lmbm7nv7q9pqxQ8SQV2444P6cdfZQtok/T5FQ4KHhA3YXZDvoZCOqpJ6R
YrgexoqeOlmpNNTNSUAPW7/tvRIytPA1ZXaXFHxM81jeZeFr6lYRNMLbek+q2sSm
WTqdwYXBo8C/lpvRyCn9yCLaVSOTConpfZdEe3EPSV7fFU1RcNkJMgN51DiDOhW4
lb5CrDawAm0dC8NNnnPVXj/TE1vdEN7N2AoomzwKDoBQzmjn0LgxPqQapuIfz8b+
LYmzi+yPnhuYBveod0f3cCGInAwrpNFiNvH4ec1RBQsdN4iJoCQdF738VDhLMz+B
JvCYnY4riJYjmjoO/xyqXPHyQ1x9BJJKnp4CaF9q5lX38kmYuFPQykm9Wkut3AhB
jLk4W6gAcPDffCUHOa60PPqvy3rbYC7ll8+mCm7KwR6HK2hetAqjQrWOvj5QZu5s
3jYiudOOG/+s5s6nFB+FL1b4ffzbhQcpRVca3nESjQEOYVZZ/FOpaTqaG7cVDcHy
fAFavG4udm5RrvgGdgUS+cPjSkwOq0Vnpp+7TUZ87J3xPRnwN6rHV6NlOwgIk4DR
uC3H4BtBPgqNbe/FbbYR09W/GC3bZh+4ZEVNhPyND76UkLcsQA1y+eUjJkJOwfvG
Y49txTfPKyrvpo9Z7O7hwiXSPDHPwLyTb1uBzw7pH9acx6+WkyQFareK6KiWAtF6
hr0pbHH6Mfgk95ev/dUAVPfB/gdsdYGdJOC9yo5rkdMLj4VXMdTfS5C1KT9EvTxp
lzWpKyLsR6iHS0s51UqbrRmugukFCbwFXEeaziU0+BPiRqjbX5O7l3yXm54ZB2WL
RtS81MXoqRCh1XBI/TUahUAKY395oV33qbfnvyB7aW2wUp90JIO8vw5hMr4Wqvbs
y8hYXEptGhI/tkPQsaJDYvsywlF2O6IigFQhbLBES/EnKyo3ukb9aMprUiWIuqvJ
Dfjeo7Dq33Ga9TIJpuuJA6qRK4X4d8wQAQPnMfGom0Pzd0zcBBasJAzCMGczjUsh
Ak1WcofQ5T1bZclVHEUB9YD3sj5OkqknhTVDo44WRZbyDmI4O2B/iH0DWnCPglTU
RIYY5+GbFUXJCZl02Qc0RlfA/+m4/vWmqZb9NFemsmq2SlmGmZmLqJiVsEj6iESd
dT5sudwN9yVOr1/aRpURjAMngKNl3Ejz2aWqbXevbPLyFielh+Immdv2WSXXJkGP
pqK4hTu1B5+fZT0bVlgs5A8q+3DHK3N21zPqQkffAg/Txax2HOpZ81LsSpvnyg1I
e9oddwXFD1jonfyO6c5CDGNq5+xsHFTUo9cBdxe+82BJWT75hjDbiA1haJMfHJpV
y6SkypRJdWY3xVFbQiizLKdQ/hERo+0ZOWPntwNds+OYUbrBQwO5KNU0qlbfMIXn
xXKLaLKS9BtHXquuix9RXTab8uydJinE6Yw3YFmvwhDQ/wfJNSwePlaRiGeT873c
g2cCMo33Jm2OYZ478iilz8z/mn89o7rL0YZu761k+C+S5rwHCO9ZNyT+7fc18h8u
baHDtQElaW6Vos6oj1b3+e4MkpgMD+BqvYItie8k+yE2SWniaOftqezoo5RWhWFz
aEUXsDT2Bg5pGvUT2QI3ssz4zTRMAfxkupakqWLE0pTJlTyEDkV3acdojAthPNYR
nMg0tHlo1qL6mK21bVNTmd5HmJWJyKDG8fNsp6/LiMfjBVlalc0UEA/9uvRtJz/q
UzkRvDWhEdlkew8BgAlr38e1TBpDlvHM+FnWTeuvGb9orpOKozzoQy+5zH8RS/2e
SCb69rtNn33d50UYpPw9tasJ3OC/5TpSkLYZ5P16W+5/j8HMaZUcpku3OYGkLNyZ
61/qmjefmqJAd/vwZYPX7r0qJgFTxjxaDg4tBgYZf6pmo59jPEUr791MqlXTmzyM
HQF2AgctGykA5M0TPStmBMzYFM4thyKCXniRdlZ0FT6p0ZBH7KG+EWqyCmxcH8kr
woMdL+P4N8iaVLPKiUL2isGSxjYKbr3MZcOOjmgxzHoHWTeWNffnPLlsI3fGhJph
IQYfc0FpWgUikwamo4WtO31gXsUgPF1LYwLlG0yTSWnLD88VfpcXpSj21hgLgmB0
wgRmgDBgGk86l0iMEQ14NvhpDvMnWDb47lQjAkD+blfvlUxKezV2jrpYEbPgbtY+
cse73faAcFotZmf6grqiMfLAaYZRZpJiiqPrkTU8v8QDj/hCtxiUHeXgPDRkeGVd
lZl1ayyrn2RibT+13ShFtUfkV339akC1atPW7u3mv8jNJZejEclmmJLuhy8D/6zT
3/nVhD21BuIB1QPgIqaPbPsNTTx4/9wmUGzMYHFWnV/igMMT0rhjMET6Cu+OZ0IE
0486rosY1n6708kmuFWVCp4P8q/59EhMmS26IwosIsIQOyqIfYLX8ixVLD2+28/h
H/KNHJJE8lQkWF7B1lExIrQIB4ocVNUrRwC+rnAFcXBvmNsvYamuABaHnZCKcO7p
coapqYWi6F93GnmFfJNBLEqWIgXCXuPHPqU22ZbcpUhzietLYG9UPUCu5Q8mqpYg
fBiEmeBswi06yxhMAslZo8J+2p8HJaCpCQPG0RSmV7UzbYdiyUouSUhCCV8QPpX9
NpLdj0z6+W5QV8+GBKLljSkAz1eP5XiD8YBDCQxXyWUYWNMNqcgZycMx9UtGHXDP
liMG97dgC6fmUPmCvO3s39Pa3aeElcSZiFR3KRcSjslIoGey1VtUmMpV+szq6D0C
r0RCei/83ySv0DRFL6guxBd5U1//GOZL4L0n6DlriPwSouve9zn9auYDCBb/zoJF
wnEaZ7sC0n36jl5KhnpuKUQaaMhYf31OX+8WvCyh7LjBbOAfFvHdGg7F54gTVZYp
SYKdDEYdo89xHZ9zzo0P9R+bDbWXS1pdXnNkz3NoqFYpvPF8Xxn3133YzeWTLWwc
xcpGku7bcQfd9brfxfjm+eTXRHKPRpRTF9n3wJCMiXUhfzzNJXc9bHTpH4dpg0VW
AvUEBYvxpqy/ISXcNajGSgCQR7CzBWzICVY6MTDKrqe76dxkgQMbdwVjUsrE3ii6
pgR6XdHRdlbbMIMZ38xmQ5fKME1pRUiLgh6XBA46IU+g+/7qnSNEBIBH0g+htOc6
6Qv2AGxdJcDn8pGpgUC0SosBNUD+ZcmFaNMIDvg0hF9EUSoV1GKBKuKtsRaey/7/
9PFvlf7qUxZWTNaY0Y3Qj6vDM0PO+HdNIa+B7mjeZG4HKd9UACWCT4anWU5aBxQ9
Yc0mVL+e/A8oZ8OCj/4pDCqFI2Y0LhmdYCu86ZQKdS0mX4SPWeZH5eWA7u8/VCtZ
3y6Ea5I3tp5nNS+hbbkGTGjlDhG83JkNJAAubHeQ5lVcy+BSZnUklKX8opiFBp+a
QaWZzcFhZLT/tGE6xjHRzEaY5DPwxN+7X7j8qp1Bl6Pzrt9VquaVUVprRc/Qsxuw
nU5czwygdd31Bk9/8IGKI7JKrft7Z/cPXsuQsKCE5yIYAyzNripJ/j1M7ta8JYrS
Ky2pAMy8tdciBa5pUN9qgpg0l9pGIcjtZ1i9OUgjJ0ClZXMB3f468+xhgvfHzq0x
MNDWYLzFIx9mdEcxWmfvWKWlVWACxE9eptWl1XTPmb5hHgdqNgOx5JDJkX/yyQQO
02YKDZSmEJULv5XIIqRastwFeQZYzPCLWH4+/2TOiuLaycwCCK4MKjzcQErYr5Xf
aYdpe/0F1DWl9zgGhHRgKwolBtBMXyweNl6uHV2sSCK28TZ3YpjdWbJ842VzvHwv
/PWFxKcbydsHb3f9rfm3rxkpMICDXyD23FrZm0HoM1A7juuqOt4MjFIIZiYwCJzU
qNXCEParor7lO76GIL/fmYdlLijrPjzT0cfLqgCPP1QOrF+ebuI3JRtnXkeLQxGE
CMRdfbkfXTHuCtqRTBOEJt1VsOD9St1WM3zGX1nZBvuYP3WZhD6x+m5Ei5i2hIPN
VUBtV2EXxYPL9AES0+WMbnGu+APJVJK/I08q0qx2Y+MQ24Mlg2lu2awpQ4QWEt22
JmgNKqdLSnn2JUJ7zfle5YaIJb5EX/uFakyzoZgPhqDgUPp24lbCigv9vF+9DJu+
wILoZWSghmyv10x2eQ1rO6oXXAS7Q7ZTreHeOjaXqs3QTeR40HURCvx2IT3u+e6t
+crZTzWRqhssOAhxuvM42kVMQB8bIPlJsvRWBakOKX4rBp1nbe7qu9D9Eprzgtpl
fVmJUJDFufFHYVA0ww14XAtvX0Hnvvunn9AWvfzfSqIfOr8Ax/E1zjTqm0giNnS2
N8FTlfn4Li1WDy4Jfpd2F74jWirkQOnIyHy3OON2c95wlUDmMqg3pxvifMlniBeO
A8UAsrUrVwkptP3YzDo/IQXOa+EFC5G1LCGlKvtH3ZvulbJkeNTI5AtUiDT+Ixp/
jnN/Fal18wQGz8rhaZHVUDPlLl0QOwB0RuthVgplDWE9mu6oX9XBsGncV7FNloce
9JeLb6b81Q/XuA1zuopgwUny83nAtPjW/7gUJcgOAufKchv8jw2e0jBXPnlSDmqn
myIhwyAAr9i8EW78uNYqpzNu9s3TERxmwBfLUVnjk4hwfUv1W7sTfjeNoyiKMqn6
uIJyRVUxq+jB1EIvox9c6vGvpwG3NDil5VMYKRvmYwIP0f2I/7jkIwbM/ZqLZmoc
3qiNYMRg1P+MQcFvY3TrPQ8L9pkmhbXrLvjmj+CqyQqr+ouz4HX9m6F6VfZguk+7
LqDiw/2yIj3R6+l/p4Ck1hqgw1ASxFuRgsOJBDXk1mSPaiRpkj/HgyzjT2M9J9b1
0PZ61vYoR419oW15nqR+hBIPyk8kUMzP0ltH35ofhMvExnogvZHfTMqaaIw6CVho
z83NcjxNsFGY2BCR1cEKRR0YPUsHAjq4QgjuwMKs93jyfg3ndh1+KOcolhTkqk42
maIBIptxr54U8wCHdpmS8beltbWWx4LQ4Sy6ex1BTfZvayR/QRVrrbT9aQ/74o0b
AOHhn7kaIIp0CTjwCgpjbGoaPrduTHSI3gqxDwbzLNMsG1KgxMxTTrY98lsFYaS5
ILExZ+jUlDHID7oBrPHeHsipycuzJqmYqlKfzGkwqlcBEL/J08gHhueknk4RI8vl
czMeQAeuw43w0wNI3hjdMvYHj15IyjgS7eiCLQ3hinOKYv//ei12v+ofJ4bs/B5F
T6V9vg9OOn4ZfTrfUxG3kOc4xEbSn1rE+zxCqwn7jLMe2Ik2vZhiyn7QT51y+MQJ
Y1VngL1TN4w6sB9+C5zrieYgHY/p8aN21uTTdvJYBf2B4DXBJU0j8Jle+L3hmeAt
x7ftUIPU2GLbFufakShK/+giiJwDsn72Ostd8irFIIyo58m5oEBr4O4A0HV2ESPB
RZGaQCEd0/V+gYHHedkJ7W5vUh/GXk+8MuIc8uy1SOUdmd3QW3youPYQ3aMEmFot
wy+84rHcuL/6Y/6Z7OR002yibl5p9x9tmL7DVwRhMkM85b7lBGtq1TOvwt2RSe0h
4sN8cQzZwUplOj3HH9NYWxSNWaNXE4DHlo1xQAj4RXApBAApVRtuTWrKga06RMPE
KhaOKmkma07hzALUz9ImvGOA7pGBtrOxMOLCu67us7W/oIqxMx+CcBpZIy7sIB2A
/RV35DAnSTgiSRe16SFdaQyEV2+HP72meaMpGfrLIshKEPA8bSMe+dZFIjUYRFBv
J8F1SyZ9AfCUm53QIgZ60jzgvvRuxhjwPasZeOwnJGhkzskrqYUFwyELBqBFHVJu
amBsPL2E0u0448oFcBrW2sgK+X9+anS/mozM1pKT3VW2YF0sVBzVnje5p1+9o8bj
SEcGdsSLLJ17UlXH+qP+XTEAaz3VjhxX/IXIUwaExsaTmG5CJ7OCB0Nf7czojVWh
ZCkJL7fQD/iyCrlKvxHQpLlUsdZIFopJBMUFe0hRjAMtFtpR6ICqvDlxy5SNgc19
/KyRee/LQHemU/dqRgNaoFm4cjsAm+2CmXPCHzpOP1kkxNXv9UWN7KNtYCWq5Nwh
fD26iwkbLI+XCAfA8OOmZ5ZIBEhP440mIHcz2eWhPJEf2y6zCFMkOq8qQsfWS5ES
inO21xy2iMccC6MdkJrJvb433bIymRFfVGXjUMlcXqUwieRu1FSKnGHimop6VcaK
BWVWPsB1L5fvsEFOCoB+gnD4O15KrRuS4LyqEn0UDcVTOg1hJlAJxumpUJchr08V
yIOUugNgCu7Jrl+SOxIjEQXurzFZPUZGJpFtBBDkD17wSel85+iEnqFUP8YeDp61
d1gkzEa3VrKiEpCQ+W+XXK//3KcZ1c31dCUV9EYVRNgmLpHI0p6hxQ13aovoM/O+
ShdAzfJlVOUCnvmA/kuXslLtviCHDcolqgVcpD+x8W+DipAsnJjOl5HMhPWwDgIo
ulTpkDkfEf73GvqxpFoNknXTBwL+ppN14fQvZI9FjCTYdnye/CxwGguR1MKrhIsf
qKHLLUWdIDqDs7wPY4hzd6rTeI1AvotPp3leBSOW7E0ypLyoMFy3/83ewx6gBSNF
ZFqbyah2MNZmiyf5nvMdOgQ6fXAEI55VEDfbanedv4fTo+NFVPdQr5dH8mQosPNx
w+p+FauFOz0x9XogSnl6MnkG2qiknS2sBpDaOZ8WKtWm+tfnDMKiPxuO6GXo6KWT
Uo1bLLemyopCZ/PlY2BlKb/Tr+DGcE3TKTAstnTCbIecTF1Da8LTikvc4miSIi3K
2SnO7ftbZWuOSZcn/6/xVlH3mNiz3wvou3Xj8U4W2X52c/VGn3Blp4DIzSvbfv+3
SLn9iKspiv2AClBHQ0z3/hdVBTNYxisIMP5FgRtlIVE7uBnypOkptF38xNxHs9fE
cfdcvoufBMlCEEzag9Qj6QC8a3u44BMH75CfmkxHcfP1w91O50Yk0INUQOo9Vq7R
U/qrenYpKM9D2A4YKiHce2hM9+uLZVPM6+rLxvIglFt9wcrbq59pwb/sJwSn6CGh
BVYBOKDUf5fPUBC4m6uIZc3QLIwsmIz4HXTZrl2s3khzRkk5/zk9G/5czEBIp6Lh
Jgs5NP4bpCd9fw4VM1XE9xX05PyxeKKouFBZSVuqdyUX98w3qrM0aTn1EUrSzzkW
YWl9Vol5Bz1wOQAaDOwo5N+E0RvAdDPt+oQQRUk7AmhN81SW6XeEWYy7e+LQH04i
7Rd1Qs0s5hw+UG+szdpYQ1lzQBCkg3gA7B3lAo/TVTrPdZlrlDBAdCRGOU3P1Npb
xB+OoMfwp3CQhDtLUmf+zjdjJfYeguJMLNxjKcrfNu0q+dNImQs8E9vMnqqIkCvr
PSKzWtELCjOmH59BzzDlYnQ9t2pEjBi7VKH7ZCBrrrwH8X0Smgl2YBSPV9dNuvcR
lUwl1fZl+4Ae3H8X3FtiNm2mzEMthf9vS4c9su0hZr0tHhHTWyJDbS0vFFqQfJ9l
7qKs+xglN1YvuwenLI2bNQZECDcL1EWVujWS9xGl+em8wDiojVf9jFtPPpwxcFjT
LL1xFsWwCwwbXmc/tybTKBlnYG4PHqLgw65IILHjveIdqDVL0zkWeMxUciZc6mOb
I+eQ1eJAOynoD/VTKLRJztiaqAVpg886dlh+4optL84sESmD3m9Vyn1h2k14a/r4
CaNSMJAVTomDILp3yqErxWDEcRDiTZL5X8OjxMNfKtKXErxZ2PpeX8wVcNNHu5V5
JOIPt99e9nyzY6ZUxomThvpuF0kh+55oGFd9bEGtvpWzsg2TIGS9wSaeBbzMo1St
TWIApsyRpPuqPBSbBhKBQbG4mqCtzku6OgzWAOW+KNfAee1TU0zF9k+antnFsNI8
rWwjMWqcxyvULqdNkJzo2gmsbeIuC+YCKJnzQ8vHyliZEzOeoDIRp71GWTUVr5fN
m8+92+oz4VSFSYnDUGfsHzq9D0MQyj1wpyA94n7vNeqhenI3rlq+KjKyzgCBJl9J
Bp3CpvmecI16EjQ9T0KtoRJKv4oZW8DRbt7gd++gDzgRXGsFHU1iy90+okXLvHpt
RmnpV8qXariY+eVESPzIRWLZ6RwL9XhgotXuEUSfVT5z4jcTllbR4MV9OhbXwN8K
LErrn6+Nr7iBvBC5LIgmKitH989o3FDzHZsCxT839ixfKEU+GKM7wHSLwPKwVqqe
28+k4X/S2U/UpWfPj+M7K9dJRzJdKPh+WnFjVERdn2DZUhIslmIo40O9BUx+QId6
0xF1m/55YKJmW5jGyC2C84Z8q2zZ91eUPj5C9mE0dY7ukPkS64zn0q4cACti3DzP
iSuYRdJtuy05pnsMu8rqhViHOIdTnkarCc+uVicNcuSTG9BNJxVXSj0cP0YYvx7V
BPtCRjwqsun+ImzPdWgQUoY+90DfFSp5ePX48iqpFDGOflWzUVyiibZpVLFEz/IZ
YoIBUuNj1QDGt7xZ935Nbh++lB4IogQMMByGkhWOWSlQtsu07966w3Hhaddnfb5s
ixE3e0ahH3fKV3ViHYBVIT8eSfbWDVjoo0fFS3pPa9ciEaAGGEqiN8baVHsiuFC5
g9GuBAk2AIxQDrcihUIXdcZqdPIs7kupLYNczoQLLfPGnqmuKUvBVwqLM649ph56
Tg0CuQRRX2KkQ1Tfe34ZGXXC+OzaDUSHO1zM+SYUD562ftD+YNg7V8LgBDEz2Eqw
pkevn56x2Qyna5J3Os0RcXcSGBVAPsWpD+RKeCE/9RxJHo4zY/dk2bY4knx17HFi
b8ZoWYbwDmaJVO+FrG01d/X8PcjTr9ESbYZRH+XMdHJBNa1EF5gotOr29O4wpDVX
oyE3Yz1ATBqemEGx3fC8UhsjlZbvKxsRiFwHNykUAOzXxxsC91dizxRLl9DeVI11
GFpzGdJGqtFn6y/mLrpR94wj/JvjScMLqHvBASuEjMc0PxKEJcAtVwbX5R1eWgl8
YTGOXKhpk5Mo/sroa8Yd8GtNPzxCPiMaw6k1w1EW8SRlsqtLw3akSpVOAHI5TAFQ
VfBBxS2Yyk9/7N0scBVlo5fS69Q2ankjVtnsStyc427hMKhd72NczINl+Ym77tIQ
KKx6e5CkLXEcnaGCFtJsL84BF37eEUBa4u0+2eHOcfNUDT13dDyGPdO9BGAbiL/Q
iU0ywAaPdE9PCaGhXqojSfPj7sxqZN4DFRHslz50aTSQIPfNTgxcDkCM7PH4uBLa
mfoVNu1jmCJI+IVaHtBFX7R3nk5PMbi6cZCrfKmTC0ia5FNex79i3sdhAWzei6of
NXlEeIhR9nAbCTbF4pahti2sQpqnlPi9p4HqcmNGhGE=
`pragma protect end_protected
