`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XKNLtFj8yUv9DTR5Nbd7+bTykAZsfCSMMCGsxh6RrZcV2ZH5eH/kWl2zQy/a86/s
MZ8QveTZOhArYb8OAaNaOzqEMYA0SbR/5Th93eZoGUhw0781S2REJuPLo1ZaVO3E
8kzKtob3Eb4SRn+/6+n7zj2VkP2arXQwQVRi6Fd3zuQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5408)
dR0FxD7W6LqLgEU28s/uaZPe60J9IbvR3fjM1ThmPnJiriVcyA0k5VHclgTF1xCp
aS9Ble+kURHxHSW44caONWmMOWFbRbMx6US/Xww+A5TlwHexpJD7s9Xz5qIOiWve
hZMzMopTUqTeVXE0B3dpVBsPeRj6LZyN18ND+34o/LjhhuaY0aXmH+32XR/I/mYW
BKKNyauiztvVXK4wtkRUlM1WceM5X3TGq3k3GoMzc/JUeIdtJvW+z+THd4nxCXlh
8gA3q1LcsGEsDLrDgoCuoXavuhHBIZUyIIkuvfa4siT2eWi3p+rxxoOnbMXdM87W
XOPqP9nr1n+Ql+r2Sj6sn2FXMqX5UQIzOVu51wDNsw1s3h+sTrWktOTEqo1yOoEe
TfZb2i2rT2BuAfYla5NY0nSiAr8Fp6cR7YeWIz1QPbUlvl3XnxcPZpWjCzrfc3Yp
xpXXM5UnN6xBaYRusgvaETXdpZtXcOBtKeGNgxG2Q094Rj7opd9tjOy/C9YOO3Wg
QsiIGqQAe4A4dDoE2GHhsY4u/ibcvCFrJ1Q/6VyZljgTMXRx7wu+Tr/cjvnSr/3F
J2h3+/2Ln3Zb4vyKiV9jWOW0OOWIzslO9DdF7NvTTlnn3ScLZtzt7XzY/uHzHIAm
VFqvWz7LLGWF+/02zfrxNVQKC0LeQJF4ZQ8/3UGk0lCz+trlnYovmGHnMX1fXq+r
vMKWDGgVawL5m1A/gwsPLr3pGJbmFXp1gWCBRcdK9IDfCflV3RPe2RK2QBJRBn/0
C9lBXAcMPoaN5bCJQ/65yFDjk6EVRDqEV9uRWv8Mb4rFagrFco6cl/c5AwygSyxw
eEF+K7PWTQTMJZxGG6xzhuhLTO35yZVyBXD8PNzmgG3AShCRbAHU22SfJ/zp/Do0
KEMMSjrqynAqXiXGZJfQiNbtoPR/gDSWaAHUcYCpJWFtxUT5QhUMnvnNxHzNLLnw
jPVhZg82lTRySIt9GDh+WDXTBIqrW+LDKxpQJ75AuMFbywEpuCm1y41LFwEDDsh0
EYy7zavx40+AV+FGQoKRgUKaPHuZWDRK0W/asDNlN16fxIPJrYrgRIHqLdFFDdmj
+gocHmu4A3sxfQLiHHArg3OJ1vXR+bUZ1++DbD8kLqbWZFdHMtcatKoVF/8yGdaK
ZYaSZ8jKojvYJyc0Ty8wvIMv4qDmtqFJR54iygl25rpimUNN1Xn7sLC5m0HyTKET
/ZwePUni/wj9qol4VH9e2w64RepdO+n255fio1Vbtp+EaN9qzo6D9XGQGrZQ3Z7w
PMOhcuLty0IpvODSDyVYYC+zKVhrHeSYq0fopaCj0FK8qcXOLJW1TJM6eQ0zpWK2
8ARwyN/F0XZLUc2jVuqJdw6JtdZsCO+WqBQvSXOC3L8fylGcfG+X8dDzirJCbjAh
uuf07ur/4RIU0JThdReYPWTgUQnRSg6pp8Z3jmGvaB3eQYlY8k3j9P9/FShLFsey
VYewAxenUvAUgsItgd3cC64YFZ3xdaW20aKke571OPE+eE9JsMIAEWTph2Vd5UqQ
okoDcW6l1qIx92WR3OBeEHOFPETSEhQ+rdrvKa9CQD3Xf19cvXQAZo4SS4GrXD0t
+Ba434O8pFBBq8amwtmVp6P2Ybtpi9dIEjba6l1XH2lZW1UxFTX3EtmeyCwFeZoc
X/zRZH3p7QblOCidyj6VG21nn0WOUvF/lQabrU6hPB6FhazRRd0BHot3Nck2Eb/x
dz0j4ywdgumEC53T+HSeCNdfSSrfU/4teu0aYP3ikNEt9pBN9kmpxaY9xEpFqUyc
wpYuwS4wSVX3T0OBTYfx3iVUo80S4odwNZ7/lb+x1qgh0+xX3wuLeBgNuR7SWOKd
f1AH5pWsruLbe+SM9GWIFJiCJ9U8twSc/SbOKyBa56Wf5cPCxBKK5Vtx2xdPNOmS
rErGMDxT/RUYZ6rksmSw9+N+yTwwWJOh8Aw+UoL3zX83sU6UIk9xlnBvaQopCxgE
VOVEwC3M1IuH5Yss2hl4Fq/01o1ohno3TtvFYROQ92NqStAu4LwFp4VrKgyIM7vX
8CXB/1BCokF4ijFRr9uYfSbQg5clc/bd/OcR6u0K4WFgz7zXfkzRlBjiOWdLn2WI
xeMRAd+N2bMmJmodebTb289REkd0Z7RjfGJuIobck88gcoYjJkLCA9KrrjXE4pqG
Jcf+PbQhZhCzMTdcEmFVmCbwzfnQ2WH2q9j1u9Qd2Q+RtJIpR9OuX9DC7GsyZvKY
G1I3fL6tGmXQXXcMPoI7hFWtGgwb0KGEVsdDBdvd4cOa7WL3AUcD0Kctb+8nbHa7
vzb2ZO3hRTpP/ll4yu4S0JghXAUiDxv8nKpgb/kGaFrjW+0mXr54UVvqg+7d75H1
QDsD8IP1KpehZkxbEOsU5MEQbwYl5CNBB/p8FPLvIIWB8rYnBz5Ah22kmTFIzYNR
ZeCuwD9vUnZezg0swWOAqdFTfi2qBVwvAMT+uc6ECUK7DXjX4j3NApQ7PIiKsHJs
PjnI+ixvt2lVC+QpYf3gZf+mvc/pzl3H1zC9AVPA3zNeTjC5sy01wY7ElbaO5swW
Fnw1WCJr672Tk6vTYdVNZqNjYyLKY8KEC8ZrTML0QdyDN+pNEhr8u66Wwv4lLkk3
yuWjIHfvYiRIRCLGjlTbP3dQvzMZRQbzJ2mw9UO6HO+m/t6jSVeX96Jn5XReKRoe
pXXq3oZAgXpf8XbVnzEpwMW4xZQ4ANb+l5Y7YtOvH26H6KUdfj3N0KYLGfIdSI1S
a3yBbExXPgt6IohwW4wi0wwHJ0PlMSGaoewpo+PLMYkC/wensUUMpGQ4euHbJ7AX
9x1iVGpYGtDwD9seGFpSF40vr2c23s7SO+IKAtEME+LDCqbCBv0BcSV1hta9u4Lk
1uWW5xqXCDrgs+2TO+yyi3isAfavCKLWPYxIVgzMD4XW+wix4aRiwEfcyDWLkcmW
T0hANb/krwleln/X3COjJSJpSHvey5OJGr+d85T34mc8fx5w8WzUuiwujMSzC/WO
a2t/ii3+jqY3zpZzjFic9ZJ6F4wUdDCko/80eZvNPCp1alML3nm5joXheePds3/8
vkXYvZjQ+BM9Y/EYwu8jvTLVzJlGaJniVkgE8heK8cp1nd+qIqkPhHKM5p8P0bkG
4BqLS/sebLqQkZGinL04woglPVkzPNZYSL/Ckf08AFVRvVfvIipEkFa+UMpsJAcg
N8LTdwmj7WsgsEgoUa0xge5rZfj8o7KohyeSkkRrGWzFPUr4FlyG/eE9NedaS3Qq
KB4CXOPtV0xYVyfxrLfktAg89tGtAoctTXttu6wdI1+f2dtuE4aLMDzcqlcSTsXU
tcED4DRmMc61pgx18isn8xJiYv6aiiKlDQqW1BJy8RSk/RT1RmDbk0RnYX+j7j3Z
3SffsLBv5QN6lm22b5MxuYJvkTjAofQYAgrDQU41cHvGW5awJXl4KHEbWWf+xNh6
Yso3/4AwIuUG9Tvjyoq94R7hwopXiz3DAMsqI+hnaXx3UjV0DwJjVl6lcavwufdn
UxMWtpG+TBrLmJYKMh6J1wu85jORP+PZw+kGRJb4lEBx4Lb9pnamlRRPVfRG1PAk
FcQqYZ6mOdIhlCROeCAgHWeLPGFEXRc9Ed4pZlN3y04UK8xCRnEvbkrKhNnxhuXN
yMlcF7mKcsRf8BGSdzZm+eiDRxG+Ix71UAycgqJ1JllHlT4cNDRDkWVlSjOhlh4V
E8l/x2LGedQK1VAcvbTUcGi9iE6yZZ4Jetxt6p5rXrNofY5DRt3fjon6E7pbDtCP
rE/gYTyD7yTNF8bKV6JDUCCzTlHxAJwwOJpKCDTauw5UP8sl68CXB9b7L0+QwOYc
vVQLnbo8r2lnCa8Tjsb4APFG1/uf9aE0zqy0EU4rWuRRPDc80Q73a4Jdfe08sGYZ
wcQcjOrI7FOguSux1HhrJUxVd2rgj4F0L0WACvfHylUhzwsW+7DKl2XvXtSAdAvZ
h4JadZ5Uy/g77TtxEdukRq1tDdSGHfwEcUtvLEoaXSs3RDsdIPB8fDCKIMFGctq9
ovQNUWjq8eO2wZXEuTUBi4on7FBAvtkHOQN7y1FT8PJM9pXZXOInJf5tt/82/1m7
uE6CIGBNekuuCC8vcIAjiaUcyLfHDUhto6hNgNBjddDkmXuF9Z8og46F2Gqxt1Dz
iHd3C8bZK7iST5ikhGcdUaGqdXMMFaeJ8kwlxeIHK5WPsz2EWat0SP5BKENkiYEA
Rvbze8dp/1qiceCdH2bFAwEryoByk03u/ue3uUd4M5i3p+bbCRie0hsqz9owfE0f
Y6A/O5sKK/XEEa/71E9MdhM8JicTfJgqNw7gCVR5qCvTTsSQs/SD/PxC6X/ItZqE
G1XQeuFoBclNpmYGv52MXcA6uRThofTPbavc1CpYsZ4zkN7FYYIWmCKwyXdqm1sK
rJH671eepq7Sx02nuADHHWBuc68THnOrM1IcbfkSUhlJkkjkDH+JKZY7A3p5xnux
aaU9JHCj2H/zcbjHtfNESTXJurn5eYdYjaKKt41zqE7MlGRUAUZ1ocydhJkX3fdB
OH910JhzRmzAYpqKiGaafYoxOQJB06ld3cKDpljWBGPpXbmHiH7ZN8gF1t0gX2SK
4zoCXwQfCFVnHKTn3vvTuY8IwNGbBSOjKTPsGndhpLTwNQnWrDzv59MApXZcK7kF
l+Kx9um4p5UhqILR+QPZPkfAENd7e6l5Nq0jCAU7cM/6BgAgPTsp9yE9WXAji4Q7
VBpxkzH+d8m4/XJmWOI4uSMUxdCYhTTgmCotZ3pWxInn5wu8wby8n9pAdpJ5jxEQ
Jocr9UmtIa+/8bs6juDOSGGxcgsLwpUdhmJNL4qwVazwkHYOTodG++4zraW4NuV9
RrTcITDQSgWT2T/URkgooc6z9ae+T0BbCMJBv32y41P8laVrnxZlRaZvFXupIksx
lgG/uJ/rCbDO1te4t6VEXRLDy6bP9j8aOt+6nhQF1UIfyx3iKfYV+KGTjV9Y264W
CbmItbj9Rd0dvGDeqztGQ09nFw7xoFrvI3mvt2EJ1HRXnVgJHqbuXhpSryQZPq5n
NkBYudESOmMpPZeBSPhAN5xwqNKocqymrzZtHTp7OsUjCYqprPjU12F89I2FEE0c
1kVBDXHBxXNdlQtPIEZyniFQiIwmN3cCQ2/ilc56BaRxFOLOzaRFDhNqNVqr54KE
kKFeyR5lv43Dav4J7zkwY2NrXTG3bTANh9C9C73HVclEQBc1IzXuN2cQ6KensBDU
r6yVZQoCjg6dBXdb232fkWXS2b9b7b7rj6N0TB0OdNd6keEUM8Qr9FQj2JgFCnCj
ewRqIRBWjW8ahYAX2prUWrgb7ucNdlPOMV37P2mTI8kcBgGIFzBjUmPN9Eadgo3g
7FyQI/Aoam5O8cWTUIwNPuSh9OnEeYf81yHlt4jV4MBvSih/J8vXV6bHmhuQuBu+
PwcSgf01Stuc22/JRtKGSWqdKLPflFwi7APDCJ/Qv71F/CV2mtTfiF8vaYtnonSw
vYRwCPZjI2GDTF6cmuI/FhLBvaMmfqsQOYnYZZL7LxXfGkPJC+Ek5Ho6QY1aG0sb
WtVr6SHD4Df1RwISJt2BGmzEScoedQvO2WE8zyHx4BiT5Cfj4U+X1yqfZzBaRgqq
naGazo8tm3fNTZhJKnVamqQAqbRF6UMw2Nsn65TU8ZyIL+mjBYxA6GZVdunLKzy8
EO9n6KlLFF3+V62tRyW0JpgywTUo4ZBgxbBSYzAaWEt2ztr59xkmU7olc2jgxKiG
CzW3O3IC4uPPtoZ4AVHHlxFiImJFhC4OVsgrD/Jones78jeuVJVmh6UGDuTQjYGD
23IUr/fUp6l72bhDQYXQnZY58wD05tydKkgJFDHsqMrOZSu45T1X23lxJcWr7E20
ME2/LEDg5clxZ2moJNl0eQeEO+eh1naQGiTZej871Wwv6Oa1QF9w8VS61RDaozjc
pHU861uW3btdO2a8N6J4+N26MNz9chjmTigUpyq50cIcVi64gmop+71Qp2SMKgWU
5BoKSO2n2fNz2FgFWv8Jur1GqEiEVlBi1ds6fXGzTnobPK4BJKK/B4XYPKmDM6r6
7GtAfkGn4SwEPU17AFDKMxx1nJPKdH+s5+GjuZDbLB+MHhNY93mkz5Ww82Ywsfii
qoLSVCpMG/aOhU78qIRJ1HkQEkshsUJXdAg/2tUGE2SOzdFHJ50+mKeG3A/KvghA
0QZOositgvfFTBIsxWh0WbOobNLXYc+FklaIiOrrUKnQAkniY/MGLRRPFy5/m5et
RotFmeCj1fQ8WDAktB820pN/1K+aEtiz2+BZDwpxeAppYLSvh4TIrw1azf3wQ3xh
XncNw3MQQSndHaroHIwduu68PqDre7HVJoMpUUC7pyUtdi1sYnl0LgjFoKSx4i1B
OwsW5cxlHHZVphDD4FE9VVj3rQRGrL2auTZfbGZWszHg8r1mGFhsg5hc0Cjdgc7N
FViB9BI7YJbqk5Tz000/hnd2m6sbU9HJwqraaC2VH5nNvsUauxtV6pZdBXjTmZ6D
Yj3NV6JVR8XQwoftlAEDnAona2iBgPJiPg3c9IHbPXWKT2GwJEd2ojiCxW5E3012
T2w/gNbUdTEXHlRB8ooPr4clwVj2bpne9WKA9z4BIArm7hqiwgaYIR2aB4CbvJ50
2CdlG0Yjd1KjJf8FLeg3rTJUkMz05Gc0hk+MNmQD5dvHXlVrb5d/H9YZpwrslerb
VTb+OXIFo3W9CVmijbM3yIART0DO62WE+/0w0iyKJ2XM5a8RC0I3NdF9WCxEE4xc
kDTcmorwrkLhB1YmFMHD00eC1br+ESd0CBeevLHWtladruEHNX/OkaUddChNQVQQ
9zMbUndXFEJXIyiowRZW80oFOWMdWBv0v4QCiD1iJPJh99rkWQmU285UwqA/x3T6
kDe0ND+MiK4evk9vejmsDxWl6nxDibibYGGhvelclGeMcuL1yHuqbYkrEcCqJdKA
vCJq0S8zz9XiAiIDf4Tq+n2n8wJOgkM0iCpud5BbeGNOw2bUC2Oc1sNWdR7HwU5o
3XX7rqADoGwbz/r+9Lp6sZSDJ5U/lpqmI691iHJGHe8EcHHWlLFkkFDu8zgJPlGt
QhfKM6UlyGzV3u8Tl/Y8kJr9kjEBt6JdsgWfJzWG1cgXZZWzJg3sHy2IUJ1fEAC1
rwc3mhemEti516qApXW8tq3VlHlO88m/3GUyRzLlCLI=
`pragma protect end_protected
