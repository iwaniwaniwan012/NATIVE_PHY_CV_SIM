`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ue40a2UdOUYXNBsUusg9QRnsp6yJGIY1Lav8cIYMqaIQPcEV7/JmPo6BYV4cqzUN
lNDXKtovVwFfwRbCjXpQh3y/noVqa3xePnqOk69Ot/1JuGibgEyyHBiJXgZCxuCB
qH5Naj6Qkmdxomxwemos/gwTe5Zeb3HdpOTsKD9xaLg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21904)
sXpE0CCGxk0XekY22Qm/Y/YmUwzqEIYXms1PRncTQjiAAsxcKfPa8sPlTnKmW7mt
brk0xUQoRpLI78HYB0x108JDJ9sn2f/hJDwaInO3Xpd8tfB/h6mOrHaT2HPyhEg7
Tuhd4bcT5VgU/FaY/Drsf+TqsCrGJILwRCVGUsU60EqgMq2OoFqEsfIUOpaGgFLW
GXMesyQlgX496e4KQTnHBjf0eeky/zga16Cmt63Y3iARX9rj0Ar4OuOFJGUtF0Yd
9h6aPjiBEWzntr1elwIVMPbPsxMKakXr4hfeHQDtyPI/g+P5xR+sHR+r5T7hotjf
Lds7s+cz0fALmpDFqHXJKqfNYvK+tH/felsen00ToQ9tHOKHEDV7NRxPpQQO6lA2
VkEpn44O7ypVgfC+sKGWtAN8S80XmAcYEUUpgr2xW7/ZldmCliKtJa37u+vZqxOH
l3VqmCmctZdc7zLZodk3076mnLMl4IvFBC/+Qph1ir2OhZ+9I2d4riToAQ9GPrxk
pOxtCOvkUdM6/pFgRQ04xsyre4brdNraek1snRqAouFLrq8cIg/oAXAx5RopTZqM
tD+F2iEvAOmVglB94+ywEdWZM7JJydJehvCo+sAFTRm7bbdABH6fFjuxxUopuDv5
IyImV/rIaACCKHN2cDSeJEbTojNrc7dh31DiNU1bzfmdm/QwgoWMMCJ5ewH5kC0P
NiEiE1Z2h9YIh48C7F+MDc1OZmsR6xcoOlIhNsAQQ7y+/kcl/CtccfclE771VZn+
r0IZ9ioSfItt0isWM6mhuWycoV4TZgvJq+x83KmxUXhm6BuP4Eg4EI6BP65dKb3H
uw9NPpAkaSxv7XP9CbWbWKK8uy7GVBtA5FGKG5yjKqortm/qkpHhlaFseD3Pow/t
70Hp0U9Ze2GFfuhld7loYu1AoYNa1wmT5QCLgvTL5+w3uCUQrpQrmsGXHTO069b5
LDMap8V4nd8zm//eIat4J/XjhGpu9vKYokqMWxT8Wcm11NTHStl91GgrIuYpE90e
JStJNTZi5WJzQh94IOwdO6Lsf46MMeJS8tBdKjRIbn1lcbnwaleXEzX5a/6Ciy0A
sIggqO/uPyDU0OwHdIY9dsK3mR0Cv9S/d87uNG2SIQeB4eWSljkpI9VYoO4wxgB4
yAzWUvna+AHdHVGyXs35qyJdB8H3GwoMyuV6EiESyuq2V0AUwte+9VPoBqXlqZnK
TxznKMZKQFq0C4K9Kum7h1u9P3ytwerg/oSq5VkeBvXRuoTqG7ejCIfq023CHBnh
2fa4DTUYBJTWNaX3bsaMsgqiF7u5NXbo8r05sESq1XrmBg7uuLgtOm8B8RI3MDpb
Etz/tXR/96L/7NocviMwAPPWo1+RJxlyva8AqO+t0rU/E/UpwapYmA+3t0fDNMYA
A0vcBZ6FAGsKyNJDxYWgKV8zGL/sMv6s1hLtoWhyIA+Bz3orM/mrrI3GDwSwR8Mq
hRT9TiXQFZY+8YP5x57t2YvoJ/ax73lB7+lkXkdjX4rtfV7wrp+LJq6f2usRj/MG
WyAXITmnbS9Tmch/4tE1DdWaD1w14Cj23UFNczlT94bD48efliLp/i0DeBr/xhWF
YOccW0u2ZT83unQeJYk+CNnfPcvT4Vj9DcweL54KAvYZMp7iFw1wyUjwUD/qjD46
cO7EtsxGrltjZwkUl+U7yDf9mtxk+TND3nipJs713GbBiUGcf/PV/jQfG2cbqqwJ
iWWfXGDoMI64WIhRUV0F/1nG2rciQcSOuhwHmi/nlg2JA8HDfZwEWprDcGVi+OuP
mzIJUV+JyzB4EuWkOSK3tlYtqzu5mZyRvgitMwmosytZefOzEeIC4RWBFaqR8Cuc
2JQTM6OQbSmmKB9NrMFcfH19TYoNo/XFpSG9I713PAbd7Y+gLyUHFZ8O+IheGCNk
OOfh2AER2O0jZiZpNLoYgKZ5UEAlFdjXA7PzYdUUHcqoyROcLNtqwRQeAfSAoXsM
3VZzc9JAYSKgG/ldV7UiQqyodk5zs8DlOlI8M6CsyzW4ovkE4awGDvRFsS2FJ/1l
z1UHP82t05mvzz0L8KD0XFSwAKj85bhPvO+x69/mKkj7a15GXGuzeOJDE6hGec4l
gjw5GbpsB4en3/DK+UCvlCFoYV2YdTL1wxr/RYMmEg98OVEJwdZmXZgRfbooQ+cV
mHdqDGri18zn1vZeZ+8hQJ2qGjUuclNTG10VoyuefWp570YNIAH38xDJbgSYZN4a
pQhQ36+i8eN0wIyUwsXIhrWzmrG8bsHx8BwVMPRHG5JQbVw0wEGHR5uPSjU6Devd
g9TO71BeZyTIjANyY8SIH/aFMAfM/nFul93fkZHVZvu7JqlXeHikCi7I/OLboMEK
T4wcZbsQcAZSyMn5uQdY2s3XnnAcBlzC9ckT5P9m9N5tKZ71g2zxoMXytDKUCVUB
eOgxKEI3hZ4Rk6rDs5H8C4Xv/qxvyijnjIkJ3gebE2Y4lRrTu7VvICeE0yThsuu1
CGKPgh+LEnI8E11hUUQyYsoSiUPxiu5PpoAjZm76iM/EvLT5UPAoeev5Hr4zEma9
K+CC3j69wZPQmUuadkrVnzUR8eZrGwRJT7blns3lJxV9Zd42wEjX9mRYvD0m5J92
zS7voFyAAOeBJZlwkhF3gKBlpRsvUD6JKbKSjWzXUEKN449xxpVM0LOB7Kbyur3C
voN3mWKpJoDp0kxwXSPpzxp1uIMgwk1TxdlmzkD1ZZ+BRw5jTB/GXB05lZh9fuVw
S3jRjr98BYR9AWK+05PCa/GupCnVbQGTrMWfx9Xeo0y9iNO0QaGgUKJ7q8vIUs8m
/rCH7JY1zL3a8pNyAK2PI5K55xqUPLzNTklwGA75MLQEb0ACi7hQa1TA4X6aKDiG
3V+OzlccOwfNcT6n1JZfRhTefOHmi+qqrqG3fGI9T8MPdUTaptVegIxwaoeP+BWU
WZ3hDJJ5sj4aUJA0umUXt5PQbzLHw3jp7sGYHiMayg3Ub8SOxHGgk9EILkYRsURY
UZIt630vgRMPrk63OMeMaiJWt04Kec3jEFHo96eogQJbLiFlwfYPOu+j55hMrEF0
axZNrrZaeGoBrZG6wLVCOAeOXrspPm0snHDBvOn/fJjW04Phut9G6FV5GTRRIycm
q5fKMSMxk6cUlv9IfIWBa+CE4naP+cSoxuFWlvxr5A3ZJT+a2Ex561At+1TFwuQ2
vWwfvXO5pfqCxaQJOkA+PkA0qOIiIa5cuVWz78NEaNikxVrx4VZ8kxvXvNWtf48Y
1I1ABtv+DqPEVcRohyjhd/d351YxiD3iljSpIpQiuqRNcl004UMXz54c865iK2Hq
PplLk+4jibWMBUSf+TPjdYXeH6lwp+ZGO38N3nqcwKyWKDZkBhy6952k2fN/FEPy
c6qvsUHBug98FBdunJwJUr6WPecMIyOgJPvV4z5k9WUn6p+kloL60DmR4fsjiitr
R5iHMf1+KYwkUTOb2eg7Z5Ynu7iI7qY9fAeUjdCmhfXjH8jfLydfgdKLCtanxqCA
W9gMcuwcEWkpLdAv+utxftZHWuTfUMyAIAB6EBm3asPF3qK1RZ+BQ86tI+AK/SQ8
K/okiSm/0K2OjiOhUFZ24ONDXoFY/QTI5GRAnCBQNYvKp0ng6v3X1LNCfQiY5Gfd
OwnKQPqgCgVvAxQWSCMRDc87TdUugcbgkhc5eKFs5OXvHvieYvW3Po4L7lA9KdYg
cA8QyJO0nkGZkmdHTEu6GVXGsTpeo3X1X7jnJRmbf0LEsVr5L9PiN0ZPmnsgCqYd
eZmVd/VAxM6GHJvJuRLfuhCFNsBHDpMJI7MMF9GkxiFkPAkWNakOmNUr44PRneYe
VKOuqt7cA+HAL9zHMDxkqGG0aGNiW68kNpC0plAoBaA5FfbdhhrRy/1wQvUbVPir
rQkLkhdIY3rbHGeZvZv24i4BEFryQL1U61nLjEjmiN2zhVlpovc9HdL6SNMiR3fS
SRhaC+YepZx4kuubFXbtiHsOZUlQZRwEh/i8DTyo83wVZGje3fNJnf2wdAfSohy4
Qp/rLKpa3nd48hgaAjl2aZavp68NOxxg/6Bbmj4uqTRZUsPPtsYsc9aUwqB3peLj
3UzubgbI8tqrvW1gr7gLDKYgwGBgqqkRtjKAu2h6HmaXiSR3h3GIlYIoaZ1ler/y
RrbQ3j1TWM1NiMASA8FJJ7GnM+5QeP6kWZ10NOg4juqRLqNJ3vei7bPmCelaurbs
1ZxDvSoRaTlvto2xL19xwbrPT9sYmwmPTX/VRViUPNBVwQa7T68AIAtMVCaj90lK
9HKlx4DbANtUPgxmOwYaHz0rZkiEQQE/1ec776RdJcA/Xjcnxgl1a6eKOjlimn2m
RQMhZORtZWOy17SVqcBOdmORAkaUhea8qDeqc4OsQ3V0bpHfykQPa595vmEdc5tP
4OiCbr6N0V4WMY3Bo9UNwXXOra1OUe/+XLqO3RmAaENq4qIfbnkBalRXgbxI8vdR
yTFjIYwFqLTF6uEFZGnk72kTJut4IMk+wEBOo09rfSrJrFAogIDkbAj0L0aX0QG4
gycxnhyM214KWAc3Tdnnl3GRda1f/1fst2YqsaKTW7nraRfZc63aQ9IC2uyyJUv6
+Zsl7g7sWWmJ7dMs8nHMxcqd1R16EOSxgD/8qRKoP8XfUJ9faBxH91K5BwB+peP3
dDtzAn+adCNotdQ0+im11AsJm7GBs9XJcf8CoPTmvWMnuHrRWLdJeJadzUpZVT02
jl1TalNW2AzBqQpJTCa4zD6pixmS9ucRQJfAG1Bf3G8m/m9MY3t6wWsr4/M5Uj+p
2DdznfUSwBLCtQa1t6JWLU4RSvQMo2QlzulKFwIXeytzLGJPF1E6W8MaM3b/pBC+
rxsxJP065LleA9IVcVjz12obovdkJUekfqUG+ScwsYvibhBrJ2At3LmwEbMIGfJc
JvTUaGfIehDUszMG5sBuu00F1QCHwANH8yR8SKqb7d1mb0oeGaeEBc1kIiDKqu5B
rPV1S/J3DiJjKrWT07jlYAtwgeGbHcEVzTZeS26sbEqcCtZWlmJSsSuZ4wLV4Pa0
9YOyyuEbRpU1PVdoVhEFvsD8BG/sRihKF4s4a7s241O6y1gZE59oTEXT2YsY9e8x
SI6Tzivi3rM6UxPoFeIkYykTgnZWdS1eb4FxA2PRVOkHyLysYdsNI5YyLamiJo8Q
tCpjw+KGV3nbwhg0pe6hqFf0J55q/mdhErANj+RoKrOXk4YtS9jXp777jSVrlfip
v7/hDSrWGoFeW9aYbhMWLWtXnws2B5B+38DgJWDmVKiMzBfcXohI5gpNzhMZx7sI
n0UDa5Vtc6fizCNR5t+NzlUM0hOMvU5jM449sBPxz01zTnsGx7xihb/63VL/+XUQ
FYq88Y7GebA0qU0oGaBW7loKR8Ic8pqZ+2qkwHYL4iTU22dctytwjKzJ2Vc2wlki
GdtKBZ41KQ9fOjpCnI2bD0Wjocq+j+Rpgt60xcBNvj8M6G9g1lrNbj+kCnxUNkBQ
VBA5Q+hHyUo84PlCcieEe1bjbFqRMIGKUAp7U6JTArkVP2nPOTKCLZGr+bfy8nU0
UqG1CYz4+49Lsbn2RNUnLjN7mak8u57aRY/ExAurkIai1bXftAmBYhOe19CroXvV
8/rMr+5jP/jd2qs702vz+6sXZdYUYYYlG7I4wlZqQP/opqUW2ryMxbe3h1vQzZ7q
hamWWq9etgNXfpUqveM1ssjLURxjkR91qC7eA172rOQQEXhUQ9cLItb+ntmVMkFm
lxpLttB8P66S5WP7GnHqEJC8GMPW80CuRCEHNKhzugDwWLk6pU44xNkP9Rkujw+P
fl3TSu4B1vo36uqDGk4o2X3ibS4TlaQMoSPoxdP8Hh/gD/XDAB74Q5TrAVwKNS3C
8XaTSDxSPpVawdg/r/hvs/eIk+NTkkv62em3YfL1gR5bPOv/euEs0Wnd/NFHPeZ6
Gbaw/mDzYEkkfud1GP74y0yJ/MoIi817JY7kMr7z3phzWqCFmYTZHx3Kz6q5XFkX
hYGwNN7RsjoXyIkq6lfK7IqVrHbnRS9dRSIw9y4IhaDBiOKx3dCle3SN1iQryRpY
NUI2det+FAADohBBEZMZ8qJ155xyd/JsIWgmWaHGi1LYCkrbhAEUaPYlpz8yGdYl
D2YFed+5ZzB2oKHD4gekNKbdQCPHru1srE+q6IlZCmzei2cwahejGGCwFwwLUS1T
XDtziNzYH7GB5T350YSt6u2AIPGlhBTmn6mqeQcmjd5cBK2FrdTIUyH2SteTxH4u
3nLyr0pMgc8odu1ImNVYERpiRwqNcAAo7rIDX0iKyIMRSqpVJRYPSIdAwd1jhZih
ifOX+rScghwOSfly+QjSiOKwmBy/vIp88Q3M/jKNKDAIe8oYj5T2bik3cdypd1sC
eVgX8yAniOgKZB4mTAvPSX8JYXm4NHw10iIFjicl3el1ps0Rm+iyJFdYUboL3vHO
ssSjbG9ZTszCUT3UX0glT0RfChretYeY5WZMKEzQt0Ea9WJW+YTcje6nCKnaAVr/
muRx+kMD/q2OI9pKoqvWEhnf694B7JTKLUJJ4zGq4505kVJwion8EJbddlXyTVdg
brTAke5OFmJ5t8K+ZArVLxLx4CEZAL6SJ8uHkbpbtLV6IMZF5M/fYMJI30qk3sIj
wJ/Y+qcd3+3RNNf30NMyxS2ibqBaB3oFqnPfX0pSI0xk7JNJXxUEdj/yh6t4Q0Nd
uX+FPBPm+RT9QsgOXwQA4Zht6MQ8xI31PjhrG+MicwATxyNWfaMB3v2PJXmSuRoq
tJ93qv5izTIbAncacBS9jPHinKXjUXefVxvK0X1OyxrlT+NPfbNtplQXeY5EXzem
yDYSDD4Kf9Isk7jwS8MFUTlrhS8Z3AOs0c0eQ6eCvqwNwgJEawOAvujbAfchanO/
6mzjJ+ocVTeYClX+Zxz9REfENAYiQ7HbxeTPTQEPgSFhoTCHDbDpFxjrWAQ3VdEP
lwUhfN2mY1ND6Id9ez9qZcH61aCCuQuyfIJN81O8hUAJzi5B9FK9j4drzRS2ZQjU
MW6ocUgNvXM9ZdIdK78SGa5qV761805D+BLUCiCtvfAjEjdWYHIrxDsseMK2taV7
B3SG79i/kdiw0g6ujvBCDEjxwHh2xMYQENaApPABKRckzylIiPFatmYwALLBN3zb
0tukZt3OSlCdvXXBl3/4bGQocrb8INgQxBD1JAS9Rxdqc+SZ2CXeU8U/bqBgg1fA
1mitESAEwmx+635sAT9p4OXfdlVTY5/jdvwFMxBgmdBqFhiKvXFXuV/PFT7zXSfw
OSi0yOdYccOpxOpsvhA9upjQn1v0261A/Zuv3+dXo7IdtAdfLajPqh0MdCW/0OzA
AA9Duco6uFS9W+zmwDAIlTnuVaNAd6ZLaSetWxlO9gQuz/IM6ktQ1WcMOMqMXHK3
lt28XmgAZX36SyJGXPmhc7uNXKgZFWaE0ptdqYVYNPDNQhi1mNTbp36lQfJJr+vf
a7yuRD2HOiC2yG4sG3sRAchSGd/179fFYPD8+J4UVP0EEuk9RuleVr3ZMA3317vP
3wwN8d3O3ASDwfcsPxWG4VkcOzxqo3nt7jNUsvOb6YlDaQEfocnQFCt1toJQvQa9
W5uZCjoQZXbVXGjfixGRURPnEJGvreE6tuPYzBOJiLzbqaOvJO+drHiXr98GmS9p
PB+T+asiRw7ScTykzD/8iIyuW1rGG2ohBfKG6S+MOdhleB0RUEuRfYCrBJpa3Hi/
UHcfDISYFJbLeA96KkKq7WjDlO986XffP91xG89GG0a137TBTTr4+q2pGC56bIx5
6p13TQYDaEa84RvkP2jlhdZ8OmJ1wsvrEox7ftp1EcTgY3MswVNY5cYFMkoy9DEw
XTo2XJGa/qcl4ZTSxAwvnMZx8n//GATdPq4ZVyqHwMQX7U9N3QjEHs+DO1F3RHw5
FBriafHOyJ1FfUYDtgRmn9BNHmp/Jq6bjFs/MnmqEgRShzJ0y1ABJ9wJQZoO6bpE
uG20OYrNFh73DleDSHC0uTZwsy9kEtbTJQYF3QlUIvEj6qjdS9Z4uR1NZZHyHbPg
lvQFILplnGsDtc4t8uxvUP0Hzj8PJezLAnZgpcm38FkT40DcXnVmvRlnAVwvrLHy
iLQ6UuJLEfDNdQarTvzhRts4H1xDRsjAYbAJ9lT00NjOAS/vczSkUMs2p1Cfa9HG
Qy07rPsxHgbiLfSArnYmUX9iJCn/0MQxWcmfOYNRnvUmU7WhaZfcjrJ+cHjX6Xtg
sJgxridP2reMNDU4SZux/vBz3kFHPBpSfoDZ/eCyJQKAMuEEqnf0j6KJzm16X0gd
0GotQCwt+x6xcaHZ0jq+2CWifzlCp0K5FVxPtefcv+an7xDT/KEd+UBCvogqbisE
cIAmpnK/taWb1v+eW7oXsEkOykWvAkfpytN7lWng5xT9hYtJy9fcm1KbcnDk9XVB
9ptLqpt7rUtI57YUAoJPjXTtH3Tu3aDTfV+BTsHKGQfbq7SFvcIPY3b3FuwCyuiW
jGLAe0QJgkDEqjleG29X9G3Bgr0In97UBAOT+xsvXrrBXkkiC7lDGkWCu7XUHWBn
BHx2XzSa1zsuXN3jCIiSBw5xS3/w5fxcwK1XW0CYs7tg+1WmMNi7uhR9TlNeFpOt
UYzDLjUpc+oWfxKoqekMKqRVNb/aOdP/k4Fl0APXtWEPNsonS0WkKqbeVu+60yIf
6f963GY8n11HhIGg0KpDOyEluUd/bJy+k6wzKID/mPnpusZj6H+JtrbaqD9RLjHt
1TUDCeI/7FRPeFpeGby0Ih3TJHxU8DEKbM/MnCm7dZYMuiLlbaSTzqVQKvnlZ4BR
A5VtpaXEP0ESjfdK4jAE4Qbx32oLR8cVupBIo4KOZNGu5HoXLxolJJAm02DRv0QP
MTdEiVApEPba0OORVOQG70KOgGrEQXSKCmrUrCXbqg7Ccx3xBEoHH3a0CmskPO7i
0Hevte86IDuYRbv5qoHbPKhjOyCv8KtEfRENZsEhwE10rzAXlSJqk49Joh4nBUpF
4uxYSAuqhgoWL/n36JGUeyjbvY9lH3vF04ZqHY5Sn1LfRZiz0MJ618wxv7X+jtIp
p2DeVqgj1liMuK5AziKYI12vEB0yIuoDqPELzK7YQwp81zNTk5a5QKCP+t73VWq3
IN4/xoxNn5J+pW/8x29hj5/eQu3+iwzRLjZssmfk1sMb/949DM3obyj2b5V3vCZN
fokrePLfjX77SbrZqoMXHOlMYNsrh6/QqRe2s/muWVGkkT1Pa5txqhqFuSAvAdxw
5FCEAUajPkBO80wzluaiyDQc9IomrsVS4TrLQqZS7RO57qM1LWjvWGkEbmVMaJtp
FoyhqNtk4iUt3jLtMZpAhAccej7uctJnJMmLoGmQqQsUFJCzI6lTeBlQQG5AVFG/
pLqBnpQDuAqz7uj6DBrDbfwLZgTTyduA0UkQ5f+j5Mh0OSX+39mxESq4uEcoIXCb
twRiRdQ2g4SUIlmmNjrGR3SsankdOaQauw7OHWGIvQ22Gg7TOFXwtr9vTbXgiZqu
go3NHy+jNTZ0hHN/oQVucLf3KkUJWVNkqRUDBNEQXbJQf+LL12hyUajJfTxy4PxC
irlDs6nqQVFNNcBSXk9F6Q/DeNL2lL4lifoUtylIEY1Swp57RPQj+XppkCXiDyz7
Vj50DtzZf+zEi1sNiFiQgmsW5/6zZdQP6W1tqLffREqcbTiL+lpRK/8zLWSZKvFW
SczhIZSNCXMxjo4mLdM/c5y/hkoSBWfeZRWUcaK7/r8yHkQ/lTRO0lRCgN9MWYRc
xh9ZgZuRFMlJuZDOe9MzOkkwUFlmnaugmHmcpX+6D+HdCND13plcHXNO5nfUwvLL
x8zN+jj0bY5zeOaYD1zN6GfN/Jfyq2EnwH8e2zCMXhHrZT0Vy+QnKnhdARgVJR0e
bzEo2SqvFZz8wb1S1WLR3Fp1SnnLtVEy55bhKLePLIlvRUvtdoS5sCITeBjppIXZ
xMyJnJvWT3MRdTBAqp7kSEV/OLUguF7deXJYNviMkoMBJ/AcLNZOnqBYUSp+zFWO
bWqEFpXZ35GRPePnaChTGSpYgbxiDn7Vt6W4Sr76RAsdUmjYHU26Dnd86lm1uwWu
mww4ieB72QXcTr2D27iZXuuEkBFCFr6ImZJgOCKyKrliC4sr5xAaEel2iVKWbJdR
u+Af4edfDaoFciYmDoD97SeaH+qPTJadCnu179Ao/kSKPkec+EjTvLIvzEESkOha
mz4p0dBRazv4I7thwbEv+p1pHy4H9ZtaNuyUakaHGpAoUpKrGPdj6uNwTRwzmiKs
jgxUEU5i7yw7L6aOazAdUG66L3vJUyAwWjPY5WNurZbZz/WIlIcsAAtryQysKO64
szeylOZYMsu7UdER/2hpv4g2xr0nYSCN8qCt2Lz254FzK7tPJCYJqoIQ3ff0LLXU
CjEDmDmIzTBg571Og8hcH8V+qSAdpBKPYHFhcKo2/ih6YInFFL7uVZ704pqBjPsb
KKrRvMu+x8oeYz9uTDR84C3tYUbETaBtzvXwXC8KP6X6vhLyEoXx0ipsFhc3tD5O
fVklXVmBlRN3BumpO9jRZymhb94RK0xEgDFPn5sZYEkBK2swFp41MazGtdN8OdS3
m2KNv1L0rbqPycJRknxADx46DdyvEFWSiHPWH64iNdCBuFsrG4lPRThREXFEVtn5
fZ79rRS8wFI/SfhlQIxEyNigRNEvcDMh9GbYx31JU7Nufqoef3n+HvM3FvS39o49
5ryXKs7GFcepM9907ztCPdSVeYc+bUnzEDqhDoK4ig10sUYoguAqTitsoKf4LamQ
zGlPhmo69gQli9Luy17JNeyblqhE+Nn6YI8ZUlEpHgxvIMoyDlmDrFEnMU0A1kbO
0N6VwVnzJI02mN9Hc4eTh9u6ZwNiTZVp8QY76GBNNk/biA00mVcWkNYI8XIyjiut
MH0+Ua0zs98bpnoEO0gIzM2d3/dRFwLjfLeq/eq6DY69jvBwfhxxr2Cpp90RdZ5P
eHAErBUy7KZFMNY6gYK4rMgSuKMaiNI2BeQ0OyG8ZYG9QnEgiE7l4MMGZLORwf0h
+LyTl4kU0lYMNFrTXPHUxABzRMr4I49Dpaji7be0nEQHoG55ASYo8BHzyHEqrLcR
aVIpshfY4PAbBFOlY5dH2B8i9zwTeGJesckObzNcKDkJcd42azBmrT64f4ZnY7bC
yUY4LNHKedjumXe2cKQDxXRnYBzGDosNsVEXeFk/9T63K4/vnThzlEiOxZvx6Ll6
5cXnzWN5i2uPRYbpvtPe/jLZLWOyzYBhNYJboR7Z1Yjq9sh6Yg1bnEjjLrhxDCOR
FWZADyC7lTfOkufpoCeCkOgASqDjmZf0FJMKg35DfwfSI1m6aykCku0o7MXc04Mg
SMyu0kOTQ+lRf27z3I3u6iWVyQqkjpWqhb3nGkD57HAuMm6rCKIr0eLasoMQ6tw7
efrdIn4lpenPoPeW05CqsXcvh/Yn/5sQ7Z33ogCxlAZJDS8bXNB/tHpoo8lhB37b
CFQx7cDJ+/g8q9JyAVqv2VSJZufw5lmlRnV3Gm6Fn0PyflTmjVUz0lUsoCnKmTqw
YnIuubpHIgHXvy/9+eOVN5pGoYlJuKuuocyp6ZEudpp/Hr/G8BPVXmiSNfhcEVH+
ElqPKcw0csYM3O+fjIawO3Ae5UnAoUsQt7c5pKDyxliXkue5XHVEUGXrCtcQv7vE
om/knpw0wYvW3Dwvdr3D5DdkFwUfexP9C30RdNQQ5BQ6O0Rf9QzkfqC/tkcedjQG
MR3ShNLb9RiZPeLsC+qZ97mDCRoAR6P/9l2BjSyw8mhqZGylI+cNVrymrTeiWfU4
ck+QO48NBW4VPynChIeRc4NKPoyLCHliKIoqXd0Hheco25NlCjw4JciL/vvRZ4hA
7XsdwPSxiSnjtn1eBxY6s2mlyQSQhwJePBu2Ot8Cj20G3JJ2YlBVuzrufnGFyFvc
BO5TrMhOcoZP7ruwwz3DqBqp87qC5Lju/wFZFDC56fy6xf84EH0qG3gldp/CwP3B
4xE3+OTiI7eFm45XRYI6ldqlah3hl1/i80x0uV2zFqMyy05kuJtHYZUIrm4fTZur
dPryh1kKSE1O+jCWJ78cY8odYNj1qOwv922Y8CmiKxCisdeNqc2LJcv+Do1hK7/9
wQCREWJOA70ncxi7htP783KMTs6YUMtxcKI+CSkBhhi1wT1MW3RgGcGBD4ieWeMc
KHdbi8KFmaFR5QRv4vtxFKsGQBs0je9esS5OBZjNShCFIHHH/DlYiUdYXms7LU6Q
xFrFFG5BfQdA+EwE8TTpy9Gj5D2JCOYXrlWB40uG8oiH6xGI3LHZN66JKGoWkNng
BHWUjYDkJjmpwI6e58Hmj1PFcKn8PAMYw/hS8W4ZyCYY+SwQF16S9xspswjjAWSz
jpxtN6hClbeSuisc+tKA7NOOd3CqSK9uwyAZuvMkLuY5XY0u2wfA/vXEvKssfiFB
Q6k86Hw3DB+Qc9xOdBpTAbotGoOpalGAOtrbKC10N/Qwr7JXdPjqgTE4DXQd0QjN
Ajhvx6yyjByZ2JDHHKRHO9XBJHuAr75Uty7tS8App0kwhbhdf3erH9fG0ZBbM82D
V9etd7kKvjZH1CJCUvA3qFNrHzvPINgJBUUSnvZr6BKDLa8yKX3USeQ+m8VjvbNf
i6+LOAVtoKohMAQrYw6AM44p+r6mOFgEalF8D6W8UHh+LEj7mz5epXPWcEYtOmE9
hBvHZe6I6EHiuC/0qXXcrGGPb7AQfCiUF/cHsWwNvE3+Lw+dy+TH6qhrmPM7SOtV
Gw1igh3EI6PWX4lRkjfx05XuUQeiS66NthkrjAMtQIId2q5u8ix9fx/49Z7mHUY6
lOlC/ZRKd6WsieVkCntTeqHTxttz9vANtcCBQoRRqWIIzu69/Ci0T78zb/RivpNa
yenwxBMDnvDJxE4FY+Sx3jBQALDrcmRhuQ74iEi13yfHML5DBxnhPKzwO4+KqnH2
Vx/lYXw3Voaumd85e8xvvDLeAbUafTFX758MVqhZCbRu8jjv06tQ/VSuHDdyNPmQ
NUnwRzmhQXc9QMAhBmvB96xB7/sUYO32EAblI8x9LpeY+ErgkSx25gaUR8O8UYDJ
C0VEkngE792gFp+TXVNgkBcqbpW4Q209y4Ha6cQxkEz3NHArddzw2oVt/5Sj5umb
VV1+dabgAHYmluv+k5cLiORlAH6dKs7Lbkp4OGvjlVeU2DXjPIqH1otwQQbOxEEe
hi6wW/TcBs0MHA3vV8oeTTPy8nI91VOdSSIzzG2SaqefgM2XAJPAF3u2uY797kFD
8oy1lpGkJ6YXkrhZH2FbsUhYo8ev0bR8PahZG7XI/BEWOFA4SEOU5WtdfcCxOhx1
Is1YF5W/4b8dOCy1c7C5patsn7q+ql84jepeZcNescb1+hmq1MKrGv3eVx8CSfCp
D5GkbhQDqkvSo8aVpR5MHrdLD05uDhweAuLJXBNTuRtT+ZiN5V/Ene9hjTRlqiMK
IL0+yr8xYOB15l7++q/28QHf/+KHWfN2GcHSOadLxv9GlUQJPapkJid/dz3C3a4k
2oImLqMRMWBE1CiFAMHQ4UXW+tJUdq9RYMwxgvteZ6Dod+V7bn4B6v++OKWlLsvA
0nBaZuiysVrdk0fzO6cPXkz+8kx+getPsxNB66jopg4RF7MwfLhmF70QGCS4OboA
b1h5gwsqPry5BbwjwBSsG0pgbtCPjDUkIy7+so5Vf3Evb/CEkJSRJYkRn//YhCoJ
0useO6zoB79lGb43F481U90bGZGeiuDEfvztNhucecX0llGfic+4+5EAFzNYxTR4
GHxsJLtvDLTMkNkPlwdHpTO4usO0RCyzDhUjbj3V5gDsy70QCrmmC5pdP69OZwse
VTh1bjUaUjlu55qfgGflhjPOqjfg12kW5AA7iJix9y1uGXy19gAWz2eLTvGgyG55
UXb8TY//MRWe9+LLbFwlUrAnBUZKZOT6RuQrW/EjHt4DjiHq4FzIN+9bUX88hQL9
/pBbNddjTrlPxRp/3pkjer08pnMoJXWmYFFc2y1w3rLJwBAnlgbw+PwbRftZwmEq
Bo9beDcCUTo/80aOgGqucahDeSU+Tv/XxsFE0NdLGA/PUeOn7ixsDooKF82CL8TG
91d6k5cHB5GuwCSINmet00DVxI87bhADqZGvOzTyDAXDoVbI9IvXstN7rR5UR6HM
VvbvYu+EElZwEiza4O+VRIyjMDMAICB0nVYqxVAVeygATCRiQnr97WGxY2UcRbTY
edSg9CZOfaa9lXuA3GKEZDsv5aBzw4uHP82x6AEG3tj0rPvjToZdwMEqrhnVDF2G
yKoXFvyauzIBJvj92iCPws4zUrsLgq1hxRrdjKbIUqm3TDuZQ6HJkLDWMhFm59Xc
p3Q/vrmV3VVwpDqfp7QbKME3SP5eqw9NY2cEhSk6axi2tmwXaInqBGKpexllQee7
mwSSud7gkEJigTxYYcnFzcBrQZTk9Y/IX0GtoY4uxfZjUEiQRZguHVq9tTv8eU9j
/rPq1pjxI+LdSbak4LxTnnmcYvFb6dCSTzBEwoAj6ofMAbUfJfOBS21ml/lrZD5C
UTtYEuCn4dxK6LPQsH5ZZUqrhKR+wpJyCMo+IIwEwSXN7xS1rrvcBZAGlUhvKs1v
uSyeMKcDnKEM8rGXxIapRmaS4UAdA/UZVffNN/ddX459K4BJLh8JFmx8oRkmhRqe
F0ujGKvQsSIlZL5Xug4RWC7c+o6OUQ6YYApHB3I3DOUlyJGRhoUska8IKiSlqkq5
Q5YdzxYg+p87bpIiKXci06UYRWJjNX6D9DphS7H4abp3tbOGsQFcLAvtqGyR4gp8
P2myMqJv0QrI0RxkNkflvhP7SYbwFfU4XkoAEezOBUBx6YzDEYH3bjucZpdBZcdw
j9mjbL665U14S7esLMflEUd+IlhASZChK8mgRIZ9w9rXhuRsaU2hHyTY+Onavptr
xm388hdQc5en9vC1QIP1ujEmXLrhfSapeINsD5fx6TwFEmUXGsq7pAEioqiW63o3
z1SKG//YbxdWdI6c790k7KwHLS6b9sNWv1nl1zd7B6HhsRvzaaoYTjvYlIRUBsBl
jSoWxxcDItxpw1nVuY736M+P2k93v5RHaZCTWsZhNODa5j1VPF+Yjksus/5c7c/1
X9HIs70yRxkQD48lu8oxWQgk6RYvE/f60zD6WBvo91QJJHblecKQ7XYgfJzjg+R8
oJsblMhMD7ejj3xoRt/fAaZhRS9ixmSQeiu8raPGxXzNCbuc/mtM7zEi30EZRd5B
qwZrcBTMO6vp3+tlD0EbJbQpCMe37DBASV+csZl7gay+OtQFs0pjPeDu4VneWMl4
PYlSoFTROWZvDvpUstjmG65lhAEMWMzD2C6n0Ry/TtFFwz52hbE/+ge1YJd6Jx7/
Fy3Jr+FkjUWY4XqyKnHzOALj62NzMURE7kpKAYNIRz59tK6w7mp6+L/J3IWFrEhz
d3FrMvT8ArDNjQE8/UpO0ALCUJXHsCQ27Ppg3lLviXvnLjwG+2Zscz+JRw6yByY7
sh9MPcamRbOPFbIS2xhagus4h8RULpbEanBK07vjNRgJC9SDeUk0BR7fVo5C6g+7
3QT7TQoA0qdyl0pGQ7tCdIJEk7sE3c80CPbdbv4u7BdPyXpOejDRia19qWl7lgVW
ImyyM/vgfHFcYjRVGvolxZpYuHwXDA7penOIyhg/79wDdnTUuNdrqRVnz094sO7X
Un8W1NJqdQjg1QTgIB7VWoW7ZiFjHr/FozZ1f66zTHE5xuA4lpgkLKUTzuVI9O+L
1zBFsadqjq/vuBi8QdZ9h+gDrsCPdGl/2yAnT4AXgE8Nwqj2f8rO7dQ03S5pheML
uAtzPe08SJy4JXRslfgmjs7rNH2RTyv4c4PHnAYikeuCjBR3/25yLvxuEvwTcBZh
w3i6BQz5nhK1TBS7liSXUGoqowNhgYE61tRH69i0N0zn6GZS5x86mx6wealjzAmp
rQCEoe3ZbObf5xOeNW2bZMTd77Sb6DAEilyOoKkMpJdr2G/pzvETQcYh9OfbnUwM
IKQ+vG+CjWLg1gk0u4LlzSIAzL5QUrc0ZRcVR6wAqH2zACu49iYw6/D6TgEyisQj
Ca5+3EhN8vfqGrovfHxt0gdb2HJ7apoWI+M00N73Nsxx2ogiZvyMxB07fldaHCI6
jgcopIPQNxVZUA/QgqLIa2PHojmHxr2BX050cQN9P0Hbw7f/rMRZNMRJjOahCcBX
7+ZRCBDZ1Hdps+7BJ++rxo6vhnUxgUrzLqzwQY0Cg83/O/dQSo2lzuV2IYXnAjNL
sU73Oe7avoS0F9Dal9RwXFXT5x3/RJxABrJX1rvsId1ShisLwWHK44lJM8wt3P2S
vekeBiS8EWcCpH/lFd06c9N4S1g9TPGzSrEd4GDM9U7h30kYhkBO9UBaJ0t1cSQp
p4tDyQEAQdw0DpGd8qITXKzLzjOVJZamzpREk7J/yGQWAR+aG2bRKWo1kuD8WwoH
ZbFtPNbitMVKGJqHjrvLFPxlkUgTwX50IKrnIIaPCe9ubHR36ql46I4jryEWf6D0
AAqVLok+dl/YjTxwvi5Kib47AumS1cJUHTSb7CwxY1XDbYDLYO5gH3LE09eHw9uL
8xOS95DtczbY4jn7O9cPwuRAkPSV6u2Kd4p1DpX8OfVnJyUPYUmI2EI5vBkM7z1t
m7etT+MIp7zGsqlixydVdIzpNZ8dp0J5O7jqWdr8DukW3viYGm7UmFJjdb+lAkYx
oIA6bTztUhZBTeLEGe+AaSMI5rC33eqGahV/WPGdW2g+UJJBsbDNnpaDWsXWE00F
KvQWb7miR2lZiC6UxNLbewGMdEV7lryleyUA1k5duy/8bjaeMHUyZnSqmY1d5Mwd
oHUF5rqAf/ZDLOMV1faJwLM0Y9xeaC698UtrQ9BDv1w+9N4nOP8ADr7dCDcEssGK
RG5YjnPTkdB5tAxIMhECJweXW+tE/uGcP8E/ehAXvLNgZQlMAqSODqbNRRgWEid+
5rVIkWoz/wywNNkvc0vN2ciaCpoM1VhO+mqC/35o/myGn9OsA/ijagCzj1aiOJWd
KFTitaFy5RhCbUsygGap+DL5TmochNvvukc2Hv3JeiM5fcW36DjAcv4B+q4QXR6W
humUKgPCEHVIX1xaI9Sda4fE7U7vngPZ+HJkXW7FS1ouh2uNSEZ5FI1S0BDmTMZr
tYECUorzuHNtElbIJ6yqh9LMGmivseUaz/Kb4a4kHYC8kLSosIhs2xcnZr1iwJ89
VlY+G0P+1qItIwBDvFFg+nZ+iO25F6Vd0zvRJlEl67HQYAHDU4g3vIKQomFbi91U
9exBNuvWXrsg0kCUhM4rXOl2h4yhlllYv+zNeF85hgBw8AqFRJ/AuX+7X9F4R71F
td+C/wxHbpo7I2sf+3+B2b3Y+KqiQTRpaFtaz3D7wyQU07YmbnjabYm4ZNLyH1R/
NEKY0IvexI+77PtggCxAFIQ/Erf6CjGjZHPvZZBalGlzyN/YxKJQJ0kmmDWLTHjm
fnnduWILQ6C8BaACAkRQVs8lw76brXonnDWEsbEoQ0Goxpdrb2DFZvbzP/MTKq9F
s/kQ+JN2vkD34iisTFLlFkEbb37uXN01Nzp16Icis21Rl0dRzAuZ8VgLySp3OI/S
1mDqKVP9dlvIivziOHg48mRXdnfXDneoR/1HZ83n26CkoKGxC5hxKCVm5Lv7m8uL
KWQ8UlBzuBau/gZdsmJJCUuk13ioKGgfgN0/kES0MYoF0BFESDPvcUurxG1MHpiT
x2+urIXFzIi7qvbVmB5XSX1G+YFqXvpBl3nU2CYgK9i5ctCf5Drjphw/oBpJTS+O
Vd4Xe+1fF0MBma1D2wC/jMngIQTygxB2LDFoocwoaeffiH9jGlFEh/YWOKjc+JFG
yyD6PVVKN1o/6Da7JPwKpufHulg6qqCBKCpfUAZ69iDz+ohusDhGio5Yj4xkyqGe
/tYQDNy5L3didF+M3Ctot00tjLfggqTsPUFZR8bp9qAb8d6GSXCb+9B2kksXigbM
bebl8i5l75JbA92U5qHgADyH/686VuMdVXtSya/x7A/CfLOZwqW8NTGEOFsBc2HF
tHXXRzzSxHbRblnaHPo4BeblJpsSMVSfxnxvTCe0lPB59mr7llPSnsIaii1u1WFS
P6/21aq+0hoQb4xpyOxVXL+Z7WwDErGnFNaoXIW5AomJK6itY+n0CMFLVS2xwdam
7/5zsAp7AAxAztK5QkR2j2JhU8PgMwaIKO1p69DXyrRZiO0bpRxITwPHWw0/Ne3k
YYkLZcGJgavTchRS7hX17EO6uEpOwUipUzWNl0E198+eWytEcUm6wMpvB/HSvP+2
j9caabp7ZmfJ6V4zj1ZlWb3Uw7KMi0UpkvQOqd6m1IQH9xIA3wy39EpeDWkJ+cR6
HfaPM2ERfY6PulnGnOmQSrebhEsifks4JVEW9zTflpSFF5/Gqf2J31MOBCazHTiW
xesrv2V7jhV8w2CtDCSJuAfeg3JnpOY/DcEVgdHnhSguAQaFVQO/Mt0wcoEY6+5S
kMjp+NTwr2x9MQ8XnUwI/865NT5iFJlDc/Z2PE7/UBpvUjRo0Ix1B+/OgVMzBEOM
YoF7n1QISkslpOQmwdJboqada0lOCvlfThzojsF6RQD6d3fB0B41HZPpiLY/mM2x
HhyI5YEm1QXTrKe8n3tDfywsezLhGbpXnu9l2BPUP+iQWwlsmMbI8hPelxew2SuT
f9eh/rCpPPe4Nhi81XzRoD2vrYbiDssrYu2rppNuw06UzGF7BJTml6hbB+ffbcSx
3ByVOidY8UWdAbvgZab4qq3yF3G2ijxcv8kCsjX6PK/Cv13a/ys/GVe3fKNUg4OF
bzmGpyfgERsU0MXQHZTOikpueFrBIq2NRpQflQglOvX/TYl+42WSVoMnvOVjBK0K
Ut3wQOpHIuIFdPtF8V875WCORAcZHAl6pVURr0jVjqtHshHocgbmaLkUy73gR33D
pmLxbWLOWkkwhEcH8s8A16MuH8CVJE0rfM6UMDOwlz+SikPkiR1Qfvr4yA9lO4ZJ
fk329eqHOtZlR+/BReDrh93A+I6ld8AF+IHo7GOXnvGJu69wdnu3Gx/plJThvfGO
e1l/cPBhY5Flk8tXWgg8ATyeqZym2dV1OUmulvLmXokDyU0YJxuKcyo+IacDhe/X
qM0cd0nQcln8jRYeQCOl7SOKpkmh3BMbDrj0VFiJRR0++idVLkuyL2chAxcVV7Bv
sjgqIMJnOxVobZ/lUZeWG+d+qnKQ4xOyUF7ExN3Ev+pQcJU4O0eIeAA3DT/Mh4ls
nzDWNcJ27nRMqCnTzzaBsujCpjD8PAHo837HUDizrY0lfnbkFk1MStbwa4YnVbeg
CdFbIxuYRPBa0QjDlxR+ipEjR8u2xsoH3KiKMd82vpBM8wSD6MxaFQg8QaU53RuG
mCe3O+V1Jgpga/HLuIVYc6EmvpxOJUeDntIYEs8iDiOs4P9i68Nj6iRcqjIPATje
Y+XAUJXSzwQ7UECJFlxa3N69A6XIThYOM/P6Po1+dW9nU69u453yvG4CVLq0+kDm
b8eAwEf5b9HT15kSJw16kmv0/cJL9fenxCpqvgvvN6fUuPRqC3ORMsjvlI+ko/ew
E5R3atUSkiZ0esegAEkMjniLCVEphT0Lpi3fMW5x9TkFp/vkCYr6JHGOGPWRYZm0
pDigzZ2pWiHaJZ/fMPpT9tTX4TxkMMEz4JyJPj6BLcgUdMeyl6kANvGPjgBqk8Uk
sR+xZiMbzpDMI2Oa0Sc9dflTUTDk+TTgXF24cOGw8BKq2VS4kQwX9lVTfYE0xK6M
IDFi47P7CkZ/C5KYB3e/lXxXmFrTN8BgWDw3XL4e82cDjou7gJcmesehTDIgbyzV
EOQ+AmWtC2SF0WV5fOq1MpxPnUh1Uer+S/V+UD0nxFm0AAAfWsXFdeV+TsnAMBmF
6wD0gfkNIz7YLBhcCQ0jyqjXAbdnpym6TySFa/5AxJWu3IJCrLF1hTyRrDriqIU/
KMqrJQ4rBA6aaYAKZmcoNAa4gCwtujqWpF5pA0JqSBTR0q5sMs6avpG6aVsOU2lN
20yyn0DM325gQAaTbEa7yd7hRf3X/6NfWHASsMHB6l5FtYt2Fsh8Xc5TXZXiyuWJ
NsFaa/+PcLO34oULTuO6jU+WXiKmBCb+YOn+xSZR5eULTyLueFe4yWu7yRZzVR/A
V3g/EA8YccKT0D4dYP+4sVg3OQQxPYiPMZy4yapTM9xYSUZc3G7IZ3dK4+j0F3vJ
6F7r+GEMDBepfduLWxUL0aUEAd8gnScJM5g1KwXEqwH8y7imFtCo0kL+C4fzOXsR
DGnl2vKhiDviOaupAk1BwMu6ghG+6Vv1uxbmT0T65GZblSJh9FHUwwXm4l+nprvu
Ex1iUrtLxl0rwsyQ54WQ1PNLsoV6oXetY+U/Json0UZ2cTwV/bpcoaii/8iQFsQN
+H/KzlNlmXYCYM0UxSdHgQfUsjx7cGyE7Ajwk/pg6luuRs4EX0pDwgTORgqMoOVo
pC9MmgPXIuyqNUUqpRXJx/RwgDrPlI/HBkLlJt+cnF6fChd0Lk23BGcEyDNVw51u
k6RYm6zno0vR9UE3Vl7ac7bqMN4s3ZXTvu7so02R/nsglwSmbia5aQhZj4vbGTVe
hBzPhmvZ1KRc3TTPNRPldpRzl2vVK+m71V2tiG60dU3ibQOnL3Lq+jw8T14QXciG
xdgzhtPA/67mAVYe2f4dXA2LpBiYGmc99NaDg7yUbL+tRkF25Kbv7D4+bMX+ndLC
g52f8rCQTJHSZA3KbnAZOqTtGCm4hMLKS9Th9Cxj7TDTo9Ue6VsFQ1NGARjkBRiC
0/GsSeBZhKl0rGlqBgWNyFomax9VXl05MnZ+icPcDAvixVrZQziMRvICo5KJv2Ki
oVDjZEj2viKxsbGeY9Ng0QneYURdGZLMELZem0/tytNz+rXLy7DijMuZxaKOLJvM
vm61drMNOvv34EWqwAf/t4o80RV/qt3KrOgyOI+seJJWgcbNACkT9oHC3vzTdvc1
VW32tRqDFtupfgYlIEbniznu66Sz6nePTtpE99oOyCojIVNph8t3fPNLwaqO3mc7
utOYzbyBU3f1IBfO8KXHVBA++BMnUuv/toYRvWFFRtb/zjSqBfjrv6fKUxF+bffL
VNjfZsojzIN0ddVz+I+3aLjtQkbVu26BcwWFsnSL1PIyJP8ahoXY73hDW1roMNq4
HGo+BDryOUCWdxayO5tejV0XLgIPsc/CQeVzNkGpBXFYB3xldIX4Qxco/y1L/4hC
ARF7H519eeaZh7XQClHiDnQR1Tp5G+7GSLFeuX38Q1/t2uDgg/ZYKXXBUJ5Bl4d4
x+iHkcqLwKPZpgoCnTGr5wRK5z/tQfj/OSbzUIPA6VfrGitB3EOvxXSlyrXjqRWG
nwsbDC4B04bfZJHHuOqD/GUc+etQBUyHG/fZvE9kEAZ6mirTmqeiEWxYV8ATzUJX
ktAku2fpxhoyqsP9M7P9/1Qu1y6z5ZxXomYXIWekyVt86d1WhgjH8CQuPjxOHPAA
evBw1rSnUmamyVKRmFIXeQFwzLNalG0iYTHn3XA52xksDyZpCetEY25wHXQAqM5I
ochzShwjjd+H1HOgiY1m5I0YPqOy4en9qzSYYVKWuY/jrLP9XKNY7diI9ZVmTcPF
EeD8PkgOyizRsnkHCTdigyk9HkPrbppGxFAHzSsd7ylKHHKL66fE8Ne1xilNgerp
GkFZ6auGmnU4YFHWyRPOBPlT3aUiiGOS6V1mL9Qrko3fxqoqlgyV6OUDKAaQ28Wb
bwBiScDLZXNomYD+qAxOK+txnWip/okfg7Bv3YUqFTE0TFM80iR7pAM8cKnPC0X6
XCFLYo2lRIoeNUZGpDr6PmIfedRfzMz6CBDd6Fq9a3QrQdER11xBRtll9aY7rZhW
fpPaNGNEPE6Jp8dXut4A2RnkIf1tHMWiMBGOSf7RTvqfE+b1ED8M9mGmzQi+Kyv6
eY9shOKXj5CroQsBvODFcK/Ef1JEmHoc8a85lyknzymKKn5rNBokw+FglMR+plTV
A5wyiYboKq4z4/iVGzWYTKbLs+kg8nuLSIWmy+MOVCtmRTE2RnOahVR12k80Bu0/
Qfyg9hEKzUa9IhznIhjfIVOqRTvw5NJSrMyglxynoecV94WPp0ZXGpdlxkf9R/JO
pdZZzr3clQYhYN2QzD7Obk+/uVvQkNQmN4O8i7UiqSSQho+9lEhsFaxJsrHh3g/Y
qrkirfH3mrCWE2eAWqBW6dpOx+uMzIpiQKK86BJo+xNaNY8Qr8+5eoBkpWzYYZBI
1EiTAfRZFGLB5VUGztUUScD9/RkHaz/N9qcCaFWe1907u32HXitMlCBp5XzV+JD0
tSij5My7OAe/w7F5vSfk5CZgqSBGEHoftJFtLJFgP9OC/JW9dCWIjbPQDqocDJjR
sQsZz26+tJhJkckY16i0e5dVEPS/7S/NmoKWFo6LkRq0H5VTxW89MCMV3vUI/b2O
OieR2Nq4oqrd2yTnoYjifvh142oDrXdsEhwuyQh5cceYnKO7ExGTGg7+K9KvPQgd
qMRCmbFcuxJsyni92nPL1KA+E+5FH8Xl3zKwPA6CzLBOiCAryfAZtO415c+nBXPd
TiSruiUHe/wA1HZdSfKeyCYXZ5snOL76FOEZEWIf5LvGxMmM+kmSCwWz+oh8B3CB
CDDUxGw4tYFHV5E2AgKdPc2N8Uixhr6ngSbgil85OqiKn0sJetOjkPoh0nrRnV3U
aE5MSuyrHGEr0PLTzNo0a05gh7PJj+lQqL2lVPMjjMeSmDZ14QmjkInpLT0etblh
5VsMTSEjkPN+/m4zINtrssOYyHweM9/eCSzGoVUcYG9d1+pZpd0X3ZvjrnvPf+t0
JuN2fagS+f9majqfX3qPprLoofaR7n9jgCgnJVoYcTTlUX+ZOdYsk0HhDSU043Gn
SrU2fSn3QEq/KFJo2dOLb2FIvdF2p1V9yypsIEAj6KDRZN+cmEG9h8jiBGMorofi
naViegP7k1Pxyq1HOyuIn/1HtIcwkYJk/J/ZYB1FQ/rYvY+uSXAJPWqSvaW1Yqem
RIX4nTBa0VXEbazctVgaDdPeq6Wa3gC9p2R0mXOMFJuJlH3UgANUZlWXHyKxIbJd
3OZKZAvdOUGqsNc2OJPBK2KmZA+/eSXeFwp+QDbLCZa89OTkKlP12xVUH2oWY+Aj
OPcvrBRa428lDObrNlZss4+TISfLHAsagVj2dspHnKyXZ4v0LepemtfbQAualxrt
goizGQRMLOrbIIL9x6OwsG4ApJddG4ner6USIO34e1b220sSzrucyyrvnfGM6Uyc
JYF/TGK+3o65wTA7hDQll3Urz4JO3/A/rtkf3zra/Y8/k1gECyCfwCXBgIgmLSr4
WS0DLrMIQBJISYjwm3RGl867UVnfxOG2u5rOhPovhAcx6u3Xi6vwp/Vv4NJx2yl/
iAsIquCIGtEEFsmbHTB4C9KrWEOq7xEXEiSo/SBFJBOE+TrgDOKoCZEGVmdRFSVn
xKQjk5P7IyZMZleh9/xAepYJJz7HJdiI63QFUpR8ekA6+JV4hLywcoTJ0yLcr/dX
W2Jxptf+a67G190CqZIRxWe66pCwt/w3KgSVdyvqg/5Qxs/y4c7VUypF8/O1qLi7
cehtnxxknM4b2pTLXpBPFFo8mddHbdi9WzCQDv54kF9Om277ep02q/MthvKahQk2
KUDUO1VrQUwvQ1aoUhjXKWVpfJnXN751R15I3rzFEQ6blzomaoCGcTqYs97lVa3S
7sfP4Xl9Zb+dEqbEV/4aRLIstdpPNOf12tUHeR4RPspfw6RWXifsJqovy985E9Y+
F8hAKyAM10f0FZJGYroYBSAQ/rkeixAgGiK073vxn2fadxV7OCJqLLIRC4KubazP
iKgP4NZvloD10vxp//uKb1p5VWhhp8hWkdZBCv3BSr0bMk6HDV4o7XthJY7utmh2
mKfL1u8LupAZTohBmtAu2Nfcvx3FjjJYU2gGGSx15YLu8F+a1CvIqUFomk6Ck057
JpfTWwN+ycyAvQAKe3fZ9qqMGUfyskaMHkJydYRo0D5a+LteSNOQeQWT+I8TLSy5
C6jJ51/OoInWoZSFodfYx5sA7V5sVUUssLPojuHIq+NuTUSjnnb8KkHxEH091+OB
RYeA/ZkWl0ywSSZgK8gX1gXaht8ZyRhdYd18RFC0r3CqgoE4YDOXO/tFxQg1OTt4
Lbk4zizEHkTNoiQ6jVD7elTYG7qptp3sCKLZsOOcf9zCCqArVAzcVL9OOBZZhZ4V
35jbGCakcHw986RTuGQZ09bML9Dq8/eo0y31myhnNe6iq7t9myEfS7eteouOvurH
FTL42+qRo7+H5Obm7SKu+mUCFmwyZyohsTE8nIpYGuupQ9Wf3weWWNaRUyfj8hm0
q0KLItdj/DcoMg+QcBd2U1La5QIgwjbGlDIOaUug55yWi7dUVfxHvkb2aPh6qDgA
tPk+l2oSVOuulGdVkDzrtboFjFZD//SQqRCZqCut3b8166wWA9cSN21STO6gqVJx
CCWdIOKbXKS0J7gkwPfHfeJ0k2OOlH7iclm26RGOwrIdLS+p+RgmkXMIxT1DsLJQ
MgOoGN4BxSpYyxNTPKhkRWvsltSHhkNJb7MBH4MKUmwbx547Zmk+DCEG/yFPH+Gn
4rDnFBK5T0y6dEVvQTqVdU64MHjT9Ay6FIKWfkg9pWFKXJf5Qhc4fDSUXlj826Nm
CsNuaebml1S3eFlY6MraBqdGmE265dGi7NDAapXryP9vTtihZONj8YU9N61E3+gO
o6jJub5Il7s/5bIXKJxzAPCGELwAvPWDd9A8nNI4erWW/tYBRxLREuMIvb+YGkO6
IakDwN/XVzXjXc/v8Y/A/kgVCfq26/1S10PqG12ydpmcDOT0VhG8Dh8MuvOL6y9g
wOjjXoaJpmxgwaI6w/YgID5FU7aZaVjotS04Ds4qg7Pm3bD9SYlzf5r4Sk2lGhae
Sdx+JSYpcfIMsqCbXckMHKhZTZov0o1BSxq0zg36k45claEtg1fTPVIyG2TRZqwT
3jtirAm1Wp8aiJ3EgMCMLggRT4mhoo2XYC8673cz3xkQNZjVZiq8riUxKKNgoYdG
+2pO7RcEbkM4+I5328TSeWVzR4Kx34B0Nw+gwJPsYxaJND782+dxrZ3gEZI0nuyb
yDv9oa2O9Lp10Y2S9499QAeyo5j368/CxsNXCOua9Xw6cQ/W1I3iNIrQ+0QJTod4
IhgSzf5b5oX9VYQ2MgJdzBwwBAS5zmtUsiKg8jK9TK2GQ9C41Fw1QPfwrgkoIwrh
rvUnf1aJ43Bx4H5O1agYk6Bw14nkAvkchSMOBG7lxM02Q178qIn3a/QGmlqTSFVb
fZwO49jKwr0w/YyMlEnMooZ/IshMOGvZvrQg+4fvelM+8ncfnwjFyLieXkn2Wqdp
jJJkqYslNesxTPaoFP92LW9PITIZIS83q0Z7vumrWHatBXfHzE5+6NPWf36BIkAF
PGMNJZyoSh3pxvgRMTjn+IVUWk043CpB5kGu+MqvkiQxZ0c4J8515jXpSfsG2nY8
nFJmyd5Q4Orp0CKbHRUwQ0EcmqEWcA7SILP8Ay6erKWLLQtqwwLNVhOswW3O0xiS
jCoqOa/4BKzaHjtu9OpHsLfDnCKtDcOVWwFKUKEfTINk1g/DwW2INDoNLZwppAW1
BiUzHBM0OgxWuM+siTv+M1OkJZy5nyBlhbpwUBIBnwYH6vbHHpg+GC13CQS3/9CX
9ozQfctRFAi/Id6L0CjF2HauYuMUWlMT5PyEDvvEZQqNKD/bcOmoi1yPs5YE6EB+
qpMknKkyrB24UTbbcftmyLQRPepB9GMWWS0kBnue5N8+AT5ydl9db23Uss7wpnJn
AcgJkovlNT4KPBCaNLtRIJGytlPk/ipTqQybiLr5GtI0609rE+qmiomNRJWJYHOu
aCXGzyCz39wOqlnkNlpdXAMC5vPGki0HmhbUV566FDVEq5iCz+2LpccXAlDG32we
k0sI33kiCzrqdt+m3UYGo/wol7+Wb8B6QH6mOQQ2LS2SsfJUVdENkafNEhhydNeA
GWBSIwdU9bokKcbPR9qcdaYkBeAN8WfbUPABeTC4phJA+5cfcfg7NTjIv15U2VFA
uLKid8fk8GSR6RF9cth5iT2EznQ+hlaoLvGOYmMygqUWkZBLyDshsdxakafoMhyb
aH/uyPKGQKkpxg6qzUMWaQ1xwhcwvA9VILjqgeInI29fW9uMGrCpNRmvI4ULpKSu
bIlXCmN9MsGNeXgYlS3sdBRKoCjZ7OEB1fxxbt/7RJYnb9bR0p+LGOZPMTbtcjAn
o+BaNnXYv7LtJgw+eT8zup2kb7X+C12n+4MOCdbsoJbWK79NP1juN4sm55smZPjg
Q5vQZIleGo/aQlSfs5EUi/Ey+ZC39OH5fLCClDC6QXutwkHF1WIY4DNhPTpotTDB
a19wa9ZU9q+3nsRN10Bh95riLqwasGKITCvyNWpYJ3F2tWhSReAynVv16CsZx+vC
v0w1gsNHTNmjsk5Lb+plRAFKnCqLVBnSvdBzE0hPDi+L6n4gqsY4w+fmBntxICex
v/txms/oRPvX/2LhSqF419s6uVb8VKSBbisNEvJuqCc5xUUj2wNh7GlpqqLYBi2O
5I4t3o15jIPFry7rtrcgwbzSSK1eRhNrpAdrs/ZYsAJ4KZV9wcCAH5ig+1pXfE6v
0qDnIs85sUNACQWrmJlvmtnRQLoK9DyakQ3GQM2hV1Kywwm5G/yvpItPvjgzoqU4
P6iI1TOptmw813vfr37QaPbMdanlegpVYKz9pKkzX5Y0P5BJQr7wNu36W7P/ocKB
zsHPh1YCAiRpa6VMy7MK2wb9o70f7uCXz1agEKUOC4sJJwnh/FxJgjqpaJ8/gtWl
yjxCPDmtl5XSEQs3tKnEYdPudKr6riSDdPDe3zMBGEsz6xfEGnpvW91kaJqy3rhU
Oy9EpuSDpJVz/64mJh/5dGPNpcI/S2BPml0UOtxLQopx9dXasB74qd5jDnf7F9m2
qrOeu/nYE+3LXRoGW4GoHBYWKPFB6gIgrpjjZoODt52gkETHBrivFIEQDP8Lga+M
daaeoLG8TU8rWHOQa8YzNpAWUn/fpKW24wcJ/0NTlk30UFoRalGf8Z9L+pcKdmpT
L0YfPnbFr26eVW5TfAgHkAvVCEj7AahPdIZyqQQCmilzqbSR8UXp12KpCn2VS/gk
lzJi+LYAsodAkOvrkuiAQWi9eRqzLEOeOJ+ijBxfjdcfX7aRYJ9olfAk92k0by1y
hw6tIeOlK0immEXk3JprlNZUQBh5Fga9rURC4+dt5OzSGBwk0u3B8flfbSz3HdL0
jYQ3Je27jhoFYXDS9y2wFa3KeWARxfo1k7xwVzUWquN1W3Grr/JyTZAdJrZUehp6
TGiRBv+4/jQJIbALZRDRa8bWqya+1HSzxmwxZ6h7qOgcnhRuLMhusMygxaSGaP4c
e4qM0s2s66R4lH//OzhVPdaM02dZovRFcXEUMjbrrNqhYvk3sEK9QDk2qdduXj13
BMstEO5rItVXNxa6MTM1PQHp/Ikq/gjjnPNVOcStjEcjQKwhNLSWTUQwYgc/uhHh
VquANt1dlhSGKzQqRZB7/J5ZNDheONtbD/gliIaLljPSCNogf+nLhpN3ppa6gOJH
2rOS77k4SQqieRSQPHw0E1/JF7xIVvq5NgDx3Ufx7rElPqCrIL+liB8u1pGYSTFW
00YEJzxltPtmIasA4ado6ymEyluiyB5siKsW99dVkw/jqpJKWbcMrcoEEWYkLZhj
/0yut/OZXj76zK7YAKe1Iak4OzENZWN+E3obHiTjbv6D92aQ/ZUE4h0ytA3SSkjP
BGObYVgG5OZwbVEGuY9DVnfis37zcPEPQp+QNDkv3VFpF2iLmaRp1ZkxHhZ8EXI9
XIlb1KVfYnG46uXTJ5KUdJKhQnEDflU0ZMbwQuYbbJsa5XQzacEOkUoPhNmyGNHa
+a9kK2QGlDaELJmX2XuwvpBEnH8Or2E6VW9PGkHaFAxCZNgNS2+7HLZqf5Te4dYB
DBIffB4m1Ub6wgbEXaL6bHoVFmKfqKHzaWHjX6z9HCdZ8ggmccFSze6oo9yu8Edf
R3pyXt1wRhKBHc55WABPFXwVhWLkHZhznuMCEcSwI6UggwL2I24W13cTgXoBzqie
yHG5Jc96kh9Apf97++3nVwR9nHJxIeZNfDwXhTrJSznw9OmAyi6wWYVIfs8gDYuM
zGnB6WAdfHnC9vlA/bN2gwRwcpkHTb8Fckuk5B5lRwOdhbIDwnJf7Y75+f6biBO8
9zWUDX+Pj3/tq/nbcHqaoyY3h4I1PcW8N4jGSSrOO5P2Xe78KPsWnNj0bJQ66xQ5
lnWKDSKQzTwnYJNRG4lws0QVcYqh+N2ggeeTxwihfsRqXlEBqrRpeToarZgL9dK/
TepVIC+qoawH8HxjJEF/Qkhc7mu+ayUn3dNT1ERK0HPe1+JxCzn/M6QyGc6mKunp
g4AW0Htlzfoui0E7YXwvz2sDW8w4HGhy/zlKr1dK5gX3BUf7GFMZaEiAss5tM4V9
gzVNKifXium/8SPieWjGDvybdTlwD5B2dbcUAsySNprX6OkDt/wq5ZBYFWRNSAii
FRSJWEuWkreor9eppotwyc3XEFRgTRewj+e8xuNCcWHzOmOMWxcs9Sx9dKYGJllm
PWTHRzX17Fh6qQSOkW9wE1+EpT08t6BEkquc8qNqXUhXXXNI3PWPXXw6Ocxo7Ol2
nK67Zxe2kmBQ1DAnKPK7uFRevw4WZRffFSds9c+e9xQvmILnCsUH3nhjTEP4myRT
EZB5U9g0+hU/AhQLsXCmZ/jYj0XC6U2LivRLSrY06SSyZ5JJ2R3SR2TltX1MD6D9
fPpIP35XLGpSmTFm64xGgeJf332mCSZivY/1KSCbdJRgOBy2DhFZvaf/2HBr17D6
6P9WC+Qmi2ggijW1oBVr3SufpeKjge3G9nOGglZIxRCuQUx+WLfyiGRSVHIvV4QI
cd4QoYWnE0ibvJ6N98+A+BrzLGMSqzd29WnHyU+fg36AgK8gERuTioq1xGVZUUQm
OiBESJPvEL5EOaCJxPKlWu2LpIAdaxE4KgjxWGc6Nhw47XvWjeCVsZjNjAUWeetP
tV0BFdw9Uke7+todqRSpiA==
`pragma protect end_protected
