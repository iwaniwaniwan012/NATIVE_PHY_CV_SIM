`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nkmihqXcMsCZ+nLlUbt869yz8/+Ntkdp5c2G85RtpZTVqZWX2xC3UAomjM7JpMU+
bPdvspLM656JE4hbo1fxlbLLWS82BGsucWHZmchvG5UiOcattjT0JJbAtPKKzODY
odpTJd5kCAlwSClUYAwIR/qWhQD84mc1wmyIHt4UOZk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4304)
MO6uontKNQfhoIKTFrUTYigyPG8GqLFGBu7vrYcBpnyb2tBNfysf5sYH2XUBEVRJ
iDtYOevAIg3WPVQ4IyXCAwOimb3iZbitmLN2OMApkQftpi6xHctn22+UuZvyu65O
ug4k+4d795/HLDWPW7p9pFcYoeB/x6wxFyo4aDkdTy5qX9WPs7VzxPV0cGx81F41
yqbRn0q8TzZiiwkUJhQqUgQV5QHjuPQZZC6KQd+R9ha+ACQrG+Jb57iAcqe9Y1kp
hUGmQKg1oXiN9B5XYdBcBH/eMSj8WjzZq81CUHuAbWZq2aDWAvUdqFmwRFVqQBNs
WYghB+PPfhgAxGsN/nnTVFgHT09c+jm37HaRkjqiNTu9F6Ck3C1594Io+AMvccA7
598UB1S5dDhPCx7teAy/t8vZ+zb56cFNrnZ19PcpBtU6Sz3ODmPX4POTV2l6xrlL
xqpbre8O1mxNIIkTPkLdHmWCg2KPV5ynBlqNSIVQJNG9rptPpaWM5c7t/X4ecsA6
UIbHXT0mKdF9u3JhiE5bzRZHMklCiXELrwSJ7No11kN7izgKU77ypTp2vONjllpK
vZve+0Ka9RkOTgudUuviTs94eJ9KEX3sPLAfe7vsJAdZoKDKiygJwpLsYrZlK0Ug
W1bEp47FJLtgUCA3N3jyylu3TwseWljEqd/feGyiP7S/JAVRgfSINXSfvjekzo/D
lXk7x/gDDLKOnrVBRa1N6Dmp8hzpAbnPCAdXoswBLQutWxMduPnGS4yRY9vdXO89
UmzQ9sNgahUX7BZBw3z12pGNRZUkbJu6xTrZV+nmfQUvzlh18Fc2kr009wQZu9LE
IbCMs4QAKuAwd/4GOr7UlP0aaOVZKYwclAuQmM86Yxd+/FCCNoCcJ/OrZ1o6Sgu9
OKrCJ8SP38y9SGbmDfobslWShmASWspmjHB4NaALUnBMTH68QBqeQ9gU/DacRkDI
k/vvmymsC3Oava1tqQt5L/QIFS8WmBFBgjJo8hAem+qgaUaJGRggsSCPJX5rx5bj
lvktlZYotUvlVObf4ongHgh37YiyM+Ir5BLpBZj9lywADFiBPotiqrDPEqLdmpvJ
iGsVrJ4HG3bSJho5t0JNH2CuSGUzXoEJCgqbsUJZ/E1AQJzQWSU5vwzpotXK0p9X
GheIBGobcsgWfQEyM7H3gOr27Iot0p0cJCJOmgqY6vAharYNP5rh0jh4lqa6Snrl
vGrvcaUTcJgdthZKoyTBtZXLbG1qtbHA+6JLQFqRuUoprU19X5REje6XWEoqWjPc
NncMLvgBQCd/bRJH0C6c4oYfXKRyB9ASMeL2hZHG7dDnRdUsXIOwhrSOSWdMQfIY
MDpSjhnRd8i55OruuipsGtoWrTwdJw4P5/VdAfmnDDHoU/N+5rAby7EcKdJIyyJk
RfjUfkd/5+GiUToypymaWO8r0GHZEZOCHVjRG7w0XI0VvGUcRdHjTJRAPdPrEuld
eLsNFVqGJohZNI1EuUVljpxWCpjO+aQXujlJ59rnV73lS6AhCeZoHlkxBf/PotlW
VFxPBVKbHHj51wMhHcbJJNH4G6rowHxqL7jlLeXpKhHe53YHwxbK5/Zb8ner9OML
47JwA800rPI23jemX0dQog5GYBiGH1rzepFk1PQE6IFRq10vV0tJQj3bY8AcKfi3
k5JPcOVk/UHH3mt4XuiC3VFLVoEiObCIIFZ4CYVKDnrWfPYxB+iZAXlpXTV0k0xd
CiU1gCMSznpk58fefTmsF/jM64H/vfmCSsa9+4Cn3Mlh7w5kt3PGiwIh/D+Q9fzo
mhi7AGIWetaRCtizJnbrXYJ4LOUZqPywMDFR63fRFS1PBaQxLUiZ24AQxtZI4pMX
6KHBCijnQfm4dVqPiANPjSIOOwMQz7wKZEr9i8ukamE7F/eX+8MsYuVSrzEBqBIq
nhNJg/x+NO3BtOfCbAlhQ6jJFJTZpO0zvEbFEEnNRkXQylvLHTZwGw8tCNKg4t2f
aOQ5a2M/NaM744DVEJUwhy94k6/qSXxWAng820iS4cx22hucjIsPmTnLQ+JC0oh+
/nmmt71D/uvUGaWc87/ZGeRBHFkTUgHnv6pzw0rcbb0khDJlbA9vWkxNkAm+ufDc
KHI4D9QfBM/ORcmkb2DGWNzJ7xVXVtFDz2AziecfJKu/4rgbEgRl8WaG7vgbEG+/
MT0fDlMVT0RvgxPVHuYkrt0yAm1xCf7/OEydmxoVCuPs/M/OogCOd5FZrgQgDieY
1sva9xzlJgIGoQiP6LM/c2MPutua9PoD/9UiB3mDbjBAunJANqbFFNv5ay9bKL6D
hkeyFw/qypfPdbznic7TBqaKt3AjrXCqQVCVCrCNVtP2BinAGM1zSdavJTaq80Wo
ezxkxtEB9XFC3k9ovnqJ595KZqcuSMcZyA/G0kaxDPPKlYi7VlBtjX2XGvSy0Njy
UzVdCHXXKqIYzjl1oHFnCadvBJA2SGir4RuqBzAQATQ8V/C+h4nIene8auN8G+n1
l+eab1pLNJJVlD+S6fkWRXHrwds8ayuTvcKkL1n33Y556Me9j6z1ZUp9N81wWCQR
IiDU+hlNBLosh5ogLm6CsuBO1tPr5NEnXHe+XmEtX8TK+LFtlBoMQd6vp1dgze/8
9/H/4l72W4LBtEs+J49RU4qmDVZI65yXxP2eYxEhUW7adA+fXSVPTgZxaKvWeb2e
3GopsfafTkSaz1MrcKOyPPLDy4xLNs05vjVvlCWk8+uGqUuKbzvwEK9IfuDUUHjU
r29WNgkXRyEdw0PL0QFNQ/clIVm1DIFnAEOfhpwdvBl5WkJ+ms1MEzKMzZ+wQuQb
cLjvoZEjQSpOMg+End2gJB4KhHYeDAR4AaMIsImyhRgLfR8D7Lm02JUWJ80W2UrI
aOyw4O3r9izp+vtkHVecRiQrsAodKmK/upjtkM4Ntp51Frp+E0stqTuJ8zbZi8TJ
TMkvKtH7rNuRFFaGV7W6QaxwCl17hwObJFYk/Tu9UAnTQ6j8H17BOLYkz7jq5o6K
GtsKLjb99MtW8tZ4fssSgIXX8kaDkZH6RX8+Wfha6nr28U1y012D+tVfgBFHnWhx
UFDHMVMA6S8henkgyqog82QixfLjORH5XEfV22aZ1WfD7J5trV1koISC6w5BORYS
JWYxL/Pw6ovDgcHj5PwalMAIvFftd6SSxZf0eItW2cSlMkM4bLTrMe3WscElUPsy
5rvON8UGE6YOU9O1Jebc0/g/Kc8C+W6oGa0H/JbPmIxyJxAYEO97wPGMh9HgcQkU
dwJ7dIThR35+URKjI2Tkk9eytjMGG0KPYHpMyrWpwmLNtSKrQjUP9ZfRs+Ko+ELI
xMOmCatSDRd5HHm+4kOuY4Q5NzMKt7m+2KoEI59n/rAJIEBB6PAUT1/F+y/bjFOA
w9pkULnhQHqMeRmpWYPZDlDItsOhUZ/0XcDxMZ1LFBdMx8df8cwoKQyHLeWXM3SB
/7XcNB0yxwGPEWelgSZjzOnSj2aX7HO2abLSzaSnVIZw6CCzoJivndOKego2OSXg
Jtgf1pgfKqZwgqYuohOID0BC1szRIlS4iEttzRCzcX93fjd/IdY9wk2qPuJOoYAR
xnTbm6XZl/vEThFCM71NQfrguDpo1px5VGKNv/85pKvyPdyQ3KnZu+aq2eCmuVGH
hZvw8i4Xv5p1MuVsdbOAIpmQsQHAAVi8z86RxdzS7kgQT1OG5aKYa5vq2sydLylm
c0ReFAPEc1gvGA+XWsAi1Ogjowpdh1ylaGFvMFabkATh3lvMhuOjZpYFbaUDFWpL
Eao6y6DtiEKck79pe6/Lr+kFMqFkiuSmXROKQtTWi9gROv7ZjKlk4RPo5omKMHz8
apLsXraJv2aAyWCJsagyTIbX8mrDhaHU4lRQ4okSbxk94xHKqUlBA3N6KVxkOTPv
7zIZdoVLpsMm2Jrk5PoL+Hf7ZMQ7V+NHzLRv22D/bjF0XFVdiBnU5PNa3+4f5Xd3
U5LPrsix+LwObkjTJLk3+OqwGHMifZcPl8dfy/O1Ou9Mcc3r8WwPxmOYIDKZaCaX
IVz2rWbGihX85jAE6o71f69abiIqAsgKbSgEmjpZ0tF4ZliQC+b0x1HxBLiRMftI
ehKhF8wVldgbLa99biykeV5TCMTfxI67PsL2sJxDABBTfvvOecMiZ5lqlcpNJPsx
JSpO5Kq+r3VjysP447xnJREim9Yb5m1A0E7Hgw4JtCwx9VQ782N2frk3tuuqCoZu
WhIUbdpzzsfhhHD5y8kI5r+KQX10BvaU2jPZvUyMBlgRqnRGqkE1R3tM7KdxFKqP
+2WAqXgHjKzCbFT4m3TNJnTAMHET+VTpvaKwf5o4kiqumwndQlECjuVliX4YRL/h
KYnEtPPiI589WIU0C2vqFp0K6WCgaHp6d8TmJlCs5lTn0uftA0CuaoILoU7HOq1a
AXY48jFlap3MAvfB9wlek4OO+Xl58lKHZHabMHNMHWTnVqzrSp+RVDFAEXHm2LDL
Tes+vXyLMFv5JucCHCi3KI7bwYCfpzUXV4s2J1FR5QIGJaz8oHkODyPMjaVC3vnA
qxbcEncqp6fw/X2oUWlKE6KI9G/P3DUJG/EOmuUIPlf6/OWc4oVkb3dHOg2pRoov
JqXrths/nIv8ar8qQcF/tLhetPsDqic1sb5+1VFXgnm1+gkpcYAbgq1dUixx7Z/t
3YgMwPziCf03vkA5iHZNO1RNCEXbEYnFC9PCTG5moucZ5AVOCOeTdrZXm89e2IZL
2DX7CgKtFzEE7dq4+gyvM/9YpP+g2/YcKhdUU6U9TuAKsY03/ODnGol2MR4wJnca
CpeTj8zZBlknPNf+Aerlfn5+pGFHX0Uo6j0Xeh8WCowG8BQiGOpJGYxcGyeQ7Gmt
JY+kUfy9QIe2mfyNqHvhHPEQG+V2qfxX9VhBdsJoKaBdSIaETUqaCmsqtjmvrNaX
Mo5w8YElsgIEVW9YeFkHCdXi18+WiRNi2c6nFqGWcYHhlkIqUROZllnufi+MPiay
g5gEbmpuHWvxf+f5nuV6SxX8CHTGd2EJqz0BK5RDYjjPsiqtuy/2AMsCA15gLDzM
bFpxl9d4Q8uxciWM3e2+KMC3dWpeW/j9oBuAV8HaG1kYrFtDSK/zYC576Ud5B+WD
NEuzZEqktY4qnOga9wKMcWeQW4Woj6l4Cgq1JPBEOVWNnsKfjgf78MqwdHsC3boD
QG+R7rm8jIdiS6K43/WJ24SK4R3W59iTijJ726RbX6cZ+IJk8BHVbYwOG00WhslN
mvKnqzhqpz+jmzVarXSVXzEHrYPCUjCNHPb3COSt+6oZi0mcqs4ubw7ZEZa1LT8C
uHxAvdcXBeW1wR3kkS3rl1+YF2ldNw5Uz8WrdbcFvQ975TLk0eT7qESySJ3a6UXM
g4lchJhiQbJh3Do8aA8s9Pymq6o0UiaYM1L8jCxO7lCDOAE4h1kxDXQTFuUYy4Ob
genHDx5rA7rAWQZDUjgzMRuBSG/Ywiylm7YY+iZ7ga6ikRL1NTCRnk6K6x7KAjKt
wgLXXplsE1+BZbFOFJ/pY+FiYgL+LKxyjh1fzAwQTbyaPKp6Vozb2x5XXwgW4TK1
uzZNtPXBn6tlbAPM+px0+zYZUx/2pVeXGXyNdDW3DWvZ/OiJB6XQOeGd0W2qExzB
GfM0ag+OphE79FBPevBPMKbGGGJCYZS399RXq59ma+fe+cV3aLejGTcUDDbq2WKS
bUBynT0hNj2TCgnbV/vLZEovRcAvlCETsCV5ANpLCNY=
`pragma protect end_protected
