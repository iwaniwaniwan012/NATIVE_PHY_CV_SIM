`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PDX5U8mPXI1UL/cY+XG68RV1N7emR0QOhGbTqfGNnr5LBZwnXS5Pkomj0OWw73q7
5jbhE4xqyIGuThfKd25hsI3hRMS6GPsrOV3MVXY/PKdCkdVNr9u2yEbPb/sRs8Kv
lpvGB+GLbmGAg6PCm6BGYnAd2OmMsQbULnLSmZPAXZg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7712)
vV5AkMsfSsQ+gnqCmDxlL0F1C9EkyjKHbGC2ZJ/c47NClMvDP4Rhzw1hW5s+2aw7
JxfQyJVCR5v2PiJDtm1/17WtlA9Y9ctRwQQb9EEDR48cp0N/GrSxWIeYV4sedUeV
K2eZZOQll7E52S8Vj5+rYbraTX6FHF3dNHb9bIpxJ2UHU2h4fWOfTYNyW2ah0fiD
A9dY8ZolwD/mnmenKLUr/C6uM56OT0ETWbdoCgGjjJFIaEWp3Jm3IG35jiY/45cr
eThrNMT5tuGR7oA0lp1lGacA2DrSoPgQmCczFf9piEkg6tujrfXn9W8MIZWzYjyU
5fFxI35CYimAfC1FQKurnYfj4DvWYVQ9w/4mkww1N6hopTAtsD0ZjSY5oguh8Flq
IXyinXE20joP7e3Q8Sfe/u3vdgkdTEEVCapL2scjPMhvWmNlfT2S6wTO0Lwcf6Pj
uaa/v1sNacFcMIYib5cbhJ6pBpGs7Ig3QGhShaWA9P3q7vKIYaIQSm5L3NZCUo2b
kgEHj66qkU+gcEMcgfhvTxLsQnXKxGVsaB73Kt0F9hG4Apyg4cZvmR9hyqe2Ga2G
3fxx1jpwYx3uMubBfZEB5dY/42AbInLSxS+zZ41PY6nbLA8zlK8rifKaL9oxnD1a
QKpSEIyGkcdLoVI8pYl+zTtlVRHo5DerXG+NiE5asi/VuyQeIavU67VqYNq0k56C
N2mJi+Pyc4W2S5qBaqsB9WZ0gcNLHha04Z701an6KUFx1IqADRlHdS99h265d8eO
/qVBMUn0K7ouSxayNaiapBl01Qwm+y0ofM44nu8zriCqdhUPtsgJ6tH+rjIkklzy
P7g5U8TRPkMlnYbEBVhrMc1i5O6gY8/nmiqZgb8FCycwT/UF/rHdHeofuKW7+VJ/
JJX0FIppEHplmcIWk1D2HFoGFnlq++h/j/qseJ7AWhgpUZAth6AoMgrBgqKlNX9J
L9x3EFrVO3Zo8fzE7K+i7rIiYAeNVwkLbi02CnTjJFHl4y/o0eEoDJfsHjsSc4WB
tZiBI50COWVRkQ+VS2ZKA5L9IqyfkE4PTDkgXMZYNzHGqF8OOEGZ379nvu+NSZdf
3vkTgpNyfdKQ7HyCpJrHKbQeRRBL8nqIFty+DvOPLKIjqGSrHYAZqumKynLbiNjh
gWiIccxhhsxFaUL3McbHBAP0EDhNCw4KafG399Sk/Kty4ks6NeRq3B2Cx1sba83C
xHqCfDBr2xWffs+rNBZ2NAwMPJ3gHNLKR4VqFK/fAxI5YURIrZurjROxayxOeuqB
KjtAGrQk9ol9sUkQF/X++Wj8aSNXEbdOOgTsIY2h56AO3jP5zONq93mnmLDY2iZB
ARpdEYCBYbq9Fgoc9i4enieVe+kGdcAsXvEh7N26hKDNjx1O2MWQV638P89Rsq6J
uz97Gppc1O+D4gRXqQUlbJ7ExlGR2zKB46glO6gbBf5iaIVcRtENC5adjQaZhixp
x1t973bj/AGi1QwzN7CgGGJ/2YTMAD21JckPE+hqs4EShuiMPe6IhyqExG+c5DS3
BcwyUpVZutGbdgW5B+7E0qgoJukvDAdt4n51iRoKGESLM2NGM89j359SoYAQbHLb
GCn5lgio5nay9mHFuS79+FmpPZPZCK4IIT+QFE+OssPpefae9uCbaAfUUM7GaSl7
9Zo7cFuhjZKWzy3a3jvXCNurRs8MCWVeVHvMHhBZgf3osvmmyNN1Qu7hUA+Gj3Fb
5x0Oubta+7we/k2qreln0Ci6IGA5z8MspQhPzpgTXWYqV+tVQj/MEE63dTamsvz4
NoYmDi+IxyLUxNewNNBAC7X9SxXq86qS67icJn/T9368m3LM1vV0lFBoCJQ4WCZk
K9tGfTk9GTdcMBe4KM3lopocwLoX0FQON5JflnNugxaBCmL9vSGIBu2YNFgg6VW6
1tvqGUjovBpUXeBWD/ju2yllUZUON53eLrLBwehBVUJdksfQhvZoqKCqmAlvIphr
nudzHi7nkC0YRHHXrKMqQyKLamh5sEF7oF1DBilmmE8SOHD2yuW/GXYrYRlDA1xA
/lPjHHYY+6Ago5gmg9Mm889GJL4c84o8R+kASu5Wj97JVr15qKvUkzOTy/P1DO/+
Jvg5x2eqtx3ACZxVgKD7YPZHfTsHBoCFfEx5hoUvDottPQXQ26i8EL6homvlEIvp
lGx48HBFv61YSBr+LZRHDqyD2lm0fi8vGmb12qW8iObBI15cjOrPWPLnqCm8pIH6
BEDhtoLie5hM+9kZwYcT2fauusRGqjwqS9vpLLgEMz3XbeC5CT4qvdI4EN3xz9A7
ww2Y4e9yOhj4+wRnnq83pi0kLLvHSjjvq3osO2EkjBsRGh6y3+Qe3/uGW19NSrfX
BYpzkzOCHO9pe2mrPfXcNmDIcuN433+qkT1rlwjo5JUJZmAVovh3PHOSBupGPeHD
NSL8Zy8PdkzsJttiCQ0wgXur3pE/xDdHcBGHNWOz3D389sN/3OoZqm/zhbSe16XQ
qJthdf564Qf2DEtvD35qcXPfnnerlbmlhEqR2roKmWtRnymh3kAllrTtRFMAOt9Q
WWnZtO1++SdAhlDGQz0ewAAJInOBAl/9UwufSylBOzXHpx6RrbNwQV/4EkIDRzE1
vJO30TaAs5K7urybqt4CI2HSmxIM36P8TNI17e7aIMZPW+3baEykiB6DIUEUbvyW
zHLD4jOxoZiEryxLdcOBNN/zJRIHfXm0r+878u3oS3ZlR/im8NLDvHlSUWAEMgRJ
nYsZznnOMGtnUHRj1bWiiy13SL8uu8KMmMNd/0igxA0OVDOfjlMDVLpCYyKtUmzV
oD0YlhiNZmGIkjyPfNzml6M2y5BF4WaL/qDhslyDD8ofDkivGHRbQTXnQgpeyUQw
lT2NPIzGLgYpC/+7zy81NGAls3Qhzik/iUcz6JvlB5rUjlYcprqWlMPzzGadCE45
r4/lhQUM/V8AXzOB1FfYW5An/pKnDa6yjpViv+I8PMppHCY0A8wJqfZ/NFHbpJ9N
zr+o9hnson8utMP5dWsa9vcrrNwZWiWb5IUqv4fsQOtDQ2AtkQ+6sHv5r+Mc3I+k
w1HPRjrGdlzJmMMudzVrMzEh6RakN9SSyy5OtON+PF6AQq73hVvz89ZANmM5CPru
/KMA2PZ9dwh4WIBHmitD2V4uz6aEFrrDM1efqasR4KaNB/s8r7jSsaGYJ9qI7o2Q
y++dNZGDC8BljHTJs2iJiOD9XOuqptqXjtoi4EJ2IMZUW5aLti+UIhPyvSzb5Nmu
b/hhJSeoFZIpakKG07xVb9rcLcpLrBOVUSBI7SFpeCusxcNc9uctE7QBrzwewaLw
kFjTOpBEPV9YgRDtsMJsD88gOg5wDtezH9D4lTTz+x2z4CyqYfCWA5U8FtwsPjE0
h2uF94pFzC6a3Qn74Hyuodrrl0WTgSv4yx6PKvpPamoPTt7c2wPAgf5AwOJDl0VZ
6MLKrXwubzCnH2HaUfpo0bfY2CP1FI6XrzRPPK6mOiioWl81nCaVqf89TW3w+5Ui
QBUv9Yr+0Donq9tbdOtEfMIe6YhDEV9mgS2aj1Z4Mv17182O9ve3PyAyjEKpWxng
D45JIvmkAJ/K53Ow3Ilz0PzwrTRkEaJsAXjMBmib8ALJTUWu1GNUQ3MpVovqdZQG
Wtd6ndH4vvvTzisAGQ4FYco7lXIKv6qRHowKUhoA3jM2DLjnKzEMaprsRihHluMY
Acj5mQSrIWG+S/Cuk9TuiciC7LA6wnjK8Nk+7MG7YY5LcxpY+iRwmruIVnfC/skG
jujGOPf0PXFeT9eRjSXrTeZHK4tpBGTgmmyhGrZ5pveX8pAAj/ThPAqbLbfXtzgm
eKdZSlmXo0qZXR+SXj3t1zdP/bRC8l3RpleHa1VC92Tl0/xLssobueVN7hcS+czs
soKmGtAMrrrRkmTNOMIurNndL7fglRL7NFU/n50Qz8UEjD1C+xiKAUdNnsf/ZTH3
03X4Wcp7fu1qP96a9WPYWSNJHsd9Gj2qkBglHMzAeu45O6kssDvSFsyvhP/oW5WU
0jF8UOFfuL6Q8Io1NtL5FQdSIjm/pzqD47g8n2m09r/vCPlJBJWxlmBc9eiivFoA
rkjbChZQGPswEkdtf6RVutmsodJL0rv1Zh7Wg4LpbRx4MntfoOAts6F6DzOk3XT0
43saWiTGDFU2QUAbEoE/WhO78lp7xBQs5KvN3/px8VJdi/4TBV9hluAi4B0bA5tl
cipZUhh0/D6EReCqBFQLNMyt2B3LITROYE6LKb73JIPX1cbAO1iPx0XiQm4rCC9S
Pr8aJXwwGUPKCyCPk1MiRo7MMcmI3TGyYuDSsABmNwydZZMOYIcXDgx52Oj3xXEg
VTWb4UqCiODjNHw29bWzwMCW1cuSMSynE84o7xZTkk6cmLdObdnIr6NOGzym5cmv
nKP8Z0109fsF2VwtEKQ3g3AziNbINv49ZilleD0HPaFyz16uGb6pq8j9duU81Z38
mwwll8b+aq7VeUPCwXuzySKEmUEa61EnDaq7GiYmY9xOuxkGPwtu6wCsGsxxSdof
yXUoiBZCCaN6nuGKBG1505NIZ9k1duXEXxw139FHxs6z89rXAuVokP4eabmvjXYv
fo8LbTWdw4ou3M8jqvOn3WqolXq10C6N2N1L1HrisuExheS+zmYR378rnezSOR+m
97wlJVOlAoSIijLcgQzFRI8J/Pw/d7wGqQCaDnfm25VTFlbBlDnsrFc0O/C4fviA
Wc7VwwB7ikVDKsclXu8GfTz+teAqUGCth0G12luMj3dW4f2vQgHh2ErbqVlTkZRo
i4T6BXA3cfcW+JnwANMjK3LhN+ClIsVlFhUDde4fAOXHRryWghfP0c6o3LHUT0ie
B7pD7pu8nsyieKC71z4HtmcCNbFQpiDQPZyLczn2vjkwsdsvmJK8v+zh8tb5zPMg
bQuiaq6lV3AljxWKm+jRK1+8E3nf1fNQN4hmfHKUkfMpq3ZNOviEdCA49ULqORN6
7k907ITAzqBVJmAkZi0mjkHbU0WwAIq7l8pSlMIMqXK35Ea0vybjPWLz/0cQgdCs
giC1WMOT2pygbNBTAGgrAuA12mBOSglwzvGRt/ICfPWbBN8rviV4spKS8mJz/p6c
EFTb2+2jzaYxpp27lhki5Lmq14GhaavtYA/XrdKdqtNEXXSqgatzTJRfzUH7EHCy
CzSl4nBOCuJpbktttmqAeP4g3rnax6RG24d6BPOB018zKetxIZMe0YY6qnRk6R5t
GLtBajg2TQrfwc1nAhKk0roBnJU3A3MFP6iUZMyUS1FefegD90SsVyPGxrcUl8JB
Ma9K/PPkQ4BGWuW5VL7rf2bHSrOktGUIjp1sy9+lKYM94+uoOsXhnIcVxV1juoS9
NMIVZxmAL46rX9n+uH8uhogDHfgWq9C8xZh7gPLl6wgosliS3b8fzUDh4m+3hSwj
0p3iKOU51g+VMC0iR1edrPU5zEtoE9zJrgfuz7aB0R76E+/kAYVK37bUXPwoYRn8
2tUHnkf+YJmJDv6zUImJf6cC1V+UzMZYN0k/WeI6Gtvhhm97tpZ7NSkNet+DGNQx
z09DyMnqIBgUWE4E1TRF5hfouKQSLm7Jvr0uSAqGN2h0hpj0rSpDOUdgmqw7Pjhy
Zkk+rH6KqxumFwWvxgLtg6uZ56NsFVbgv8Fvtz8brTLX1LduofXdQcCKKwBjaHL6
NVh2nf5huBFT6UxyIZe3Bcnzjsi5/WAAIN2CaTMAvp43O4Ps/lbltJttggiKnRB0
AzYDKXGaNDkkicZjkUARcrrvahIL7MsuJ/p2040jz0JDdB7MWZ06+NABpUC9J575
gqUns6QZZNURvXoE3v8x3u/G4jbRJg0QwYSmjzUiKr1PI9MMDdhpLReZP6OeAWi5
2fS3dxYVfMIzMn6xgkBHN8f0pwDycdnTOJb8AVLvwWcHzF6ER6LPqRZyBChJNdF7
TzFgZf7+kBe8E1NgIZnauoXrD+zpBQeOAQ5vHgSOsZaVT+CBP9vsvTIUSt4OP9b/
XJx9zK3xLs+TbFI2vpejtVakpLv2LhjZvN6p8PBsduH1qoYkqxgNJ3/2etDTWyxg
azcQDUoc0Ft6cMXohtptjt8MRu0HsRsD/YsKwXVq52OG/crHGvZd6H/8t/CC0GBe
7GZzJApyia7KG9Wlk2uMkJkw5qN82FSyCNCCicGp/xt05JthlcOsb9u3BGWAO+4w
2JWfpmKVzK45IKGlFeiuZKPMhrUqKM1nKoThHNYMnelFvWb7u27f91GFq0obAQBV
46cfC1B7prkulIPY1WdMmYBBX4/NVb0z3bwXcFe1Ma5+HrbTb9qXGWGGCW4YjyeX
Mr9dS9r3sj2Vx0g6z/pbtM9nKWxuFBkEe8FIZHIor7ySLoRNr6KhQrFz5B9TlV3g
RkI8JNDOcElUaem12VEkAGy8g2I0F153+Q7Ye0K3ulxfBrIarh9rihyMemqpObIy
W5GUBpZIRSxnUZSjIldOMYSjD2LXZSro0+zUFJarhLT6luQldb6mogAaAhwx+hZv
LZZ9reiRDJEvl0aVHQk16rom6jPoB2VKLyZ8z+K2iD5HYHi68QN8FaRp+oYfxZIU
KfhZSMl2TQzYq4z3OqdQwi2d3aRTqGrbj4+d3i0+pKukvJVsRU8Td/xIr+JUEcB2
/4KZC9YVFKipz/klGHbdVs946gYE9YJVQR9uCzGOfyixdJh2CMWf0uBxWW737DRW
+Bnbj/kEc26GG6go7/Ojfcf2FMTWDOmPuC1a96ZZlmAD/bBzSPfEm/ayrByvaeLD
05paTdnza6XcdpasX5PY3P2V6hqX95AOin+2Uv0NJRu9HHfTk31YSlvdRKjMZn8I
9a2pDTYauuWHf3MUXQa7XfNQdOEu9tnvmboETqSuph7xXJvlT956RvfxUYakaOr5
VgOkVJ7v9QrIm0t9ju1Xnr9WmPsPNqq2y/xLoviQUBHZRMt24eZRQmX5XF42jkhq
XDUAM1KcL03+tBfGms52rS8ze5YYlSRDObc0aHb2keVK6+xZNS8lgaGSYQTbI0a7
r1QIeqwxUk0tICIqLOFC+xS3xhhsHWlbLXi0Qa3tY4FIiAKwu11fRPx+iZZtvosy
Plvu87K3YxULga41UA8EKvp3YFaICsSDkTUecbpU9E6AjkcFolQ3bhuQwJn4whdg
z+oqzDu9oXP1zLv49qbnjN5gUME1+66Zop45tX7kMSmSymwOuBUwWnPfneM1dXhE
Og9DSZtfaAaBW/JzwiypCUoLKlzhsB7Q7GKZF5BPKyJh9KJEMjMCLZblxm2QyYlD
BnPfY1wr8yyNn199jhTE4Ua6rkQAC/rHFHWlfsYXVfe2mD3iTXsC2LUFEDru+Nyv
9xAqmPJ4sEgL6n7io+Uym+Y0yLzdi3wDZV3J67HUOiWVmYECpQ4q9GW29PTrQ7ii
I7Vivkw+6bJy5i3Rssg25cYTSkbuj6JSrFt4KDsosBdUNjiLT/ahMGTWI/e13Mpa
5dCpKuD/7XWRcTIcWZhcxGzisCiECo0+DEITxotloz5LqlzRRO8TMViTOnN17hl6
BzeJo8VnJJ8CCwGoXj1EO6Av+jSEZHQj1RrDIMP12ZW76DDfkwRDtCNC28Iwmo5g
a33reK6a9FOLg5cRA8U2M2kAsjLx4BPs+YZJETnCJF2zWLCnGBF+KrDDRVsvAdQz
I1i86eP2D+BtlSmOrHrIDv1/yidQBAn70ptw1b2FBMBwzLySmfK9r5hgJ17sN7Ti
kkdnS5Lx2xqhgNwTaDRFDZ8QuzMMnd6jP+SbOaNZ1ueuGE8eE1f9OmeGvGGnQXDE
eMgb8xquGcIAGjWkC/YJLo5t0JcJCwMM8dcz3Aa0ZQa53I4ibjLrV9iAogD64+i7
+RPqLFiA5flcnIGxoCHIYm2OkoiTLayICEwdGN9CVxGFlanqRVr6/t2mUiVVxR8K
QdsbkSrHF4WEuqsDKDttTztwxpvOfGOmuYvZMGRC4g2b6wsblnWBcKyf9dQXsKua
5+bax9hAn3zRQb1PTmRRGCmIekYmk0pBGtcup91aol9HYMb0xrlfMhRZ0EyCRkrJ
+SM8WGfoQvoOcs+SQAutOGkEwTx7BP5xGeZKXvbnScmYiDgFKTtqkNq7SSzNDQgM
gsFvGD2aBwvgHeF0hnnOVCrjHku8d4ue7TNRIREJjlwQEYIPhGCc3ys1S6jkl8Kh
jepVo8ZEWlgBwDce/4BdECu/nHtOde8x9AUzDJYz9LGcuDLPKktC8bBjDKl2/y+m
4Zwx8T4qzNIgg9H/MlJUG7Ryy696wC+M2umMzJwS0kOXWH5YZbwzY89OMuL2NGcV
DUPPAW2HfB60p/JP4DT20l5jqfxWv9+OAEulAt/diSi5pMJyPNxPd7ma+BZG5IaK
pP7cnQHahAWH6xVuQO37aFCBHY/RuxpZYEYOqP5/yB67OIF/Zl4JIpFjTPvyZlr0
knhp7oUtFQHTw5yFDnumATvn4SqQq3r82bFWMv/Ek4m922xLW43d6g8suThFdux0
t/7/7/L4o/Y6AF3/TzDn9jQD6QK/aOkH4nf1iSTTzddBGYcHpr01OD+9q5q2umn7
hxRW6h5zhrzWU1NECrIzhwb00spjymLZ9El9vk++hIY+ekEwTx1DM9TxnpWfB2hO
US0namQZalN0GCbDx5/3ytSPgtAsq6uxzhHEEkCxzLUxYeOzVaFXfwqJpswYkFmw
iVJX9h6ad6fDd01CZqtVTwSDXaFaMoUg/C7W84PddSCyNRWO3JOqVEbigboa9yo3
R5br4Chf2J3k2a923Wg2WNQBesXxqAi9RJVb2xDWljwWmGu1RiM/VCMMj1KmMHK9
8oEj8zC18e/4e4vMnf6ujY94i1RJ5aCvOMoiaguNi6SkgQWwH3yk6cTo/2h8A+p8
cLo6eBCPxxNIa1dfqut0HKPmjS0/7an/GCUB+8/r4qbS9oni6e4dLZERLPM+yNY7
laOnrkNIHWe513DF5++kJFozpvkzqf/1UkccAYk0zHMoqpNKzUPZCKj+2djKCPwe
vI/OuGk+AIu8YihYA6dnn4nyP+YTYe39XyY5BF0yP7ow2v97OBXODHZSfOOnUg18
dCg2c8P7MdHf5qYErhxbqHshCgTbZjhf/jE6vqL5C8Swx/UQvxleL81+b1pTBLQJ
izkKKAGl2uEEY0abs3U9ItFMRoUHQ9ktUpoGD29VuwqS0EnSb9RiLlTM0xVMNCPA
bzWthF4Mc2UkE+fUV2Q620FKUg3XQ/NbHMvZG+ljbW96KAB7TA5A2zJIR91P+rie
vkEt9SDD/L+UlPLlqZtTzavSwkKUcIyURj7lN5bWewTcmd5OWRUw/ZKLKt1iMXGT
wbyDUrbaEu9YKx1ViWrW5dQy/xMqTojn54uf9me0/lzaeYfR52u28Tb4Iyth8KeM
ywNzbScRvX7BlWnJg4CF9WWbZxJ/litF4/MYDC0d823pwFKhfUdeSAiGFrQCuFjT
cY//C87WQ8ApMM8yech+YIORgoxPbGOCuseYN+qEDYfVpjb0Zpjz8EjXoM3cLQq8
9uEBtccaI0QOesooySXdbKpDhj1Byenw/FX1v0GNG9KMhAGR6RXUeXRdwUKI8mzS
khFscyUshYa85e+HLPm5/5AcyaoDMSeGKA8kW6duMzFpux49DH29bOpNlPGNufgB
LqAmoNldHiP7DRsGvlFcgVb2rNb2AmhiH/nNBJW3SOLSSMgcuGsGjJRPWnYoZGBy
zPZWX7/cLpuJgp7/nC1OQqgnRSK7S3EQDSI2rJrY4DqvNDNKcfn6ZuqKyWJiMjGj
iIwIInOXwOB+R00INzFxRYzC5L0K5+NRXIjKF4Oo+pgNfJ/Lxk96iRZzxQa5JDlu
sqyMZHCBGvSnvq3Me1aL7VQWvkzutW+QvRPo07hJFWxP2J2W06CnoN457cQqJEN+
hUucA5dPbQG6/jELwNRAbpYrSV0vLK3Hds63SmdZExTo6ItUd8P1ZXMqt5Ri5iHN
wiYyEqdFyUVVzMceAG+knozqbjkcpazhIHZCi+6uewJ7uMZyoS3En7rFvu4AXLyj
awUJ+iKTg0+rwIrtWagLz2OsBA9oGyvYOMErj0UP7cSGwJiXeOYJaGnOwb0a8Qxn
JuE6dkYBtMvlAu2sC559ZiWQbZ8IAU2uJzhLfyRcDyotOb+JzJsJd6u5WxF9LV5D
H9XgAbi8X68ws9d5yDmiNsK9yQLWSljdgZnt1zuljwurHAwFx93Ua3WPcXbdcQnL
wzf6Yd34snKtrxoNRrgNsk07PXmsNlvs8d60il1/F8M=
`pragma protect end_protected
