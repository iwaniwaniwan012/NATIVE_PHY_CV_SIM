`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ObBf6hi0iVaVE+1ayToVMIyFe0nGIXgQ8TzdkJJfscvmmqgq4JYZhYNP66LZvZVy
D09JpC9z0eTpAMHHAFfxp4lISeZKyCCOV8aX3GbgzlKiJFZ6dMS1wLfM7p0vr/Ta
pROZWFf4Uo+XoRtw+c5+YpCQoavd9J1NAPFQwgx5Cdg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3216)
5CcGB+qKt6/8MKNDbwEpDjzGtUFSKaCBEWzneMTZ1qtI1+NRcJzdhddy5jz6eL62
EWKHAhqZ8soC2PtM7398a8znh+HLS7Ycj1FiC3m2+Dkbfa3iJox0mjxgPvPUW1Z8
9oMiB20TT9/YEGvrRR4zxJ5gMvKdf5DEF1dui1U3DLyyL+xBJpJbyFg2YMD/eQN3
wbaNw7yxLn+etFrAcgQZYs6dZNheS4+yaCqOqstwy8tIkcAIXJNJIVKSPCN3sZ//
9EFBGX0m7z5ftfUageOE3VuvOMSWqOw0xKDB4FzhYYR6ZPeIgAnHnaLR67CxWMMk
8x5nH1nvHIN6ICQ9etvvlfp3Jy0Hvbh5n7ch2f7OXeXms0y+TGDfacahDYm5Ky4F
SAV57Sa7w3jWUltGrLoClcvWwqJVNgznkqwQjHKLeerP614zVtegnUp3er5Om5Le
BCjGwxzT3s8sTyORWxLunYW8i3qT3nPoYeT1E7gXsfRLPhqkbANyxnkNZJ7KWw5h
AfLv9H5JxpG9kF6sdFBSBGSis2iHlk0d84AwHI7AnJc7HQBeFq/MD9LcLrRmmACG
hWRu2spgZ9Y+NTEsN4bBLCDq81t1tfJvLTTgxPu4rPjxmJR9LSoHOY9Mdn02PDzi
jgIlcy5SqMIwgBFYJXNHMZKxGRLWsiMQ98HBpy1yz3Pua7K7sdvesvxpuGx7xmvH
y9ZqH5K1Zm8lDWDtg3npQh6Jh0uyY3US2VTRevaR/WKHPPV4YduelAmmv8qn+rMK
CRZPKAgebQlVkNlMriJ0z0fwzFpyj3ZlwHintPDeG5iSBFGXz5JzTCFPJ4UvjpIe
NjCRC2rc91Gc/VLXvD9kimIO5xtsyia0tEmhDLisheJaXrZ/kKin4J2Hnm32KsN0
tPCbNEpDw28Kssz+dthIeIdOyApwFG7jTe8cn08q4YpbaiGZ+TDMFG/QZHUaOsm2
GfXOg+SVv5b0KwNaotmkLQojjY7P4Ix55co2CkuEa0JBpzNS9XezbWzoXoDfD2OO
Gbh2qFbHagG8Qk/KQTy/dRjn8ZoDWIxKnXYyXBPoPZjBfbSIsepdPi692SWiONjo
OyJU1aYcXzpmkuKTEx3t19HIjPIG4xTt/l+OgjBDE9rgbDbfSg7VssnuXSwbx5+X
6Z80ElOmSsSzTYDtjMUqh0QjIuxDQ9eLbNbGXOwyCghUWDrZnMQK35iX2Sh4DzSO
y0sshnOyBL7RtlurqhE6/vhsJCPrzmjtU6tN4Ay5J3aJ8AV0xIz30JhZEpT1pKtn
V+BbPX+jiLE78ZQk22qMnUU3J6aALS3xsA8Vus3mVhxQZKa8hElc2hSL0dldukEY
5YAEWwIDBqpD5XbBFNBjLbvNNQkSSRAwIQ3LXe3QO/tMBGSDl0/g/eJw21kr6vJU
ITXxnC0qjDQKLGbxJ8z9dg0ksh26dozXAl/XB/2opF4ao/tsvqet5fEWQ/tKjw/Y
ioMPX2ydciErNRUWLZUZPojgXOirpUsHe+F3RfBrmP6RYhgVkUY6Hwimb2uqSIuJ
GD5ds9wRjMGCJzp5ZUxeRlO/LdWDyIsT8/dDguiGbuHaPC82gS7mYyz6Qjdv1LRq
8/D4RSXG5ouqGnUwpDaq4VeFvfq9fhiSD+5AjGxYgEQpCQGx4+roGiyf3i71RiHL
wPSOZRVmquwvvlYZMHnMy+IDNfEgGRME0cOdhdbOC76bX5YRqcC/AziGdYDNw16S
EHnu/TUs4w4O29Dk0phernICFnopgURBByuWiv7XwC+2oMIAhy+LKsr2OYjQb/Kj
roQLmyxrOxJyeODu/pI80ucEd+Y34cFZKljaTXEz72ezMFlYEbjuw+0d8H8zYBHV
b+MpXGaRu267kNznAusjVp3p98zs5mCWc/6qJ/66zBwFJHCBbZjMb5riRytNGE7Z
d5XQFJnLLqblb/G2icmkyei2kqgdS9AAvxk6JPefakK8N/iy4iazP1gP8MQgRe9z
etdhS4/xF0ZMYk2NW0J5lNBXOeo7XDBLc9ri5au3k8OBGBKWR8K4lDQLF026MTT+
Ac39EPnJ6tc5onH+TGXAqRWlNCiJsQgtztEbIxA6BxMC78vx2HUXDj+h9imFuIcM
5uW8asdxXAHeChACjUbXjn3KX/QRDfYoO+c0zBgqub7Dpiz6ko6cg/0vHfJVCLmy
HmfvI0wyt72nSz8Z3tEiKBW4vyWYLhxVW1gMdlgIWOqxTupSqvHbcD9/C1s/2Lhk
WlaQcWJ9iVMt/qCcyuSXEZ9vWNsW9CBbv753KhQsEwRL2tJZXPHY7/HU01aTidmr
4gPjQ3rcFKLTcn3sfLMtkXCmoktd/GDVzi72iUJe2MyDzYt9k0NPWiUjyV3I3uT0
SY6/5Caow3bL0nw7XnJeyqA+fejyYPXrKvm7I0GIysmh1kxMZyUA85kKy2oQTGoM
s5wNmMe+Cj4vsq/MK2zdGpqAxG2o8OnsP65gaeRu4nDmM4onXfOtSLvQ7urpw+y2
fKEbORU1zdXRMtLOvkbOnhbI7d6tY3e/lP1qEt4AXu9XxxnA/JyCZTqElXvvRqia
ltVbtlB/kiM6ifFjzuPxtbXBAqdMwZWi2Y9Jma6HmK55V4s17YRq8a80gMj/WXvA
nT7093s+baNyJuLTgfrx36GOR2ibN+5QtqxL67ZuAVBzE40tNanuGTJXWjyCmaJU
P9SXYC9FdoSxVHGG1TncNQrku2hlP7GhRMTrYiNzcUG/aw+OXvtIwDYWKuy8vPjG
+jJxHwtiV3EbgAs/XJwxjshaF8MMjfe7e/j6g5m5drL9CiJTiCdhon1ybTpM0sT3
lnorkp8qcpd+jYlaDkA6DzOLylt3fD/MtvuJTi9sG2M1iegqX6T/pP+BJ6Zo8h4T
I4gilOB4y+9qkQNMfxQLHSaIkCJ74bU56B5SH6utSlDB/PMt8JphoLLKVkqbUoE5
zq4hNaFX+0gE7jL2/KNIEJ0HSFemcpx9ZcNospCS2kZqtE9dFvzvP8azlzhRkkel
65XZ2g6HJS0kUpGw4g0PV8vel9Hg8qlVVByzNgyzPv6EPOsV21CRGXSjtTat2zIP
9tZuytFkx+Ncr0w72TzcgtkKMdv7rXg+9NjVI6bZGnupN4LLycJ5BBSF1TzSkU7M
D2hiT8BudNaQ0RibWPQyEVmu3LPsbJu7OlbD0/Qpze4zB8Z6YHn6FQFNFiRcB7WE
p52cy/Ovb5l548y58OiuDmsrQuYv1MElULG+Sg15dzW7dKtBWw+Oirj4LQjRStf9
9JbyTeV/At5Ws0J1gTblHkApaIYrfO41Jj2tZgvZAD1O3tCdNJegkI4oScRnf9On
vjcqqcz33XPjnQ3MTNLy08XyqEvrpUFceQ6/UWfMXFqegXjglBs9C3jmQ4Jf+jAK
6zx3PY2bdAeNvTgM3j/dfFqvhHPYN8q35VFLDTtdAjStLs2vM1vmuD3esxkN6sTy
iBzWCd99o6b9bIQ3cPBWu/3kFFRsQVoKIxtsm1m2DXrMJtvH8tw4whH6WH+HV+D2
1r0P85lYin34Hxq4ZIBoZPJwkSfPdxkqeg532GwKlR9LEMIsgcS60W06friMWq7L
66QnvK5VPi9HahWcuOd78b8qARD4kUwKExguiJqtq0Ce45mWa0gWf0IrYSlrhnic
0jy7kJmg4MpBjGjJrs5+UeZTgjewcR13Qc17QycuHspjkRDAKm4Av5j+m51MmP/F
Lr9MkgnA/YDAMNVLNErF4ApK85IHtAtf08PGyFgVjbMND2X3INELe0ve6/lW4wIe
MiObzZ9tZzdGYVgiej/sJdv0JzB+oNRABJCfD0yxNGEcGAp8mXYGEFg7PpwnRL8h
OID1zqJO/O5Df2026PtwfGU4FekmibDGYLMGMQpfctCucpV2JebKDIUXarh6tTVb
D/edpf2jehRWNG4pOEKOr4RUzTpz2gI87Nvoh0nqxJrBC44PQyHnSmhaPMFiq1M7
OJvMMyeQhNID0aDu1MceM2IsLMc9D5nCzzmecVmM3WLC4cptBLP46bEpcdX6w509
luxqc4FRpLqd7xGvTeVqAWtPOMqj61yd0Z6OK/O7YMVzp9L5OP3mi2MP1DjWgNI7
A1lMJMl01i+TeVNLI98sYBEXT9vk2EtxYW/LUVG3MUv9kbY+r991dkc1KcIq/cCd
dA801bSnmT9TUR937SBtDBOaZUApESs/DM/ID+fWq8OJo5C2/D9+5wvs1/hRqf9T
4FLSHis1tFjK5FI8bxyY2LJPlIyjFHGJfEvkgv7a0+DhQBGcmn/RNnUxvsFJgblM
`pragma protect end_protected
