`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fk7AvQ5qD7je6E97wVAYKYAHjBRlvOnBbA8/LIhgBonpTJSbIMVfEn9l5eais5a5
agFksSJLufWMj1sLdFa7k4lzw1ALOnEiHO+OYVk22FWj7dd82LzlQPedknQRBf3I
uCas94+sukC62Ze5d3VLjnZ+jhVAqwqRTJc1uGEpx6U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7968)
Cy1qNJLXc3UZkz+uT4o40yO+RxmrerG/ZSTfsE/uZ7Pub4SWR7DBBI6g/Te8+Wy8
UpJZm1+LTJ6dEBuPmg0eSgLY309GPcZxT1W6KPc6h3COnHz0ZT7YsUfo58aG/oDf
X8swYVrexxWqbez0sGMF+jfxsn5/K0vz6kReDXym3NoK9PruEJ3N8uF/MZr7Oo35
vxpWOlhHyDjy7xysUQ8wCeI5xXTxCko/mmJkyDoAsd8ECg217oPJBlKSnVQD3qaU
FcdhtEGHSm1GZNCJ4yf9+n9FYtBnBzr5yZNKCqJ1jezItXzd5NVbVeldHT9ZfbVw
3LkQXbhJH4KY6FfW0Pj0xWgeMySxr5dhKfKiWUagCU5CCrtPKIs7QoMkXxpK8/v0
7CoYfjVxrGSzvu9zGizIcIHt8JwRH0eMpMLUwgKl//4jVBaaZVXIQ4GLtmQiADrN
nsmOiCnxHWqVlli0dww2Z1q2N37yxoRMzqACgBg2yc4jycVTDK9megfHMwnQV6G7
oCrTdqLomzUimbrdJwwnLc6MwagKqPZux6/oo62cvH/Bb29diTmjei2GaqYHhMsJ
h9IYUicXkHqUTANkCXQLUZA5k+jK2LwnKkFDCx+1/5QcuP69EuwsKT2uM0sDiE1N
J7UE0bx7NtOJRg0T51lF5tTDRl4I8P3veRYAMylTKpRLhtabEH5H6d+okZrCKgjC
S0SR8XuXLkhyHIBOoAK0PC3rCAvE3kOLDvg4m7UgFc4gQDsiZI9+8u688OEW82c/
jEp/oGWW3tNJJ3EfbBO6FOZuWJYSp6ZI3kkqywbochO/iyiTCol7CsVER9s4v6NA
Qf47/nALrExcpFBu9e3pQEONU7eP1eEvb4aOdvzf8EcAbD0BGtfGzJ51eRy9+1y5
5LcFcnt12YtQn0vqJz52ZU10XHh4EFKyVPLF8UMSzHNuzKw4DmvP6GvOmz9eTC9f
tOhLPkoBDEdyBRpiOXT2xMtAh2kRwqtdYAug7d3WJwVdJ1gH9uVqr5KC6+I14BzT
s+hahqakx6taOgkXgv7Bw+wtRqM79Ekw1WnTTxjDhIIAKOE+nvuCms+MxBbD0Np5
ttwKlpDeDhWEtFyguxDXytf52nm8QI1NSdFXC4BI8MSenShZXLbzr3EQNNtz4UNT
S188Cc0iwEjc6j6swi1b8r0+MWREkeHlvI3rPVmstN/eDOjO+DjPX0cELy3rTk0B
ciOp5L+HW8r4BfO0GaQesEaZ6By5RdM8GDiYo5sa/GniK4fvvjrNBLlA3sRPjBRP
D7g9nJZybW7A51P14WZh+PPneWEN7NmuEeUjxuoXb5O+6wWDa+4TzD3CJdftndaF
Ekuvole5qVxpcyAmU8acGDfUXk8gz0AdY8jD1eds50piLiI83w7BgmG8Z/lKw2CK
m101OSO9bo0l8wcsjDmJO7aWXY/CokGPsQl9omMex3uEhIL5PiEvMHQZ31bCsM/c
EJYcpNxnXBmviVB5zxBW+PgdlOvnly3LcsEQGhx9/rz0iOvD+MGCRUYa2QlMMg0p
eRiQHBcCwn05nG1nXb5F8Ewl3TSPdbMIxNkjD6JQProIN1J2uxA2ABUZuS7MfYs0
o/0OGCc49GQOLxpd5VvW932lyPA+2Sg3wy9WJO09hzlo7QvXAlOHQjh3JzGR5Ozx
CyGNWtX69GhKrnz/5X0OS4K5l4FGMb1XYfCvzTJHbOt0wfrVcB90l+iFGfPkccIb
YGX4Z4zHaB20CrNKAQ3BV3G/EEemZLHkq1QS7sKq3GTYD44vtBLMPiwbPl311kja
eXStWFTl1rRfNXZIrZus0tmRGtG81+CTJxBRTwLR0qVqQCXqBByX9BQFxozQUKhD
8TrSnjWyHS8NHnv964EqY/lH8l3zWO9zlOIz2XsCyzAA6JNhFrpNzQdK107xkP9D
Oy/KFdwBLwLKjSDHywHnhGVAgjBvRkfDBu281GrOwFUYqwEhqQlna/mt+DTmxSnS
RZGkgH4k0tC966FTt+2Da9Ea4Dt+B3X7pygIrQh8JyTar5FWT3neKLU4Pw6i5r50
Rj2Ef1P3XZSpMQp3Rp3ct0ua1QP6oXqEtISql6Z5p36/Xnvq3A9d2tfMNm2w2eWB
5cl5PP4EqNwkUPa1u/9ZjmZUb4XSGkmfb7/AgpCZ3XG2wJF1qkvX6TStRa3N0IO5
vmP24EOp/R1c0d8ZxLgPSKdU+mnnN4JlkdXYSVyJOAqqOHIIu2atfQi6onlW9fcY
MxMQyfo/WYg9wbzmbjwimqU3AXDSbYeq1A+GrTcGWtExsr+PocV31dGCCsfpDkgV
omTrts33Q52p+NoHhI6W4wsceHuvuRrXfwZ60zDw4zIeTmW+L37TkmQT/DTyX3ZN
7rg9+DMq9ECFrhT+j6GqysA630DB2A6Fj//bMxrolXBtJB6mykbuVA+VF6zzHK86
UegzbThGXUneyPsafUOb/PBILZbtZqdM0WOgOh7BOBAOWmEZ/yYKv2FCizjRMbVJ
Dx3roNl0wuV2D0yV+3OvxkhaOqkojrYGdS4gEMCk2XETtQnUDvGGbSBJVVlkAIJN
4RmGBlVLhZGzPMagUptff+014U6vYNnYAEGBoatd+EkqMCYmr5r7PRzKZKvZ4Zb/
7FF0t0sVaDS6vy3mUMV4RE4QPD3tFmQUHOUdLSM2FbfgizpLOGLzcOxDpwvqUsiD
vY0pmpeb9bkLI+lvD1k8o71f0QNMW0QtCetTh7t5d9H+v+YEdSeR+OQXcT2UvGqp
10ob62X7W616t5IB8GTgIEt/IBztDuiawgMl7gQlm6e5JrcltqLTihQ4w23n8Ots
2GmNgKMaDr7FMSspXuyUAJSlaxtJVBgmCyq9KZLV+8nFz4QNB34RntXe5Lr65Ib5
JiWkrjUZuMwLr0H/WcqX9Pn7hJVGjAHH7IWc4n5PrNlBjNhsu60NEqJKRkM2jG9q
jcZ27d+ufY0xaVK1lIAU0IrpY2fcCpwEzW040Jg4QGQC7sSMCPL14XN+iR+QD+nj
zyQTIQol0NK3GPLddQoWjibpvRGkapmsFgKyOgEJBuKbB3VMLdK7gTBGmoA3aHuv
qfKpyjmxJ/d8jK4CR+bc2F3edVpvYCT1a6GPSs9TmWUyRhSq4NPdAIGJM+G5e90/
+xOh+DFVs4eJWnOjbQwUm32pjNYzA3P/GVzsuB5zFipcMj/rug2fTMaUrDy3X8l/
xXhNqnPaSie1eQAcEl+7JHCab+JreFeqZSgFSxyLFL1gGzBGWvMgoj3Y9cxprXHV
/18ZFEYO17OI5HOBPSqF54f91L4AKN/FpLTtl7/PiwYhohKXjyegQ5m7xwZLxD9y
ibvfqRhr0ae7kIoGzSZazdJYtIuMWbXhLpo9FfHvSSJZi19A0nTHdwo8+/ftXprc
dagH4d0FFNdYOSOZgHpru0b2qeIZJPan8phI7Pfl8mPzn84Zwgabajm4A6s45pyY
ioqDfjWu6XR+4/NF4lugbHidfKvtA+lrZgVR696Ku3ZDnvcttTFDqElGjBBpfzvY
2jmCAFyw9FFcsV7YhL3Xei51tlcWpAu9KXlY+bf/Z8e3cUCAh6+Nv96WRcrQsj9d
UITvlKGSPwb4b9pJ5wkjgPfzx1JoaUeypMhGyqvizVStp91/Ws7Utubju4Cf7CWI
RUB9yj+JlCbsi2rxqBVrUVUnCLYVTujEq+V85Qp/dScGcK2ejomSsOvGa6NEYCSy
ZyS2bsFFsGrzMln6b9nxou/Apjv+PQH4m39QE0UPnuOSMN04Kr9GC1AgDnwqevP+
E0ZTrz+qNWu53XOdtlk+q6zAU737j+1U/1AMqcXjLZDJ7KHwxZEes0+LQDy3Ldd0
tInqHuIndSSGWCtKbp3Dlx2S4nGnX3Ar3z6IiWPPZMBBYITAlI8ZSr8oqKTsmKvK
7zrvp2q+36kX6zs0QJ6/TqeoPDrxI4Y0n8QG1hN443KHGD+s2+UEjwjgoPlmatWU
SwnxER+JOeqSSmZZdKxhT/voY/xsTUjfXD7x+ixD/6WW1ZuX0fUVtzRDQty1nKYQ
DM8KJN5bfDcqdAnywrkA3tbCor6h59CgvfX6pBn4wvMXVmp0fH1hNSzO/cto11hj
wuT1LdUxyOwl8kyl46d4/sQW+qtAZJ1OBsOnmupxzBIK+FOpGZl6SKn5fACw8KEA
C7SM9NcSbsb1+yeWjakSf95f7dUnkUFg12OHa+bUV1GdIGRoMGIh/IIVchqzGaNG
VdRl+e8JS2U0chqf/SJOKRnw6jSZUjlxyH2LWxDUMPTlwqbBpo3Fgtt4Q2shgNZ+
tCIhS84HwavxWycEKbFw0zRzjmHIHba/6UKnlWwWSkthK7ZNfADSUdRrBdmcIK3s
rtekPcfHPOK8PkYyGxS2RuqXzLdwhAgPzS32Xmst4OSF07q3MRkBHwC+sDpbtiEa
F248ejeVV5F8yzU+BkQW4NZjz2m5Y59XM2iwz836I0CuaU8ua39UO6qb0cCrWZCo
2ZDuUcg5bMAqLby7hvoP8wV5iy+sdgIwAxaG9RO/QbVQCckYlZnjATBcKrh3/LmU
IXvY0Q3FEj6N6VzcTFNgl3qoTOc+bHvD6Oa0WPHe6aZv5TovZciGcWvZtekdnToB
GLubhhk5RXp0f5X4I5q5vOHvmZct+5R/Okayc2KTg/Jesg+VUMKlGrMBESvpYFBA
reIqsmKV2okuD9HdW4kPMIXMXV4ldPa5mY8JMljK8x5lfnHfPnqYc1kNK/gX3bqy
P5BOkT2ifXEdqp0Pt7hol19d1jWAyMnhHbJdnZJz1sG7ONWJCAg9KHaoVXF5LvWj
gndGw1idYIgjYJYqNoIIBRoKqF82zRo/6Wxgqe34WpVXBEOIt6Kkw69c+bnKLBLC
vqy9nEHwiP24be+14y5yQ0Gcu81YdzHjUkFodid0+ysH61lV9VxqthksBTczPeyA
omfhU6ugY+qx0M3vu15JiNcOm0FWf7TBHfc91j1yeIFlRQPXI8YmDv239kxO9GPx
Pan4OQhiqxMRbjLISOyIHiH4QIsSAbqf5O/cPtPREhfQe2uQTS1WNIEhdFJab1B0
yiGkzut9bJ7damfPt+A8g2USFfiuKy+5CflrN4HUpw9CZjMMO2AGevGigmHvfEHc
w5oBvO0zBRwtfzi7FilqwqpuUEMfX9AQqJt0fS/r9dXQORt6ctb+CLLkxIXmZSNP
gO07deKTH8HWEsaronkQBwUeX71NYyP5OYcEN7/dfXHzsBMl0lXY4pWA7pZV3SdC
HaMcXHug3S/muIoPJrJK9muzj3br87Itdo/dXuxBm19JFSyOfkNjF7Za59lVKapX
nIrGk/PcXa/hbxOAW1lRW85osnN/M4zn4dV9aTgp/wVwDaxtabq3vUG0bXqawqDF
MTjMBRBz37idYWRj9vqLJpZZQxRYgdEroKb5vAm4x2n7irarRKq3KOpBJ2sOX0De
FdlInb74TIKzZRqK9NQIkgrKyNrqhJGu8jaMwLn9RQpLM75k4Qmlz/kLe+cZo2+O
qppfs0r2KDuPoSu9MnZAM4zQ0YiUXVPbDB5Biq0S1cRmj93fjbbKWWtosi+ObUIW
lDoZHUc2lGQtOaBw3kKr4cat0gdT49KOQSZhDnoH+FVywdHW6qT1Y47NqAMhx/6s
vXPr4f/YTzrcxEMzhxpAXRNWsUbtt7X07KpUPpmilDOvYKTZpzLh6mE+dX2x6xBv
gt3c7IHZMEAgKHEdSD3jc8NLsDKtTPGroGG1Rdjruu8IMagK2Q9IC7TKwO2Rpb4u
moOT/0Zt7l1Cz1vSnOG2n+KqmwH9a6diD9jFb3jMUO2fyVCy9NrRG6GjYJmlqnJN
Tv/+jTdw01E9unPcVyFx2XPnf4zprPwehMjzU6eVM1VpYfNJlaPGofjeJziswNlT
XAYASPgfTQk7kWoa/tTre0jEMp6Z96rbNpiTAfIKCEU5PXPb7YF3n7cZKGs3MOlH
f6ymcut4rgbpTEDOJYAa1atDP32v/QgvrRjGw0cdcXYlfuMTW38XzcMaSQ6GnsH/
GQaiDB4UStqItXklZzWbej5Lq9tHqpveGLVz1ThdIpWxSgASD7l011hZkIKFVVrg
6KBz06+ZatdLyihISfocnU3P1RIq6TI6j8uqLp/PKh0n5i72DRRuqcVAxXYmZ+Kk
PivQj7PMTcVaeXcaCgKXAhGgUiT6Fw9KRY81GKsV3Ot6PONuI+8UhtvOSIb6P21w
xHsur0RQkEE4EI9EKBSGpCxhZbGw9LBg5+BQNoIMXOMew5Ts7IrVMSn7R+bIcmFD
QBZdE6vn9MIWO7jW+SeRl4+V7P9oG/+X31CSN3sA6Lm3D9qw0TnFggOxiU6EyDbN
1ih2Q3IKjL0+rmHPpi7TkJVw8gR2Ph+M35Xa9A/ihvFupLuTRkso7pxeVVxYIjP2
n/Ie/cohWdqoUnHmn+Pkl/IMsqy/WckZ8HOqC5/DpYlreElTjQ45HInia8vu+maa
mLeMAcPHrzqVcB6PxgJ03gdS7+O/r2VrTBa9R0hnEC9OAMNSvSeHHZZF1hwO1xUw
JIVmrCTXJYwzNgQtD0m3z8UkxjUdxWV3LEoTjTNtjemXDNx6KYN5wN4DFIY66B/H
je3+5Tzsf4pliE+IuAo+3mVHmLxaVeCbc8TG3csHMj+Yrb8eizqN+nsXCNkz6lRJ
1G7QSxm9ffuiPADbZXttrOKDapncfi89BLlkHleC3dHhSS3ULysm0k9QkwKHA7OW
D0VdDeumDuWijbQ2KzzHuM33CEc/6AAWrNJkGeIif/I7ivUdcnad5cfMWI3rb74B
Y89ykpeFMOUOLJwneBRQkDBVsHkiAHdh0QuQqCkrhmknB9D6EfVAVHiQD6bvkxx4
fRrGbF7T+sqZzsLYdg8i106/PxzdIDgsshh8BbeAcvtj1upQc9eqS8zrDMDhnkyN
d1xYjdwquCf/NPKHJUc/+t8Jt5hCaTmaWSpWtVyMXfYSbeikMKGQzm4V1wRZHm7/
OJezxpHIaqCnh2aIt4mH/XSgIeLkWfL/bm/06Z1WaADYx3pOBcn9ZLz6f+FgSec+
SxmbYdvQT4ue6VCNyRn2D/QHBfbcx+ulTj3kD2cu1ES2ptRXYzoGVo3sNSDMNOaT
tuk2zeLgbEJkAHYlypB7172bybJMS7OYajckG0ghdr7OlcjLSoXP0AH7gbIoz+G9
QKFkieIWv5ljJVwFk611HKW+IfJIOjPIib6TorDNwmUzje1p2KMBU4sV/fo+MVt/
lqY/UuTaCpQ5fv98bOi0pv86xhLiBvMGLVhcGCI1Fg6wou+w/UG9QNV3/qJ0TrqJ
UeKrJMSYBcEM1MuRDJPpLN8Xn/wQDZUqUe4801yMm23je7wtUwsNZ7TRAknEsEiU
UOFxwTlUDA2J+jfFThnwrKkrSONJ7SkUH/wApwuQsvV41dl+k+RVLUtp6eJklyLP
O1/vLedTkMWRonLpmRPxPMtKTg+1ZGwTIgw/n6p7/v13BbD4N/jPpihcIP+Uevx8
CtwQjo941DfNAAnatH9d7AvqgjT7oV+NmMPQGAFnnH+HKQPwu9FgJNbTDEXd1yiV
FBufP36v2fRLWPRYM+raml1TWXZbFmBdlO3qz5Jds9YhGk/xxMH0uIDxoYJ98wJ1
k7/v303tZvxbQjuAp9Ar96G43T2BGU+jVVRLKS+my/A0sX4eX14BJzjNBhiZy/jA
PnxnGTDfbRilm3dx16Sm0VE72Gd8H1bCEyRil+HIPs6w4OQ0My83lxi5UFlB0th4
/MNBHONhg0+p2Ue2rZfmwXYLHL5iryc1BGjHgLvTLznvbmLLnGNdl1uO7OG0Yrie
b3jioLUi1m5rbiQT/Sir6wGQfdgn0MM0Oqy6/HBUtEs5nmin50R04ECGWxs/4pVz
8G+NPAxeo5VinqruoWo0VPNNsjLR5s6jdT5RTCPrLgAzfR3kBKEYb/prER6TDjRA
jUb0gwdtOFzQ7WC33r6QqFlUPEow22Hrb6+bliY9b5tCcVEzehZvJCMoc0tOnSj3
lx2QVm6VaO/Pig4wGNWQSpo8yWHCpxfIKFgKWnDKO78Gee3LgdcZr6MYdXD2k7QT
oLy2ZBc3daEJhXwiWgA0PHzzH0SI9LOBPGu+lCDHiPjhTUxZiGkQl0A1+aavEKTD
i9G9h6Cro/MsHHK6Ak3ZUgCgvW4GT/7asPxKdXvKPDoanu2YTngIMtH9OCxGCXAJ
ylQXAg2amAAuhI496sTpGRazu1dmEZnBhOwNuY4zRNtSgsu5zO/oPuBwLu9Z93DS
oQoLLS8ZX1ultBlhkvpznk0e9LQyFXI4XVjKlKD4bQBmO47e6xKFw5j96za54B0+
mad2Sfg0UzOISD98Y84eeTDXHlEru2zilgFb7BbaXWQIndK3A2SrKCkeXcdstPro
8LieBE9JdJEj/AASFc5ZQwyeAVoHc0ZbMckT0LUx38F9CgpmXQDph1PJTJYwdi22
sBsZykINtQRhYdJ0pWL6elrsdHatDv4n2xkIsvkU5K2+Q6JN9VOWSbsIIsVQ5dve
hZ7YV7ooCqZEjf0wcXUG956wMTo5CJiNFu+iC4BXu1pB5qSmYhw2KdTGlLKYQvnF
tbrYqHkmolLeUOLeCKmCnZypOVo5PP/9a8APptag7jQuGKUJYUrYQugbkVw/6C+x
Rxs2oF2+bralXwRHi+utHnCY0cLo31qzxV32w/m5J2LEHC3xjYz68lX22xCOBfsy
v4ZYdLOrQGnrfYTKQ5fEwg9XpL7CCUTCRirsrYSkYp2aahFLlxWEFYenxsJU4w37
qcW04C3+4MNzjtTnxqBKhYeLMDl+llgj0apUhMtndfYq9ugqx8OQhzJGR3mgW/yf
d6jh3UO7MceIP5IFp5gSmFWfDwA8sOUsy+YWUDL2jWDYw7zDAIVAtD+QBUNTYFQ7
zUdPEO4t+BuOS/KLgMu1+CooOXGBFpsz8YO9fw5SUoRToXwm5117405nQr2S2iMd
Ya13WM5DfZxgQyQaz0l0cpkw5BroHK43yMy2x5MHS1upn40f5fKqj83xruXRwvl0
3vbbQ/DNcZ6USwzd3aamcxGucWt7E8tiQ/btQUuabqYi2HNmptQ0O0OongtCUmUS
uoyKF8MoEfXlFs0f/YRioIOWUqE6BEXFQJM6hr+u5YRXpOLkUo3eV7UnuOohp9UJ
WTTjMC7pVF4c2pR82Emv39SiM6Ja2R6t2IMXv05WRv/QGj9SxMVK1ECoeD6m0hT2
ityZpmBnDxTtr5SHceF0Kc8Nd1AD8Wmvl5K46P23MqLDsuF0YFrbAZdBSKycquPu
kRSrKrbRtIybhK8Gm9ocpsHFlhnkN2o26z0D9Sxa6TpxQEwohKyLYnEpQ0tXPRM/
qTSVAsUDgM3g2fBu+lOcCg/JOLZ5WFI04Cv40SrF7ZlL4iIC2pP7vGiO5yAdH8iE
yazLLeH6lCxr2vsXdN4q7m75C/E1lvH6co8GboBPbf1ZyeKniGpbt14U00tNzUD1
EOyrKFzKHRhk2zDThDZYA5FCYnStJqoxrAmekWzEGTybCA6AFtVpe9NM+B+BqUFC
HKkdjvq7vn3q3P9eRpmI3E1v8+1JFiN8fXD5VMnav+zUsdtSZHsZUYkk7UnKisuI
37Qkgv/C6vE8xKBXT2JK34rohBY3vwZ/vSCWeq6lquzaHKbyXqYn7HUs6I5o0oeC
7a/GWLLy3zgq5Ql+kTX31TUm9JPDfDpfh3zD1NIQzq/ll714aj2wy5fi16yh+glk
3qoOCGMOhy5uwdHC4Kw5UiDt5M1b79+rOOOrcZTisqQxs6A/gEuCScp1cXSDms5+
bc1kL2UOuNrjU8R/Wbr98Rb/YT2LIfT6RN1DnugdqcOhnulvdYTVDwPnjYxHSMXd
CHrz27JhwFRhMx3TJbjK67lSQlfUoA83/vyS0LeQoeIoTKdI1SbADhCpr5IVEkQF
FQi9n2RqSO5JujCbV8VUoaEedMmUSPA9wQWVpGnx3tnQYRe6MtMJPzlHEE9Xb7sp
WWivfxVhDR2VmtkA21p5AlsCQOxy/i2pv6etvVZdA2Drjf+7EwzVWk95hAQ9rY4d
kqeNCnW4Xt2nyAUL9e6LstjdGckQtdSVB6BU/gwZhaUETluPLvCNXPSli6nm9P9i
MY9Aed+ZJNOPA94w4DiJzf0jkuPwisdYzkrAUynh79dwpXSeMrlh3kJadgA4NljT
QBbIzIysp9WRj9OTnBHZbz9W4YfQDyCG18053rGBWncUwvQCE0+Osv4xHKBcujPH
9SR7Pmk7g+VXb6PDP1NkH3inFNEdvJS6I4V5aMiMryhv+O0B5leNxr423N39OOis
eisRxacjP7LmGnxh8oHCdSfWV6JralHJkjyhUCOGcC8MZyUC0aZkxZwXpX+HYVmS
aDNHu0j3/qlVP89kRpR33Z+HGbe+HPetCdo4c9U0Bm0oyIJtN5zQzG1GIp9JktQr
U9NP/RPYCFyfEjSWWOFKfjpSI39wtpz6vTBz+Qc5RoggtT4jZaGQhrPb4eMaKQ4Z
cKCKFu6J42wj4E1aOuLf8pamIKfJ6BkCPGu7hQEZubZIhjvCVbDdXX8qUZceGeyg
GXCCMP+OfYqneUkTgzATls3RG3Gwe1hmF2PXNohRN3Gy8Cr7v/ePSAu+rbl4vHXg
`pragma protect end_protected
