`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Y7/56GUo723kdvkPi3mDH5LCyRgWUuh2DVVxjz7ifAJ3s8dmzdiE1yYx9mIj1XeO
OsDTv7gcX3iEbOW+W3ItaCPe96+I4O0j/EBG+PJHkHPcG4R6YPAHCgD1lLbChJ1H
Aw3w8Z+w+m/HkgW48w/z6QNclrOQl412N5c5R3JLkkE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13296)
hOM7KM8N4xgc+PztRIjU8Y4xGVJVbKUsQL6yyEOkFUrVebErTu1oSdT9BbmQhctc
vvM0ilQSgB57QWo0Psww04qTacfR+gMfb8H4jL0k1fqCxJ2cItcnge7pgNuG0DNV
GhdOSogcfPKqqaGOe7t5GtERp29lFktPmXGFwghcYtNMqnyfvyfjv7LwlsRG6ZnD
4iCVg7sA8VSnOuYW2SPexOyxwk5yFPWI7VMJ1b1k19ii90QtrNUSNpF2Y4+qTd/X
P5MPWKGOUsRt6WOyN+fzMI0ClgHSF5st0IHnmybae8jOCUI08ezO2aK9uA9gKmO2
/DvwJXNoDUIHU5cTXdEPtK0xeqSXqcS7IHtWAsj/t+j1lf+X4J0kMHWfvQGjb2mW
NfLuQH/OKTkSzjcGHDDryCgs4EuvFRyDMa/GwIIY6uhVIvJoEehavTqdUS3IWWZc
ZJSLZQsLACTVIv2O4kZvcimc+3SGCSAlMS6MvalvxiydS3UghNwxE2rKscnWWL5q
Z2PrrYJ9drfz+XwdXyLX6UZKEfYvtR6fUE3yo/zwKz/ugACJun8wz5jmax69zxoZ
XEkNUA4ViyJVbs7MiSdVFfqajAT8qeEGRlhvZfAk2I7CKr7OzlrZHp01ttaTbGjx
1skYUnXXP50ScOF0pSnG2HKNgrXNyupsP3OvUKudKDgXMQ8ZC04cGFUEE/26txl6
N3hnJ3Xkzu6V8uG8cZKT5aq6mQhbadGZicgodWHp79g9AtFm3oMI4O/WvGbGkGS3
idOIVkRdTFixpmqaOtxLckUB1V/Q2kkjt076GICJMOHZVQ+HoV005VUcP1FQfGWb
JYGCedbNXBwvOfgno52xQcPGhIoP1EnLjoCkpSdmboNNnZ+jPRiWbkOxKmwpIFW5
4/L1jyFpVHwTJEu2rA3oIwQcvT0S6TEY09066e1GM2YdyCtF0Uk+UhGTRepttDxs
r2Vb+itrr+mWRgHjhq6x44k228qMVGF+P6I81a+8pd5UxdkiIz79jKYq6Z3B/PH9
Q1z3+Q103N2u1yspc786SeZNFNgoSRm9h5bSBsJYDhv5BCfIE49jy9uVBW63TfsP
hNxxRfxqM93tHYf0XZ3H6iTLX1xPeBMpFep8KotbzkezbAbjcbocZAkRSonUi/rm
yQDpv+81rreRRyCkmzVgYyl9GKRA2x6vlcX70gG15kQyouhHFT8rO/RMak05IPmg
k8O3oZbam7FpiyC6Y3A3rnKIvDDTIHJyigBOOBA4tSMZKGxMsTXFaXRAVtT/YIU0
+GtK7E8yhqtKh5rGTsSvVA6RjoLkav3gQrJaLmjOXLCBlLkhRSXoxo6DXc+ZjK3/
3DcRWmbUhhI6I+PmxeTdI8gKk0ikp/KopoyisbNpGAatMOU4S87R/TGEhj6xYDbW
xc4dYmEVdad2QXei45zKMXz5J9UVKwY8ZQKx7VpFebgEOShc6hPS/VoLAmDE8H26
gOr1ue/mjWzgnitle/rHorsGEMB1CgSKum7b1+td5x9vx7PAiD2aUmQtjQc1AxLG
fxXwfiTJ5ry6RZ0nGxSeDJaMl7io3Ko5WUNql9VaeX4Fs64qCGmCUyYrhPYlhLL6
UTxDOIjnwbjD4DxNtIhreBJp0HDzCNh++UMfpkBN6yDGodrA1rzKLe5OVTc+0Zqx
0YZecI0DUGzgqx5RZH4qDUaZEr5a/hQ4mab4kPZmTsufBjmGb7YBHDfY4MdrrKMx
oCGTNSBm1DPwWFhdyhzeoBAKpSW0tCFqhO3LeEvOLvpS5U04i8ggH7xZpKjBsf7d
qmtYhbmQ/JPwY/9o4RhMYc9AwY8h33uPChecMYqX3rD41aOk/DybDoWCcBAs9jd0
G4TyfVuIXG3H1yw05z86fnSffherCt4pyH4+aiUFyUqyNiYwA1Z0bIGet2rJdRjr
f+c9qs6ct8xBNP670YKQRbHfNCcH1iH06ZEtK8wDJ+lVb3ATFkqwBjQuo0N2kWPy
0dRt6WUzNpduKr2cGW0yWtgeQckkyEaa8PcVjmn8B/efM0PVXh6mjPCgdqtf1Vau
O/0ySD6jo290iA0Iu+tuoLl0I/NIiO+NrvcGjWgIh+7B4Crtoa/CnA09IpyTTtZG
FLm/JrnpnGw/TWE+1Su7TXjkTN1KXSK2rh3FI2Hzl5/wYFKmcijjb16QbZ5/Phvy
1+LluKWPWrjxxayJO90y3fvGUtrQbhFpS8a7QGTqy0gshto46AZX2X97j7Q1K+iv
aw6cp3/j3ps+oKfgW6db3gCBsroHvD9Eifa3P3+g9VJGJ0GThXI4isOjNrM3LfYm
MrzqqPji3bWzC9SZ52R1SsMejOnqe6ZLgTjPssUjYpma8samcgryxwfnjpVJ/lIb
Goyv28bWkG33gjp3LyJNSpUgmVEhJyo+jr3lGnf8hx9Gh5lttcCKrZNmFYi9a5fl
VbZHzLR/2NWB7btoP+8QepDzEEOMV3qvUHbSM9i4iIAhbYgubQC9VnU9dFaOhDRU
3VtNOXxYiTekV29qxO22APQm1MHsC5FbF8tH5/OdWt8J99yfHjzmcDadGtu3ODvf
W/xDhFa7AAGODf2D4bZWunKJK7vSbDfaFo2XQRENId3/Z8qV1AA+63NSDnl/B1ZZ
xNuXBIP082tQUwFwwJdJUQz7wM//5nOv/VXLXmcvKPJO67g2Y2wNVD1w8zhK9C9h
NAQHCqLJJbHujeP7VEUaBfgqIq/QhFJe1vA5pNiu1yBvce9s0MCYdIeT8Fhe1Z/n
YM7l4mt4QznnwUafSopjGNR/NhLJTG+3NB6BYYaSS/0YXXgX0Ls/JMo0x4qtYBVh
4V+ob/dV7fpm5mXMnWeAeKjXltS4vs9rHvigCI/tHfQeWCo1XgW6FbDAtdhpVjv1
pi3QPM3m5QNDI1Y7Fo9I7lrMJKRHIkvF0mKHZyzVGMSwF1evsvBwBBnit318zIDc
43PQe3M/KtjQRli1Qm7s1in+lIdCR/knfLXT4XDfXUQKtfovCnSiSWVfU+cz4pxz
8XB6JVWHkvUagGRyeJ0AZHuCCMu2DeFvk1hRSmuRVfG2vD5OmIpopejGl1nensZY
PsF93ZuXy/U86LJWJ+hYMONuNxvIsQC3tSPJ6rxFgqx/wKwvsTmxoUuIOg5co6vb
gvLrRbMkgiS1qAUKoztigDD5uyXl840ghGUOxeHovEZJL/A0tyzzMn3oDGJyFquo
Uh2+oln5yUE+r2JPX0xGdkmzPfPRZZOO421eAJYr+P+Wnmw+5Hk29A2mSFUfSonH
QZLJEhNDuvd7nOXRQKZTo9tfLDa8bULsZrvPYmt5jvj/vVZb9vg0E5x7GeQxNaWI
9ySi6QZ11POFWdSwoDVrmW4pdNDf9OLqwtx9vlutlTrTou+SuD1WghGIzkgjVP3N
drwRsVYHGhqjbReUzCTt82URG+K61pwrp2lbw48grZ8+hRxATsip2BxfN1Hv6yLC
5nsjrIC3GSWT1EXid9E6sYx566ncYaP0/H5OjBEmF9+Z+Wye3/SlykWbJg3/TpQd
GII2wHswHI9DjevRChFuAg9Xs9WLPCVcJvfvoD33hH2o01GwV59dpV9509L50CLq
0frZ5icWylUH0CmjyQW0SXzB/45+seipi+fRAxT7Awg7akrJt/1A6k4ewD9X9pjt
v3TK2WxDxvXz/o96hrpsSNQ5YfxEA2lNuytzsxk+zJ6ayV6UtFyw+x4Fim/6RvyO
L543MMJjTcKe4ABpTUTFZZu3WvgBrsig8nwpce9JBKFR/UHvnrN55SA3ks45sZaH
tyLl7pXX3NNFBxmC+Jt0g+CVFMIorubU0jj6euvCNJSdLVE2NxNeLi2UIWoDoQyl
RbDTLHR8m+iyLYHYLhTCJGY+g4n669N7xoFxHC+RM6tMkNcvzpHnEyZUnVDSF8z4
S2R5NaXQAHJAulRVbo2qfIKSVHGwqFFpMjs4iKRr3GjIEMyM9qOe5lbNjuPNwNSd
gXEvEMC/5fmHT6nUIZ6HDRgWJRmRDisw9BXMa2OdQsswkfwqaA5q62HREds1rzok
Np9SpP1lxscmyYoQL9EBD6GyLL1OYS8InFW2O7z/2QDoyuwYIpiYNPjBlwE47rOv
sig9qLr66sONMAPR0U1lQ3wXWoGB1YAKMA1fkshI6GEqAFDKUSQDLFd0kq4oCwkm
oQdT7QVKdSQrLuf8omdQPfXKZz/A+sD3XtsWeIk3KxW+pLNBA0NCNfcFVHLx2xJ7
eIF9+XCQLoiQvqpeU5mvnXe8w89zY9AyTCSJzd12+XyYYNU4xMGQP+8upjjEABs7
oeT1+yljcjFCnJrlfdNRVw7LMN4fnI0CEbdCahKdbsOiCrPgzbVDvwVk+Ur6MI9B
OczY7eL7eiXi+vs9adCJE1zymNPerwKH+tgGdCqfmxjKVJDePm75joaV8N8M2F8V
+VtrthIWoUgkbSsu3GzwcSdoUWgb8xRE4TCU0qM6+lKgoT9oCSNSreg08D4/lk8Z
5c/L8XPBQdjAzjQaUmJrT2xzN3vridizFW1bjk6R+nRVA5jqNxJwJgHD6iohnrCl
2k6194XKy3zaBPxhfCF5qCM5tVkhpct0o2D1PjG/YYrpZaJ/Oc/XMsNk6C2DuHw4
K7xGjZINBo9waQu8PEMG0w0a4OV7MlWSIQbUdHcWNy9/0otgU22yLSzNWE6vp65J
d6O45n5Xqk4ZmHc3Uq1SRG1GTFDC8uUnltsuFa85tUXqLsEowJajfJof/pU9oCbk
Va2JkQn+fOKt1h9lC3JcVk4P8bAIyCdN47IAzfwk6M9tCyEXYp532dN3XxyefKK5
7lC54Mo04OwkFdNpT9/c7rQmtrbdjhQhpvwtLZNDDSKhjilQZQB4CUFrYV9Y6WW/
HW0sqoAyIjp1p5YDLe0Fu9i8wo5YZ8JFQ3okYgbteUIrEG+2qV6A03p4e+HkBJ5o
eAn5CR3spXm2ifY7fB2s+sBTMZDUd9+FLLGn0d/364r1rulEVfTk2YZCcbfEcQQa
xfAwikbMwReOkYt6Z+rj0xO4sJsKLdOgVqluUNU5QZCdMQWLR8nQ/hSD1juxb3sM
1lI/T6kp4SqIUwfT9UlykWn+JNk4PpHiYce/wf+g9Qqx94aIZO3u/5mWtAuML+AF
zJbyF+gUVjVLW9dSCNoYYtSNFOaiAT3OnvlTUOB9vloQWl/aQsWTiSkKYUT6fWwk
pKMxOdA4pN1G4gToRqSrpI1C+g50v0lhNrlBo3An/tY0laJ+YdL9PFop/7OXgyJV
kNxhXOyUVwVfy5uh4UacrwIBcso8DV/ElG3hQNv3jA6DwNQaU40b4OJXsp+wgDmV
66K3wf9pllq8G6n5aswzGhu6iRVLkyYLeSfKJApMg557ShlwTDeurWbVl5NqCl3B
rcYaEpCOt+iQU5AKePdp9e5jrp3pWeoJWR6q3q8IlrOQmGden9OBe2S1RUqr23aB
zZ6IQ+WctDkV6eoKL36CAU+6Gqrg1bUrlFJRxP+mWGAKuCI05d9Cdmtbu7HVp7mC
cCt25pwevzuxjMEWj0V5siVOiLtOJlPXP0VrmnsaqS4S3Kbqyv7jEwHYNbW8HH6M
oMYO3DCJfT77GRX/wLAdi+ydq6nEKN6WzPmYgS7/UImHjn7b2mIqb2RfQXuZZWuU
FaxUROdkC5saxSTAsUorvdGDDvofCDEj04DBzG5fTl12Mye/rTEYGN0EGS9pGCZv
BANYaFs5i+z4lwbHYm9j6iEfpj2/7nxk0IPoOzgp0tlxRv8R18ydUXGSA+6xLgER
wBxD0mvMjge6Ar3wQZP0fW39TiFoMvMpnXhau1uaBdbamHR6g+2VvmiXIW0oTOLT
lrCT7ryOGsxA2zNEbTyEe7gq9jEzGwb0O39+3OBwRB7qgJr1G7htkZfjJD59NO8H
GclltKgROq5zyXRPBz3UUGCukuDrp+RS0SF7vq2Ffnhfn2zuUVCw2J5EH38CjfGI
QgZQwKgxbwqbWL7KVeBeYd7NzyvsBcSqVlIkiQpNAZBZlvxuoghRL79OjAaQzOpR
TxwU/RPiFPrF5lpDWjwQY/bmQ/Ysk9r3U1pB8BI7DZ1EmdFpeC0p63SZthvhELyl
UD41y2Pmpb72iJTGWJ3SENSqQ1y2DfN6cUMsK7BfdIXhehse6R5aCRcR28caQpHk
XRIwTHHkIgB0a0WDf9moAkhnnkEPIEX8f3GSLrfk8o/4HBo53V3NiJ/rnBVMm4Hb
fArFzIaRhTWm/+eAjE0xPLEJh9xp0TtnloNaU/BJbmqWZQl1rXI8QroEATMJq/MI
xOB1FiXuEpxzrh1CCuxtUV2Ek/mCEVQOhn2Bmtr2DCXUTR+akQUCqtOkCDAODoVU
tE+DLK23X/pP4Jynb38kf1ZYEyq97dN2l1mYUJUuwDqAA13Bd2LpdzGdoB3XV8D7
/ZcFlKJinEjJqHcfjOBTpAjO37zzvid7vIoO6TsHAqlNO6uRucHTEfIeADy8KE+U
vVIoqt3+Xlc2xIAmddZ2F5hNyNneLnqDjrpEeVg5qPHt8UaO0p0ZrAAQrwAH6u7+
nNo229YhaCuSSboeIQFFtcWoMMl0+PgEEqt2FcQ+9DPRnPINgqpkmPlzyIjwXddA
l74zGk9HwWW53X3KrfG3LD2JAs5nPd1zB13qHdSqdOvOTRtiCAcF7gAxeyca5gXd
7YIE4cPosMwD0bxTc9b0h6VB+gCvI2FvEw1Y9FLwlXWIUhzfGqiwwB3rqna/y5QE
E5uzHseWTHcEpenWcyVwoVtVTDTXRjiZMFeF+Fgkgp+pTnI2GdrfVzY5V7UxbMEy
nAQfdQgBWuD4NIsfT3hOBdJsguBYH7BuxMnW6niAiHbh1xmqETAFvv7YkmjgOTZ2
BnKaDpD/ccLFkW307082BuSHy0WDUZnL5XazeODxeZkf3yINbFWUgoWus53PkUxt
+eDd1mrdqiFA/hnCssEb06DnUWmA7YupZNXv/J+nzdwD6DYHEEP/mPyZBsd6U5nf
N+XH5/kmUyS/MDcFQxgpqzx8wHTxTyEUH5zYMuZW5CNFE/v7GM3TrDQAt6CP9pbo
1A4IH0wDoRx1wZfXR23IJRk39i6yHkStFPnFoi+BqRXjyWPafkgVHavmcJ+QxZTK
kDhJW6EfI9IHdPJyI1vR89HwCIoH5fCvYrfzfavH0Ivvzt16CtINARnWcLnQk2xN
sTgyPKzFhlBkQGOnMsUHnao+3VDR2N2VgkhajM5WNdst8CKAlXmkjm52qmf6ngGI
H+vLM34xldBzF1u+FxCQ22IaDfs7tubuDZJhrhP37AOtr6kWT5aqYn3OhBdU26NK
EbO6p2KLCzX/m5jYa4U/No6Y7LX7GuzPrrOELYFzFRKhUnPqtQCVv/E9/q0K/tm/
fU5GY4Xh3wsJeqp95U67uegJ+SEGW/3x38Pxl2ai8tgeMtzI7Pa20zkU9Jumq18T
++y5ZGaFpB4sbUjXdPBBI/H17y7pCdMBLDbhrwsiOWSzz6KSzCOPEfud1p8zr81Y
TL/xoxr8VwHuAWfZY/6qmdb8SjGK/h+W9Zo6+tVhNa+SCk+QIJpjeFbWic4F3fgG
k2MT1w732RzeiQJS3pk5+a7GsqyOquxDIPnxeF8fpDqFHxIQC890S0mvViPAgI1B
GGjlyefT+2tedfSnO5N+V9YzoLCoyL1tC1GLxdfSEuohkCQunMMK/QEUdRhbEE/2
kc98Ixcs6CdvgrqqwtKuqD3nGB0d7ZoH4t1VQTz9V3B63H6IVQg+pN2iaNKVzXh3
H8igxUV8G2qKuK+jqrGThAg/TM68qgsEBhS825oj/IJHvoq0NQiM9hHPFmSOj5AA
/qv/uimlctS1DkPNcar16rcz72nAvBGmoR5MVQmcWHdsKFOEjZ7Yd/DogX5jormz
UeLcCZAU3bmOWaPZSdND+riUkOnE4BGMNOqvVwgbXgD4y5Bv/Oeq/2Mb0ZVXe3az
ISP4EtHO70+0Bw0c+hP64GPnPeTVT/rH77x0rvPX8E1DfE16LkIMimFMBRy/G6DJ
otV/jKO9ColmAHSzl9mm3i+DoQKff2DXaXhrw2osmN9+6vfc/Wk3VC6KKnSmrW/I
SsRolcwqEGAJM3jfv7fSx6B4qgEd6i0nG82CH9uILbaDbViLuVVA1OhWVnL+Obme
mA9HCUNyaO/OTe4h5jQZFLFLJAGKA7iYxWoIPi7Pf9AP5+iVgI+/CFJkEY/13re6
hLP3z1V5I+GKKXJlhuCp64gO92ME1fLshJCJrSP4RVzZTrX9AW7Iz+fPka5s8um6
j4LtLRZmTvXFwfbgBmj6X+pqA322Q0YJmFU2OKwerlETG2BxHP9yX5VekJzTHq2c
9cjCvVB/X+x2s39gljtkOKChFt0E0v6OOkxMAzOB75NB1tM/p9C04CG20FOIPFLF
qwmkLFYlXmmGXdQcZ7Tncg7IPGfQ0BMXinQxclK7mEwypU5vzE/a+b1IRJznxUHz
1ng/bh+jOrNWlTDPf8b4rgB/yY/HmGhDLZ61Mq/M3N40zHBxKgqtaFEEquuok+4P
za7Em9q4C3lQUVENPrKQk/NPStJ1wY8Jkl4JUJQNf1/kCInvlDA1SgYl7OdyDcQd
HLbwAxZi3pQKmCnjJDAeqVpfYrZiuQDh0JUjoM1AawNV3MEH7/wI61YVC+0KsO/n
lML25eOqzhWLX1TTZ2mUrzrXA3uIzhk0FevTXsy0c8EAnxzHn4iEJrwxE1yQr9++
ndOtBeiMyt3DEa/9vY5eDEn4MjWAcUx5cMwh0+ohtuLKhQgUkx5oA/9LzyUwO83w
OaKALXWHVefuOWG2ydM3Kl2DDvjr4R/h5bZUryPV62tchoUJuwtvyHRobGgfEO3k
hwARiuU0xwsClJpNOYZMV9PZHg/7tt1SU+nbutKV2hXhw0ujPbkN8R0zdH8BYze5
PmDKyzPG7OCIibFYIB9LU2aR0XtMpCkY/7d3KT/5tPPM6MnGYGJTp5iQM0JI8uqr
QqUNPeYvjvViPN2JNneMpsj3jgNZLrHv2FLcmzhKguDy9d2tQoO2KqmKETVoF+3a
wbJRQdI6QJjxU8PatOcNSrh6B7n5aEvq9MS8RSqrzYXXVsVYRanBjBSYNd4wcv0e
1+nC0xkWnZRNNb+nFC2A4WfsS5JX110DkPOSvcldnA6RYOunbShj9c2JnH7gqGLH
SRspNB7czfhPX3Jfi6xKWvYJ84FeprBMjHMVi6NGw8q5kM8AWQG2xb/bBvZo02Db
GoVv76VgKmt/ClWQtUO8h49cpYpjiq2hUkDvgbQBOt04jZa/SJYCuNAOODfixBZv
GxT0hoTU7+BAg/TYR7itmhkgVyRlUSMjxquIFbPXlahmmlnlUQ4H5A2tBQfl9Fdx
h8+W8KHbvvGjsuZPF3JaqdEv84/ASpg59o3VQ8jZSG/txO7GB84HWZ8vz099b8ti
Wea9IoftzKBlH4pHOBvhEorh4WCLUl83WmicHaiyZZsXXrwZDdWN6VmmpaAc8b78
WQLn7FN6yCAOBpRDjSlgC7PtwLqIfqEacsfe8Hwg2avNIAqO0vxmQgKHmozRzdLe
Qsl2uIB8jncGpaHF1f285pEZgcWaCkiKcD2P8zSEmDb1+Xcv+3SudzV1fQUhWx6i
Ig53oEhtqBw6xt6JhbYEE/ogqLXuGLr0Pt7x4I2fe3xlbBJADtkGhIgzuXTFV9EN
aTZlCYPEAc9PQsKGjbI6oq/EinzM2r3C4YVKtiAPya1RH/b8csoT95n0RZGguHV+
Kuj1T2EVUMXeNhMRejxX9WqSfEkI4RV/Tohr6KT4TjhJPD/bWodNjQvP9AbwR7Uv
VxtYk5zsCZWLWWF+t1ZUR25QB54mqlxGKUBlWo06/qHfxfSxtv4Q635YHEuI64fJ
Bp87G/GsyYUgu+TrO4dtZwjeUL3B/lprFmXOgU9Y061d3eTTi0THwMCGTbSoTQ+O
FhmQE9frEKNU6+ufYrtRHklFtOw6ZRJvxdbWTzzOHkNM1HiApdWn1o0FDIQF1q/X
lrZc6/cs8IL4b3V06Qy+vsy7r4ugyod0CM+BIZAIf+CykpVCeiKCfGeOAKqrqBw0
4Goqh7elTIDc5UepFLQhbYdsAfJJijQzSm1G9BVFV1/TNg8mkX0X4xIrRis/r+jy
8AqvKAmKGdfZlOtCfhHDLXWu3B05zy+nB8GCYy6Aca2ISCF/Drgy7iYlakqdVf1a
plL+4yOoRJ3iAbTgl4SOwu+2NuMOPWunzUhujrWQpmd+jfaRDAfvyXrDl6tfhA/d
6y/Ipsm1u54ES2YM0y9cnMOXAc2xBbbU3leWOtopLGy0buQs9BgnEfKJSTahZdWY
ugxxgvTjQ44S1uM4AVgrWAdbnFe/9UwTlEoKxmf84bN+FfkkU/jxingE/wA5Kf0s
7KmWZkxFyeZIs/nLBVVpPoCpSv4USz6A7SPtFUkY2FH/kR4mfeHvKNyDANX67uLr
n5dzpZUg2R+Ky5EXWZMuMuZ3ZtPNj+dVG8/3gdwCO0uXk0wHT+XsOJbxQ2a2/xs4
9ajcF7P4PO29osqaFHoupidD8Mf1Entc2etOEZQTOKW9EfBBfrWJhv0XwpQDgcJg
Jhs85I5qM1kHzZX5aQGhxTtLsBz67SjNnhQBKZYiR+0G/WdXstyhszqypbEUYh7q
xk0hbHpHgvp3SJk3ygd+vcRpjSMRa9J/16DB6xkrZp5WE/KYud2lYzB60zKFb54b
AYH47d01VpmHSxhJjCJVQZMU8JCY3ymwEWLofn261Zd2MYFkj+6IJywpkhVH3iY0
WUhX/G4cDzyy3BSsew95glYB4MfVSvCGkkAoyVPPawJLVlMw99McC3M/XdgxFywn
ow0JCxNNifmDbymJLVl4FvsKdBg2rgVqK7BAGK55LTWHRvh/SSHazSB+YD6RrAkS
CqORr66ra3KCZy9Z77zrc6LJlJlv4I3hfipteG1iOS09M2TZK9Mh9gslj0MU7IgY
WdTzJ6JObSSvbu1BMZMG4C3zG7IjlGOimY4RCanKXO/Q43MGeYW+FfYsQ/5RaLDy
Z4s/ZtJEsmXl7ldkAr7u76XmhCj2R1OT58wRB3bEm2Ta73b66dgGwzk7cL8Jbzp9
VA1Z+9LRh90zBduJx/VQDIi98GIblncKULbLLpwYpx4rpQM6yaG6QvsPRfoN4PsO
9DyZ7GkEbD4SVZCswET4xkKZHLVs2CGRZFBnh9whH5HbFH3zOrsw2HwwkYsgxe0o
5CR7R9AC5Jh0AEnBpK8S2eqz9+sLF+DgSsGBbDFMFG4Ez+pPUU13cTZt/McyVyh8
FTG9XCi4UbbeFrPqDlyjCUpP63Q5Q01CbSN+ScCKNFnDdqLDKJO2L6+SG0qjKrVN
H1vQ6eyd6yIYCT4E7ADle0P/r4jblziTwvGaRMbWH/66wkVAaWQ8Ya6UvRmxnpKX
Z1GuXbjMIyyTGyAjLOEUeUxbJBTp40ySDUHvj+h1HzfPQrZP6uhiPy+dJTH+E3tv
X7Vv/Fc9CO1XJTeEselxzQt+y3GkxiUa+WZQPoLEYYAGvcwEu3fHCpA/SWBm//zM
3K7bOx8GqA4LJmuyjJJcF0UM0Wfrpv/vdhpQ79kjncBqwSRcDeO+j9nXiUWBF/0J
G9BRgUjA3DCl52tTDJzRSIhKO6p4vahdk4K5SbRE2vj4tTZf9TzK9E/cFd9N1jl7
VRmk/D8rAVAJFGbwEGsz9ofcLAM3iSb7Zv8S+lS3fGqLu4ccHMX1ejyYH/MOti+0
3EBkJlBm7LM3ygOlyhm69lqDGSFC2RwWUxDM3R8ophtvu3JgpDx/MSfJwtBOMAgW
Y6RT/6B774dgMPa1U/RCjWzhryPH9NwcyZ2y3iNElH3YFjgLDX/6NuqAHsQ4iddd
kYSFCJ3bRJZM8FMRkMILc98uEGr0fUHX0YNUji/L4G9hkrhfmA5oNdS8I7F7dso0
JiYvHVMh52STYrupckzbTT4Q/C3qjEVotq2Ggeq3yp9gH4Ojwtp3aFjibGzQcEC1
jvzsj9aoCJh/xogweOGlzSR9V8KVeqNgvdzRFJjtvLiPWl/NIONj4Lebk6Z1kEaq
ZPHbKBzKa5F2O2O5sMEl1ENEg+lYtjW+dxLG06948W31dqoSbiG4ckn8eDq/OnCf
4wZIXTdMh0TuqsQOj+8cb11WMjxRaQ/KexsSlxuVbh/6EC2qP+vEETPxAJOvJ6To
M+7Omd6MshH3Vr1Qu8rAgmufAv4HLCYU5p9cQE0+AlcDORLaXiMu+UYp3hj+CKK0
IpNZL1MxgTwf1hcUvFtCzLwbNsuDxhW85XvyXkoQXLMq9Sjqd+BFmeEsbmz8L0GK
oqvYDmQEQ4M/q8cwnlZ4/3FAyFzOp8t8Xsf7vKjVmhwRZkoUaqQqjpjO4zTh3RiS
+Ct0FqoAmq8x9YM55guaTHGoHuYRT89aCnuDnyhRK6jZOD6Qm+xOhXZXdpLZGn8M
gMMtbAMTRhzP4WaX/k9HwVQXKEe95h2qRf6WN3hSCrizxdXrr6ytRsmVOEkX/bAu
lXxbxZERenl7qQSfRksILsIoFvSm+WfwwDfdawx1FKCTHwW5+uaCs6dcGI8vKn5w
+R8U1B8bAOf5tCGfTwSbzULKMTdiIOM1dBLgU85jEVdT9d0GkxmC79pKjsMdiWSM
KH9wVvsMqj3NcYjs19A65EOAOenALmf6VfcMfmedjLYGmGqbPPGG51w9LfinLc5Q
CZxUzvAlUrZvBiFMfAF/US4IcPva5tNkLcjHDbcWX1dODUNnd+EtYs+TVTYy+AGz
T7KU5ASaBNxBfC6mKOoUrNUrKl7ejVI8MbBvIAcZxgfl9nfU/3mJJ5hMubhCzT7E
KoncTychAWBlvOxawuEpsR0kVsIdIuaxCAvpy590VOadSUt/Ul5UEP6VQrCwfNsE
wuAtYaasqYoDG1KWpN0q1HPCvCcj+cAj7F4JDyj8mZk1sAbJNg1ML7NHTjCNutfh
UnzDUCZekH54W+0wIN3ozjNWfgw86nJ7SB41APd8KCDhs8b8fmEcahyjAD4CON0P
hkJLI4yEXsea3kIzMsD7pGy1nXayQKYCKCnncdkXFzG6TSpveVL7rCKEAjZlKQdY
eOBMkoYTc2ZVDe17fCvZ/8oYXEI41F3SfMS6lJ82NmXESWZ/c97jHjNPa4GNmLQz
GCAMrsbvHUcHY5yLrDzCWY69Mi1KqaWGQElfXByNhXVbVe/d03aH2lBYkV0M4MnK
59odyXuwuTIwqCskZ/CcwFj5rd82/LpvyrLGjkKb6lEn4CAmRBunebahF6N+8vAS
i413fiAC2BdPGXO/Fo5XiIYtZ9vNYDmmw1ijUenAegszU5Oc4ykJdmTHDTIz02eI
lK5TaEB5h2rIzvP1Js3M4E6qbkltl1fOfD1q1ml6vH6TibJ5FbEdXUSU7VKwRAgP
SvlQ101SDiSAHusEmzCwOSJ1o5PTsiTUdfhzhOJr4OVktK4zXwdAGlerN0B5mAwW
3TV+zaGqXXmyvy/GF7a7O1S01Uh9RNjARRvq+bvsQn9f2uE/d2z2ZPkclHfmRxuL
ExH/H6/UprBZJBYoKq6nJxKlqlYdo6/oCDuvXMdy33qiPf+NJT9EjsUkopVCgvfd
OE5btCVMDODKRx5fegyjVeQG138xU2of91c16gn4Mr09/r3wl2GUYGSfRgDZ2aHm
H6jno0LSI/vpXaLj3i1Gb+gQsPWqOflRPy3O5KUkMFVDq+9UUV90+NAH9SWL2ET2
NtUOFMBBtig36xsKlvhPZYw6JewhhSmFfhEJmidCua664Tn9krCsjRlWNlxGaQRd
C0NRRUVl2N1+cox50jAYNE9olrYQxJo1LWxSdICXqFbPdzwtQuZZMhIfLMnYPoVf
crSXo1yl4LsXNl3HeS35wr6+um2bwwsJr7JB6WCZB6nEuOgS2N5pxsyQNcW1BwYc
Puaw+HAkTUmdqxrx9QebyiQz7m0D7QAyGQ5K9gAuxaLPVkAii3TcHdX/y4yxVYpZ
b7BA+TtIeB3+nFJwTFRyjnvEWk59aPbnJBzAGySJeBENb+/CfVzsvUUETqAUGzjH
6S7qxhC9sGFGD3USIgwU0/WwsvnO97a9ClxNmXM07d1YNQy9D8FBgD4HIHXjJ1oT
W4bq9Xg92orOAmqmkPBf1VxGE1bDvrVkCcykaSqBDPTsVye4YpNUBZXuFqVxodkb
95hbRWAbbUrOOXR81HvPMwHgv7IsHg9hLausARYegEYUcYZJvzkWOmjX1BBou6jW
q3rKVhHljUAfgn+YjTJgqFOnDc7kFlZ8lN+8hgSeZiuknC1rbLhEf6JrQi7fhc8g
9rrccsJpDh3jgYusL73970M89brxbo0241tbW/FE0ZTwyS8aB5sEHVyRBVn61MDq
bQzlVmvVyOMUaCVTQ5qf4VNfNdbv3e0weZ2bqNRI0M3LhjOhcrXdRKHroLeSFdf8
h9uL0tMXGIpd1377OPJCva3RW7fnThzK9kEnBXxPn+I0oeg/Xh2HKs1Mymq45q1m
rz4cIM9L3nO1LrGoAAX528oLTDP+LsSuKUW4MbOFB0t5De32KgJuQy0by+Uxtm2K
DKIe+esC6x3lNhlpjFwh/QvxIC8ZWmjlcczI+YrcwFxrtat87t/7vKJylJZkMgON
PgSi9Vs6we4q/oHUDKixajAIkinJ1mPLab8+5nxo1QpegeyU3VOSs4dDxkokLwpj
I4/JSWoupB3beyR3pnAFWMzYHSwLsu5oeFK7i4ifTn+Js6FjNSnVJsCycrDfIYK2
OuC1BinEmpVh/xQ2KseehzTT//JvTTeB/9BoM1TeUvFLF0xZN6bMMIYtr8vMdGM2
57T80hFKOPI0CXJCPb3p6FqgfcDPZ0KM0tsE/XxUUM9V5nnk38iNqcaYfjFnCR/J
8KNYbI20XqE7K+v86ph2NSpG7IcHyoofeMO/K0jsSp2tmWL7HhAPzHk5uwVObNU7
TYhqpD3vXZNqk/NJpGcSjVmDFR7AdK+mB/cIOYt8+AXlHLpInzvSqdgt4peeB2de
0FdxPK3EDnufc9LIRJlKdBSHUQfREe9Alr8h6qcwerjEko82KM5Fo+kc0m9ri1kM
gqQlhKkM6mw4EUGJitVmWJVaoGQuHS9HlU8OctNSka2R3XQOVcHSKtBGbBDM/s/2
4kz/cvY9stq73VwVFay8UNUznuF/+zkUP59EfdSVXs+L5iP/eXpf/PJkLfFo3Lx1
1iNM09Bwlvf4FKIQLoM22dNTG8Pvd6kvlE7/p2HQMoaBmpkS0fLhyq++Gub+Ipvi
iyCn+O7BOugi6I66QRWI7SFn4tiFBPnu446pWP6OIKwG8NE1STDgIRaxqg911fm7
IZA02dobTdnJvh2qtg6DMtOasXmoc0YChcXptJmXHSNfpvBFahvvwA6VIE5DWCLl
7pzos0cMI0dCEbSfVLuZgi2vCQr3Cim9ERGR1hRdn1zAG/QGYz0U7e7AGy2EVaGa
SxigKLZvvMZ0FSLe2H3TbJjNUi8sgq74OkSaTuatcJjdFpprVtHgAzxpSpUICg2f
xN3WeRR1BshRe277FUQtWTz0g7mzw+DLMOblBlQuEYJ9FTZdia0nasl33AbrGNkO
d5W3SKqSjllK5VYa0Ojj6oK2jy2lDQTHyW2ha4s+jPGQP1+kbCimwl5FhgAqYuSA
OgXStyodHbSd0Uz4eU0R7xnbHtF6V8MZx8xgAH7bbM8DawhXr/YhEodwGT1c2wYI
nRzXEcSKJUP7fkUrgycng4aIDDHhcWLgbLupNIDZxqi6zEkLIaUk3V52I97rw3on
OnHnQHb6aSgN4WWTdyCwC14VZOHbg79hE1qNHFLrg77u+Fk4SEgZnRv3lhDrCHNW
/vKLouhFLLXn9KlKHNGjPvd6DnQLb1moBboTYYcEVRgBeTYgL+P0lxeKdusavf0O
m7Bg5F8CSUuo8p3whHvEl5KIxrCoOLMAJx2RNH16UrmozRI+yd8hzeT94J1ezaSh
eMK0ftEK5oGQcgKmszDJXmg2Bxe4Owb/p28ULhvd+cZdbuWWBil6vO1GGbU77ZvZ
LBeVio/4q4DcquVshQvBe8DWQIAr0BgybZdxbxBwBzm1hNCqK/XKSBByzenyMdBp
+IyHMo0619ULG9efpYU0RRUpOKo430+f94aqIf6cwfyD/ygVqdh5qJcEmj1IfHdK
GuR/QwYSjXnb8FhNi/TUqzm3OEis/Jj9PgJNY8f5ve49fOLace/UF1tXqsWao+jf
XbfWqq9JVJ5LlN+KRbSfXAeQY6r4lGTMQdxO6K3CqhQqoFlRim2mr1vUFq7gqlfU
AVc+zNJy6NJuHHPRsTkrlXlXVC/A4PnuJ3NV6nST4Haz+4T+xuqoLPaUxJE4Chdj
wbT2TirDejC2vXx4TKcNMNuIccZPEX1j0GipchjNErBCx4bv8HnlQyQCUk4p+kLK
I2X487YkRI2V+GXQRZwhG8RTxvWeNz+WMGJpAJxt8O02kRCqYOV7HSjMHjar12V5
QfBJI3CmJR+vBDb1FBFAx151QC7A1emIom3cTCGHWreHZY8Zcc7ZoPF7aLF+5Frk
TNOcKAGYJeAr5r5pWXmSIDbJF18i/PpP+Ffw17jbbqI5Dwxwki+Zwrt+7XfAovjL
dd+xKyHtC6zk4HTI0Dm7127qz1khWVoPaWrAqtyDPjWZX3kOC7WAjr5/iDVCvnkS
hZ0ayWCF4oepBTM2aYR+GmKy5G/d4iJuLcXMJNKPmrWf3gOvo7Pw2uwL/DbVayIN
m7/DmSeJiiyShOOvlzezU4umWy2ox9jVBu1fcRtTFWiN5LlblHFQlQlnk71WB9Z8
1gBLj7KZpls3mW+k+szSgE7cT1vldDqbmz1ODpE9IHL7mp8nNieVPucN3mZb2udL
sUMBzcrjryCmSCHJuTmASAPhkYLb8H9H3rujK6WutB8otpt5EGK93A+7bxWMplkZ
ubfZaO49hMOiWgXScs2+baA74PxxvPcmjmK7OLQAH0Jhex0zNvcM2H6NkenhjLAC
e5vV50DGixD1k4ZcHHM/cOSOHtxa6GRXfvMTBTph6kJA5npr4RuQ9zB07dYY8zOK
zTlIecCVIvnAr1Y8lr+Io0s+22ERREiEVFw5aE2FJsIGTQze2Q4bMb22A5+fFa1g
0HN96a3Xe84V98BRVzqkZiAGfFlLepjkP5E4fp9tMLsC8sy6sbXpVKvuudHy9Orz
gpNneFbuL57Jcbkw1cpZ+uibYgNYIxHLzqv+WuNWqMqpiUu2TcGSI4xpWY+zsbOS
bkZnpwFRyWrIjgc53nbawpzPdKERMOkU2Ls7OjghhUk9RFS6nZ4CtIXdMaqhoinu
BvbVQ89JtMrXPvpGO2sOGY8Nyk7VZsTFflIA8x1ulvJnG3uVvOOpwKOhcLZ3olia
/11ZjcStFpMJA8zi0j0946Nk6mdCogK84EEXw3HQoPzYgyW6j9+XGI+r7vqizfXi
S1B8kbDBvTKEaXS+5JODnUpg4xPTAOrt7JmHK7gASyt02N36Ajup6eMfNs0HxzE5
GYJtyPbN15EqHhzWvrIYENSqyfUJjiKlvVje5vHblzzpcErVFS7iDtBUWrxRQRNA
6o+exkPmB/hchAJzNBfrXuMrwYl7EY+LUfpMK2bHxwyPwPA7GzarraSce+8iLUzw
l2n5k9Vk8w3JqF21sOnf+1hDMgmghMXG9oIFsX/+Y/ebXFm+eZGBDAdwerAMUrMP
IXYj69Y1etm/GrWHjB3ka9KEnW1TkgLGFlv1rXUeJrb3uNfLwx69vMnTtZQ36bzx
`pragma protect end_protected
