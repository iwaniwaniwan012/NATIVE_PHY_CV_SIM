`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XSWuWPzM/qAh+HPlKd1tk4n5npCnDRabTyoI7hNvQrjX3AvzrpRPoL68BElFPXT/
sV/WSftHgyiYEmHxdnL5ULeywcgsDRs4zbZ49gampIzfvWVt8ZqR2W6TlctJqy49
ebS6Bsr3WtX3QE17M+WJ5R7Yy1TmsAUp0RZM7E4+vJ0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19328)
fIZxvBDPsiWNeLXbVlNhG4REgDgr+3TCLjglnmmb1WSOnUP+x285abYSededz1ix
hIerAxC8Iv0etOQ3qJuwe1uTvk5w9yeEdNoimeFNzNZFaTXJ3XUcw2GmU/QvVKC2
qKM3R/Zu++vEpFdHyQw6uhLiPw7wjULze1M40zegcl23og5nX9esccwIwqk2DtNQ
M0dp8XejdaUYnwn5FCo/Dpoug7y9WJKCrU6k9AMABwcdeGyFJomQATgvg7DKmsx8
FrzLQm1XjmDUdM5anHVBkn17N+27l5asg6+FVK0iI6OamlKaSQRcFyTed3RgzV0H
pWisgGphvrlSOiUpwrh2sgGWWh8nOR05uo2tHn7eNwoF1twiaw2DeZQt7uGuAod4
LTnYHCNZgZjyX6zO7FZguNKmdRUZvUK2I8Y8rXEBzFGiRnvpk7a0gPjKG9s0q8dW
ZTL7qeE75sJrjrwxg3plc9qe60Mot6PNlKMVitekbv4iDnVl5VSbvx1PSLVIl32d
c7/QjVsCpTfLjcJf9gbVBAnGtSbnLWw49xVZSFxKD2+ZgOYJACl8M/AbeMV2q/oE
BernjA15N4vVAVrdTh7kFAaVG4OdODBz77CjuchNubF31zykk5AFeo0Vv/vj0XAF
CDULgON9jLWKV2c8JpIQ57hcAJWfoH0bM4khSyk+EcSKv44S+XbpeM7zSd4fWMdQ
CFxziyvWJ066g8vQRUw9H8vtPnKvy2ZQIknWXOTDCclA43OGklvPeuHTcAks4dRe
yhhK6EqyQrY+XVA9VBlidWiwtQnpeJeh6+LaY6c4Uk4lsRMG5npeFaLy4KpteZ08
HEqg+xXEvl+a9zPPZIwR+b5yhQo5z/xbK1tHWLHkgdfN/vqa8c890Ep7aRx/AzUg
+sSxZZra5NKr9/aQrhfZL/2l92AJnz2JOYKMElOFT+peObX0/clFAVhbnGPvdUQ+
svcSA0KiJfhKi4ywFaqx4YzMa6dqtRHnXd6a2iW1MFct3u4mwfZaEGDiXSfqNwVe
4eHJCmli8Zk0ZCwiiaMdbC3eO1WMhK13NBjIQPDcMDP42ZB1DfVrGyshvW2xZg/H
2NrxVFmBTfByc5PyVgLB/MjunFWeY+5X6INyCCypz8bJO8OT3nTqGRqLd/tJUx0R
lv++pn0vDCLDX1DDFJWtiHQplo52l3OfETvNlzH97mtxrXXdUfXs3vGv+3W/h/Yj
htUvfjv0qJsXtBLkQgI9iFaJQX5ZAz7bNFtjLTYigLdu99mpuVMWqh7bNB969+vb
aUHnPPaC3vWHRKISQjCFEIIJCGKVfk5hNHvgDbAPTCy4ooNTM/sJezp3okgcS+Ug
G71gB0kjnwpxusp5nuun3VC/mdWlybNyuixVb3m6Q3gBVbuVRJACdr4jQy+WZxtp
RGgl8zShtWnnR3fRD2DoUaIpFg2W3xaEIRsZj/qzFyiM2HJfcDFhozC+MMJuR/do
MBSAcO9UW1UJyJZVMnPsk6BbHLEntOmf1UGn052KWoOVQiEqmKe7prTBhxgFVbFG
tZW9tX1ydWlfZ4Rh3kJP6zkD7TT5G+klcPiKaot6U1CBQy8peMjpczOLJVLj8Aoq
45yC0A0rEt0zEvyaLlhr+E3IAQqPqVbJ2ZBmO6/sE0P89lDnKo1Q84G/afS+J621
b68Gx7Cw9GjbDplWAK7P5u7yupYX/DyAHIKG+Czlk2tUtTW4PMgDm5NCYg3IiTSH
PAOo+kUlZOfjs8oIZ3JBxXxJ+C28ig54y/EHsATLD/BgQWRqXpzf03PWNcL8YXcs
BPJJbPAwsKQcsmF8tKKrFUhRRPt4GNzpHDm/upyljjTU9DCBq3XhtvLDFWB+uDV+
DI5aL221sHlyOkbkyAuV/Hdafhg9CN+1f7ixveBJDfBvwGjbGkf3Sh5eEfDXkol4
tIkziN9lwGoS5cd7U1E17+YFdaiS/lXuy4Z1ItPIWQjzI0S/mgJW0gCtji87drZb
vgojW9q4gub3aSqRNqakUbNJ6T8/bahc9j8GrD3K6wQ+ydczaaOWIhOWQ9v3y3rS
mlcYeosxU83DEZ2bNIVEUGzukFx6A4kiODWZVUw5HA7DBjjH5xJXWIELq8M5JzIk
F1ZusYfk5KR64tpKdS7wJS1K9t23piZ5LlCyTi/N6NWi4HzLbtONmDuwQCYoISUB
+51+Ul3H/0PAsWmk1DR2zKz6web8z7aYoM30wWIYH2LVPjAZgDGyEftG59tVk9MM
JIREW0nE3xCbSG3ISWnSBsCGK/KOUKvzvYBmZAfvA+jGfAgkvkj/cb92CHG9CCkQ
RIf7FoddTJjWvb+pXpsP3r9RAhNYHvi5BE8fauzuwUtZ4G3utA8iTPsyCg0QFDud
G2pc3JBMBH4XmTxF03kd6r8Rs8zvMI/6RwaSxOBqGo+5bhE1x4dQwBO6VxCKZLUG
s2b4OW7+UBJ9hx8ZC9GP74cAeO25xHVJDUq4VpbijofpGWph9dU4652yedQN7Du9
hdW3YOTBm/Jbe5O28G6boLxuufciHyi2v2R0RfCwLv9xxtiOkFr7nL5toQqSETKT
/CkbFwSvvn5o19A8zqzxlCmBHV7mJwwA1JeGKX3VH5xk9nXZeiJX6FhZBcaQGDlT
okRN7Gbb3YSXQyTTvtugBzW56FA7lglMNxzNKHEVbeUEJAJwjwM3+vCE2qEBXpvm
9Fd93vdPGhE0PE720A3Jd0+6BOZa05/iqIyOddn/8djU2+BS3Mqkwg2CEoIKCJOO
Bp4nGuQFE1xbuTg7bYncMGYa3gszNdNOIDOlgrolPvgp+kjY24EdbegjSkWSNNPf
SCIep04qoCGu43/GOmo/YvNxAds9qs6wzrrtG+aOrayFUB6tJxdr+WENlCdcD2iY
0OFgHV9GSymVeH4RoIOvfLarH5DcfvOOuFsia8U+NolbhHjdfLnsm8tdgJLDj1c8
MwWEs+H0xJrIYaXFNM7kDjRp+OCBnqqG6VoqTpE4FwTaPM/C07cukaLpe0rmn0PF
9sYze31ON/RK12BPhDNiP7PrwuPEHRGvXGE4HiBqtrl9DavcuBD62zAMCi6t5Wag
5zS7dVuyAkuYzZErKQpLOnxJXP3S7m/iD8gBhheKgJCnul6Hlh7tSyanHViPVV6t
0CuZI51ZtQZcF5yhpyIc/ncmS9IWex5HCYDasJFVb0fxOBzMDFZYyOpkT3yxQUUI
YiWZAOOoFpkF5+KPtKh5r3B+N6QglvxYPnGoEwwI5Q5eKYlDIxp3gVZ9a1JOyGDb
qlxuuEn14NYOUbX0Lmv5Kq1M6dzZh7jKBq0tZsPLLbI6+rS4mFMy/9esy0aBwOX0
jFa3q2cR38n+ZwBxd12B1Q0j+TwIot7ijsIRqA6d+bspVeEo8BdXNzilGunOLGqZ
m4d9tmGY75LF+bXmyhpRgFcq2RJ6RcgkNaBpBfo9+V8Bv7Ymyi5ZUKHs4knoLPAr
fbDFz3q3ilTAoJQ8Ta8WqL30FfM7sANC55I0fyrwLDIX/D4Umh4GdWMouebNOsLl
2mI0bVizjskcWTq/PUeytN7ZVceeC6nrr7t8uruHZtA/n0wDQcBe5J71ccjweeoU
aQV/N1VGSlsfK3qo236EVKCpFOEJFsR3RNJC8A4ge6Mi4DsgNiuRML/rjDqNR5d2
wgnaNRYQOv4+pqIMP8DjszRhAZVjcFoF8Fgak+63IGrJ+QfOQU9ckiVWiYuZpkMj
tv0R3zGeL3n+6Ix/FNADlrHzUJ6lR88e10TWTRlcmru6V0Kj+/4dyQ01INk5YLk/
uag93CG+/8svF8kni0ret5bl88jgT08FOd3DTtSto9bTH+69eNYbFMmVjV5a4CIT
Bo+UD/FSbIqTmWfugegfP/IzR2WWEADvJhSXrjxe1IxX/ZeRxiTlUJHkk25Sb+wO
d056DB8hkS+kpcQK2t3LO3jvUNtmeGkq3lVcSxLxqA6WhflpOC2dq6amy99h/WDX
RDXdoQ96XQmJa8pPUZPwAv7NL3ftoamVdf5BWiEs2AawjOCF33fWvdUFTuzC6K6A
rm3WjoSw9CbceKZG4ONMObAZkE1XqNqz8GYygeSvR1rXVf3XI3yg+g8wLhizOX3o
NgucW6+A8hZxw3hvt7V9/R8AvwuKXS6WhFdF+II7wN1y/3IZ8rqHGr/LTpSm+pbT
2FKt52xr7P4DDZLeILa6CLZa8OR6jx4EwvVVH4DbQtE4KPMWgVKGA9KpGlZi2gkB
OqFJNAFfWba3AOmF07B7oNi3XdLyw8+5IkkMBubfe4acR8rr4LVRqwkcbR7LANG7
mmefBw6I1/2Bmpg8qmbWcJzOfTrKCHFCfPI9+9tHqZibaBtIOmOCttXtPsXVT6Sj
EQ+Y15dgCMnsq5Mcdl6N2gRnYcS5d4Ci0TKTR1bJ168RR6oeN+Oim1k46uUH2hOM
sGRcuR0h7L3c5bJI4HJhXGcl2rHS3bDU4bO8kcd8L4GVbcmmmKZuy9jsvR2PPjgj
XynD00bfIRxO9aGA/1ltiNeQqKMB60ynEff0IvkV34xqAp1wEPUd++vSabxwZDG5
YACvLY0nsZLs8+Uemg/KbXxen+ThUx55wLSuAjTbNfSTVIOLgoi5jwbXu3n+81lG
IzXFbRkwfYVkFJx11BbUsfYuOQadV1Ch6LTbhj7w4fhffMJcSxCErTDp66uCOCdP
yqXm3rylkcg7oLL9SwthM55Vz6Qo/J5FLQHwo/JU2iXIugeG+DYYgXzIBH3nEjUo
eV137At0mNBDR2g7DRiE+DyZwk443wHzN1xf10q92SXeBuFq5rYPt9ZKU5dBub45
sydmpWNLP/KeIuI9CnVlRnYWtu8et0RuPvVRQzKEaattPxj5rcmHlE3PM0MnQLHx
gcBMP+iuS+HPFs+AukvyT8AeWTTIWubvJL21mvPqWAzDf2XzlJuf3emFR4nSHtsy
lE20/zMLg7RTfm0qCv7/5G1xFqiZWRp2lymHnNJZ60loVYFb6f1mkoLNK0gPBhLs
wqUoYyIQlkGVRgabxjP1WmXFWdC1H3vP1NsjBoNuKRw8/RnOYTxx2guTU5/tUFx3
PWjCkLUkYy4QweKP4EHKf1vS48fysMe1srkKNcYZn6sh1b8qcPCi1pz5ONoj74ga
ft6AHogKseNqB7qnm0hrypo6XWhCt5YLvvOCR/3RvLt5KJ1qTnsvDB6bnVd1S11G
2TsI66uhIyIaijB4mYBK6WocA2i3fax5ge60Hc9inOz7Fbi4N9eVVmnNGbPH+9z1
lohnDpK8rSio0Be1ds+tUuH1EXGWW0GCT+6dD6SjZ3Bp6YmcqIgy7uXIIorVbFlG
+BFMREVWAWTXyVkixh6XYGqBk2C93yrF9UG+WfjGKeFhv7BGV+12rWQ2mT2NHdRe
Anub9s9NcirSDSFW82Kzr/DLhQcfIoHPIbQKiIJk0WYN2negMoyamipivXetFDzP
KnhlL98eDYZ0rpyO85OcG7SUSI7wvhPd4fjbVom5kQKigAxF6kiyzjA/E5aR6xnD
OLBIQHIzeF2PuU85Ry+dkO0wltfWML4eqz4WZ8TGUwH5S0rTuMjWmwSrLXjOsF5m
oLJHE/x5WITlLcXWfaXFzJp+ugpIZaduYK7qPIHoRf09YBWXJwGerYiMxI6fmOgi
DexypUu/Q8Rxg5Jka7udx1UNBHrgCCXl3OM4wfVmMCVibJ+l0rcgXNp0EjL/20WV
Q/O59YYYC8ncxxBpW+TfJZAzP3qxjZb/DZg+CCZ7oRZfNBsg5XlPwRBX49okqKaI
tib3WZR/vLu4bIvMmjfX3UsOEOw6EFMKg8CDwVD2lgYdoBQ+Y9M5kwx+NP1OOVyF
SRcoid/9ZTyIhwGz9EnF8hfAuoZ9dZlHMXkzqdd+TgKmwCvH6wFjv3X7Jo1MVxo8
dliLChYCNgOkILJ10EkBgTeplQ+7O5ia7KT4b4TVo6Jxk/SHAWSyrZLRUPveyKOG
Iqw8zGZLLI+5NJWHozaEqu2AF8As4RgRTZA57VjonCoFMEnbI41zLMDpzdxVhDNU
EKdpE7qzrTOjYUWB7jac+LymdGstlA+3Z5WdbqYVSkPQVHAbpfaWUNJBrI4WP4Fp
FNGg55EkpQ5jTXuTuozwol/AXf7eXJtMgqaVJ2FW5w5TRqZhI8VMnNxqp40SBNBo
eNTwtz5DVPevxsZJqqfsH8gKVCQyEpMbi8nHK8szog0J3G9ZZXkNLfuond1pjIC3
8yRy6gSPNQIpdiVKdCKjkvoC9wv3OpkpuDZd69a4jbQ/2CAuUGhAlhVulYXxKbac
/kDuGt4FGo4UN6FHrnJbtn6u0nCFtTLNLhsiizqyzqienSSekS064QfIwx7yp5mM
79AlNxu7OZ0wL4tNjjlN8y2q8WqRDDhxPWJJ3v/X6Tbdm6l9dDcaVqdZun4Cz5dw
AjbldrYBTBtUJeU6B5c2olATPaKy662XoeYqZ3+0qFQBU+Xd0qiW5WEEqa4d9Kpi
9qBzS9aEBpp8vM4DHPTO8pyghY8Ji82i+NZFx7aI1gVpYhnTwlwrn+oCBbzYirxM
iGqMGyxoEwAZ8IXhlXwKpYEG54vmDtBBJSAaDv0Lg6GKseUcM9Gztpof2r4L6l3x
iCQ9NNWSaaOXBiTu6PmGog1QH8GeW8du3arYiPpGGGsdEXlRBG0Jfh55A5eN5Ulq
QAQey7It6e/kJwDNUMopqAH7WEdf6+SUXt7/sSl6SC3dCKchRUzcNJ/3VIK2l0uF
5hG1jiT7QQMCzUz5N468Y5jFP9GZ1lwaQHkSxBZOy9QqonWXw9PNGSEgtbWoLOuc
4ULxXWJvechXTssu4w0534VQy2LZkyXLbCaAl1UJ6ogvtJwLpZ3qgVz0VdwXEtQU
NtWIyAMmnzN6Nn9+LVKhsI1UTKI+1hNvtJ/jQ6ar7lBecKnmeeqGHI81MZ2za239
IG8y0go/EDoUplNB84hyjDKlQzqoEgIiPlZGiLdyRZ7sEpbce4p50PaOvDnrZJ8D
frWTeoyOuuiB2UqJgVI/LeidrxRSNnjNarleEvxmZHmoL2dmUBOwbUJ4zUA1JqRe
mBGZTcmJIl5CDz+cj87BCiK91wJWUI0ojGXvJfMyieHJq5zXE8++V0z7SCZ1QbVj
2CA31U/7iHafJayMr6kl/571bwr4o+xuSrgftJEN/7OsbmZQcCnoJ9Eu6xXW7O95
tdoDrpxWjK4ZUi0NKfeFwby2iQ7p65Lubio+3xacIR33sqYRaTfAbaHYWwqVVV0j
uufE1DtXM4vNi5kclzQVS6NSeXY8k9DhmQvhBAUbAnXtKADdS8uAOD4FuhkVQObm
zhQJqtxQ5Ahkvyi2W1UyzC5rQ9k5GQPHMvoIUZngAJrZw6fbCxiJGW1HZPuC2scC
zzrjAB0dno7LT9RZtM5pTlhBMyAkjn1FY14GvcVT67hbHcNMOHYdQd/ayGWcCJIK
k8Wg/b6EYia8+s/0bVZiAOqN/ABw7g8HsGZ7CEq+Rre+QBW0uEgalZkfBgzYt880
Bv8n7OpUpcZ8DWFqWn5y7Cx0FlZdgLqTl8DrBOCL+YOxStvzmybgycH/KgSVMaqa
H6LoPyL8qoYMhafR0iTNAGuX8M9ESDFz/0Ck34vG53DOPaxdcEval6bS2fbfhAL1
fXYM/O8iFGh9uYYrFAvS4ltwWV0beT7xXfvdo0WQzp76lEYTsD8FOGmJdBS+30Sn
9+8gyd3dr2UIwx8r5ViyeCYcw2zb2TnxlHHjKKtp/wBTEFog9sqUtA7CA0g+pmCz
3ui6xnAoGEQYqANde3CF9osIa2lZh4kUuB1dOe2+HojlK7Y8Lli+5z6hORgLvKRm
p2zobQhMFtdLpDe0Mv/t8KqYs7seUw0vPSy2rjW/126zEAtjMvwcFTna4weanqiI
mLWNcBfu3xKrsBzEgZguHXczIogDi6aIfgfAk0gKVEj9H+DXW33DHH+InJHhBvi0
uOWkfpEvXTPisdreX0kEJNZDMX0bQladL7Vw5A17VQs1kLjE7/XKk3CtaZJ8YJ1q
x0JZIyz6xNANpPUcE4eq+gfEPBMQmY0OuGQkwqcBegcasx8wMKfqJPg5ooGUFBoz
IaJKEdUSsirRxGpLbBHZbCPnr4RB+SxSpRGjGbw+YtM6Tk4sSTOAUaq7XWu3yL39
Zwro1crZfvDhC1XB3uJ5+yURBLmsvtB7e9SIpr/IEYAWAJu5c4lYaC4RNbUpPCtP
QckA6VCmaGt2tWvnXIQHN3/0sIzQP6Q6ftzWznaHgdAV0ytcZHzuelhIzIYoGbS8
RNlxfvu9rDb0SI0WGFTGnLjD3ymFvIrieZfS7swQiFW9zT4EroRdUuaymLVk+dHf
E0NjIZOXI6Jccw6VK1SlNdMzJS4RzvcsXOzGHHFrczIo6T5SIUG6FCWUbRKtu3wW
OBT7FZqc6eLhj+0ZSqzTXQ5Ma+u/FtEZ0oaCqpUp7c7EjTlPgVyoXv8EiGa+uOXm
NCPR2r3j0bF29TRFLuqPavCu80TszAeFkB9NCSe4yQGwvXNG59um0qk91D9qTQKe
guiZbYcW14jMFp7Ld6CvCoNhUI/CuFYhBbtovRQ2Glz4U2CHGGC3JhHn1VoKzrkk
KDtYmHlNvKFJRv3wt0TV0yxrDbM3WZm1kCn1EcA2CzayRXwaJJU5+YgJqPGoRD/p
LPVIUPWp/Cb8xDOQfXjdlt2pCEQp35idv9c5HU71BfIY92LILjMB4qn3K5UcX/mJ
fvCY8PA+lUaGOeeGKbMx/KOP29TWpOAYFu6qPLQKhvKQzeQIy5NyM5CAg0y7Neft
fEC1uJgu4IbnkFw1KTzFIW8mDjoxH67dwvCH8heLSqh5dNNyKKBmANywV9z89d6/
lzR0YahJEuOMgrhMUyTSoOwhdNNCVvWTHgFKYWKvB5Quc4gwCbUXJjmm62ehnROS
cPOozx/kCG2WDku1udcmDynBBRWlT6deUKRVBYTb9rFt4vo4bO0Zk7dEUVAoSS2h
cGT54yYZFgvL0ni3qNmBjtcn11tElHtt+4ZdCNHw+fJiwggfJj4WtN7t+dbpc/vp
bZToTRc6SwrbXTBy7AowG+eJKXoWgBNTpH5crNR+IZSZF5jmvjIHP7wzBguR7Wjh
g5SLb7ryA/4p9uD26QxoYubgBBXbcB7vkjaHDttGBVMv0Rz2C5f4wpgN99mZ11wH
KWkfxjJ+GVSsKDv9MUFAs7+z1DOLZ0domgcDgqY8AMsPMFWX074ABtoXr8eGPw2I
YfJuB+lfZYcV2+J/Ouf+h2gwYxYf1T2BE7uhoh6pm+uOrfS5fPfVWiQlfE6gV+O9
QRjU5TlNb7VuW+1f2rZ3qWuyAV6BoebGr0kKSGvjJIIw6XyTZrWlDHO4V3/zD47u
vcguusz72aDcYGwBd3xXy0V1KRDOxobBHGwk6WbQY0vQO1qyHDoT6l3UNwoDUw6Y
O2V3/BFC4TQwhdWBamAtosgWy9x/m0HY8rzmVu663GEA0qJcPJ1ZRcb3+QBUCDNp
HzKSOjhXlisw+jv+Ti3W9VQQRIPpu7dRzkjH0x8KDB3a/5QD6YC1TTg8FmttW/K4
XGpOmbXlYXDQZGipjXgA9/QnNo6l5LR0Jt1KZyatkhdxQJQksTLtxCFBg6KrCnem
m/JtCqSx2NCuVtQz/fBOj/ctJjBpSQOZ5v7kfZksccWhKy/5KoTNfWkiP3InK1xb
6eKfAbZvc/W3u1gRh8Cpu2bzedBIeroYShYnAriFtjNjaO2KoBbenENWMEZ/F198
z1Px0YC5DLalH5z78gvaYYP+l+QyH4aaYK0LoUcOmzEWox6cW0kWz42E+rwbNcX5
ff4AN/HVMRWFK7VtBD2TMVrH21nUmo2TjjzF9ur15DzlgVxZsI/TL+ZWxecTgshB
5fKIfhEg6Ube6zpQNrM8mfffWg641oqsZne4GNHeDGFr9+giBoxavqX4v+YVbSN9
HSIWEIW5qEU8wPczFC5hRtD2FvgepdKDMRSROt6hqx6Apl3Y5jfMxIXdi1nUbcnz
84djHUZujtsqN8PAXaTkmE8NAZeZL4Ye/Yq/aU03Jc173AJ75X5P1GPPIFhw3ANy
6h8ISomcTEp1bn4mTqJtwdkEYrxR96UeHBUWaH8SqhKCb4uyIWyrPDx7ovhW/uao
zFv4uYP8yg7awGlrbpdnTt1VYvvnF4pRzGXcw1YM9WVeXt2pyAx6sRrZUhusIU4m
g+8t9oQFj66HgueqtamJV/5PDmTvNnGwS2YFRpyawgW5Wg1U5PaRHYigagIOHHmB
6jzcM8+WZX8nLnnRfGV8HoYkhsDKljlfHZfcuC22v1CJ876S4C+iv94InjU3xnEw
bu8xGeRdlEMNKyAko+yZiULohCdEt/JdLdN4ahibi3HY61QfrGb9S0QhlIw1eWf/
bZBElhd4StBRdAP0nNijz6kWInE4ZszyCOfp9ew1Y5V4iBu9h30ZRFjD2Ox4+KGD
DAJVOcgGjDcSE/DuR8YJ2gZzm+kf2bNG2mytJOKI6bc9+lYbX/mX/AeyhFY+dcT8
xC14vj8FOUAofluB/8+tZD/T5+w2lV3k8jIEihif057qwtgIcRJD9kTLAFCIzOTn
X7r5ALeBJCGsj5cuPJ3bck3E5cajGXfzF/+qpQe/MmHAyPJsjvE999wyJ4pkRZ/5
rKl0MCLLxhRKQAki901NZcmRgts0i7Y2EgHKN8I/GYYEexXhCBPfMJTeeguUfRa/
R7EPWqcNii/PZl+IpyHqybCVGbhRhOquiFK0xtO3f6qVxFtlqmz8HPz/MGOsZ55W
eLCPFWrXyIKFlhdQhZJDcLpTpxsaA7jMmsnLyg1EhJdz8p5U3CqwlwsHKvKBx79Q
cJT+IQQH9glro//inFZwvTBctiXVAfYCLDxsBt91Y0bKxBgCy1TRXMlvqGurgmkg
rXEB8nEVFEDxfANI6TcAP366zIGRJUDjoV16okQ0vHFVuH/qn0OBjuYy1dC+0RIZ
LeMlGw7HG5oZQlyzsAFm+3qGvDdESC6qrdm7Pq1g0uNJ//rzZQWTNY7rDDXCngGl
XSne4I/RmFQUkX00Zbrijer7dm59pMIo5SZfkBwUwQ1EiE5Tzo4sXJHq72Thcpf6
9GDEggmX4qLiWiAVSVaQO1mgwSvyrVw6FyqoQWqDf/hgirUsGbtPT6FAijXcnBDU
l8bgRw9iFJ4HzoN+WHclUgio1tbNu3U6kNGLZHH0so6I9I4BWv9GEbYG8/EjRu39
x4LOoTVIj936TQwUYzXssnIhGJj5sny85nQFv7Kzv9S64b0de7JrR2iqcZjJAa7J
+NY8TfbgtZQI8JPJ5OMqCS7FTe69E54IS1wKl0SzcXseQGWFTypSPtoHfHzGDqxW
ycg91+XLRkC6G5hWrUP66C/dpJW1c9MZ2yvGcCdzzEdZkx8ryLmdHLwr6l9uKyqi
iUMM/0fchNTnsTe6+KZCnRoKAS0II7yCVSrwHIsjQQuUPzTc4RlK92ombWBPpXuw
TfQlMXZkYQ8zTuzb23d+Whiq9I8QS3ApIOP1Rdd2/pFly5TIuMPSRKgg2jNMksbW
nKSSxrrxPbwf7gCOJ7A3cEHFlemix23ttqnTtvR65W2ihRPsLM+3JAB2UXaSEWFK
IFJowRa4EcxuNd3jgvyMNrt3Hu8r6oaPJtLiiU8o3WDBVRzYRh8eb3Q91zIF1IMH
4KBqKJ+caCLrC/CxBgpduNN/ZAGGuu857hJH73qcULSylleJG4hobFMW6Ac0WWZU
sLg2TtccpPOPcYWzuap5PiIhS7/P1b6HMOi/wHxWUnZjaprJ8F9eCVfXciGuf7AQ
+KQCEtKWM3dePy1S/K/RiB3ZqP+jw/rI0XrYcyQc5k5QBULjP6RWI76/57tt0VG1
ZrFBYpLvLWhNgT6dZIOQJ4dzlPsKAt7ze0taE35wsa82TgK+HdgO935RzUMPrQCy
TcJIsPKphf7qWfxHzKTxIg79tRqkSpVNbfGnQF0mNx/XHyOUWe7IM0oaqD70JGdv
7B3L37Iagx2CDrM9IX9+1Ij3RtGI89H5fdelNqh9wdHp3FLg/B2uP1xAv7/ukcaR
eZ5gpw9JUcdNGzmNM6yYW2LjQfGH7Qds50GX1Uh50N65rWmnc4rANx5LdxRW2+LE
foIEKOFILkLblU6yMvqsLw9RQRZdxj9VI4d6Wb5uWx7R4DVApSwMXX5rY/I+NtqQ
CRIIdRgqEx2ITRyfpC9HlSIJj37NhRgVe+eoqGZy9ODwTAHRAmybKmHf1lGHXsTp
gzoyDskRUk9HA88KbYyxQ/7dqaDrBprMeRti5Jswcfb5wtvQPMTK/nsfV+x9BWnj
dTt53lw8YjKijLMCCJo64ruvDubHKp4+/PtEhPbTqYePRbGMBZ+vfG8LJkPXE380
cvCtVwlYDMRO9T5Fkf42yfs9HbQbzJUZYXkC/WufOlOtrH0Z3vS3qB/uX9tG6lXA
VpCIq6PHypmXj6TILgGWEhb6lGs/Iqt8YsEGhdrb+eGp2Ib0zPYwerTAy7ztQf93
/s/qcS/mCvzAIrzm12HlJkrMwWPMydp9wrJyIzY8buZQOsqZW4MzXrBEsqREZOUF
tEo1d4RRTZ+pV6yZ1frBR66Nu0fbc1dz3r09Xc2AZDkyoy2McEHJmmy1o3fDCMYx
YKhwtveTVGEldytVqWr/tPjtrusjEClKznN6dNZAsPlbKCPJxyKE9NpvQ9jNztQE
U6snCJ3l5NyQyFYUt0Uxu6MCvzlCLEreWKJTUo8ZxK9FL2hIiN9bYp6ed7EKARNy
IvW2HYFwZjWFJhG/2G9PVu5ZWcZQUxRh+qMK02bMN8b5e3mQR5I0JDBsE57+6AhZ
HT/1Ft1o8VcxqIzxEtjqXjg9CvDuB+Dzursl34NEQc0hbsp4NdGwiupYu/n/mXZq
MJJZR1rhZKc1uFSEBVEdSyN8YlYbEtwVDTEZnfKQO/u2wWGsA0k8tcjkWNxWdwLc
DTMxoM/kcATQFmvTh1jAVKcVrc14nnzmO5dW4WP8daXbxAKY1D/zuqflt650p6wk
Ey2bsp8y8Uaf9ynbgRXQIVDeJWvORAfsji89Oc7lUCnw05O8A/8r5nFYXWBhCf/s
s7/JrZaTZexxGiB7zHhxWy486HYGRNFaNqV6pzaWqx+2TYFK9i9VwUfGGcAEAQ/o
IIuaJVrGwG4yVKifZozCq1hjq4/ZaX737FkDnUZZ9b/5Uui0gTSGRfFkVB8SMYbn
krvslx5iIBI+axTLdNCKJ8+O4bSIS1r3pnBcNlWq1vPNLVWnwsgMLY77afCBjfKa
XH5jiIWgqDLHtUl7yU9jVEYSFWB14OfBx8IHw2EVxudLIgbJKNOSFWaJRzZQcQIP
EuG9WExZy5EaJzuu7HSfovckLsSixB0Gg+e7sMB6V9w+NSjjhODQ+gHJ0E+OunKD
aTrLLOGnk3v9liyCNR7kGE6QKoKWzO1dVZJjEYRFrd9QUlPaicqNghgS9oN/NWLe
BK9RekCi6FOLnbc9gvPPBLjoJ2mWzFr+eDHdfXIpk1PSES1lb9lWQiwI5DmdfcC5
aLkfM389iquPNPrBYF4MttTUZ6QaHnsAEGcMTpOxw/odSf3iSeoB+gg9TVIqk8jj
FBDlXZqRNfeViS1iFWa+yzTRFV5hFYKlwJx4G6D/gUCH6EJI0/BINEJls4AWvDPj
fyLm5KOebOrMLls7xbDhotViuPHfSqmN29Qfkeejb36fnOkF2qqUihw4NPiqsaAc
doQo/LR2qQRoxnK2iUVH3CAlBwn55UQILWyGynvzJVmV/Sn5E//62pbKbf/7XVo7
X1smEL3o07SOKbEgSR37F8bPW6NDfRKvloVN9i4l9/51q4Pet03eu3SmRGYm7iVh
kM4A8CpT27PSpQR9N672jNN3FkduSyvfVJszV1sLUJl0G6CUezIBL2Pi6pH3jc0G
fZK7n2rI6kH7eWQOC2qnRZi2qtPbt2l95DQVvK+/EoXwDJVWh9s8G4EDk5o/Y+ss
nJduEcu1G86+tQeiXY3s5PY4vCljCYILMUZDA3ScP30HSnwn1+LvS9/c+xAsdWEJ
I5/1aC0vfCI3+1zJDH5No5UGKtmmsOBdhn25F4/cQnFvN+ySHNa7r+53+2UPXyx0
X2ILkgpeL8BLSyAOQ0f1oXpyFaCQ1CRELY74+m+E97X8baDyDvQWI/RBXH9xjtFm
6JR+ZFoE3jr5Tk35kUsnwdn/wIAHBwuinp08HiyGk+NeByYXsPNQrn7bbbhFMmg3
4zVb0oJPwi8V224RzG6wlvLa+GsDCYtFIsDKIepXuRsuptKKHzQaKYj4vbDWsgrI
woFinLYoIFlrVoyymm3eyZi+VeTfia+1It5sQGVu2c2LREKWEcbc58SFXlGmbtwl
O9oWBcMZPtvwR5qMTx8t9HfLNw+96kSrF7bM21DUtEvKu6++yhTDbJCIfrHCrFBi
EhimXj6mxYo8uVJUrEeuPSv9RQBzlzrq1FlldMlPM2shC1xbQ4JWGt7bwq4w2TPZ
d8FJBgbQCF3FQ7y1dBViF45DgLsZJzOCYznlXZfj9ZMBbOuTPzT3kRpeAAGncFyy
RHrRJeFvvMNM4qpi/z/EhFcmOBhIpUg731eQvKXyzIhzjH8C3qFRxsAxjrNkTr+S
iFpibQK1Y4Qt9AyieFsmVhU0hWQfKj2Ikvs2tMTOmR1PS0CHVmC/5nhaQKMEQm4Z
38h27Fyli4m7jsnKWxjxYIj06N57LE2D5Pcdwl78hIIS1bH0hhhFQNb6BGWXCfqE
MjzBHQ7RSiNkWHJBOW4Znilu+5PUHZ3HUp+f5Asvufx0AK4CL5h8fnwkVRnGlhYj
YbVOOP30CjPp1KAwccXviiVqFeHFsayUR0oW0xePAUniexk/XWRpfjPvQ40jIWFm
5c8rzIrQflf/Gw/4EKj5DjCNq4M66VXMm+wkmrLgFdm7+yKMVZ8jF8rBWxazcFhf
8IWmHZwoEM8a0dazuI9LUjzhNN5Xw3KeDHOB68F0eXVhxKXQwHAgQ7fxNSuvjqoc
uK75fH0scEgy/gfS5MdZvT/YwFybhpJ8fCuPZo3V61XBVM3SnaDntZDyNjbWgHTz
6rH39EGeZ10UIqBkoFFFavrT9/EAqhi19uV6En1nBV/ON59ECP7wUxo9R5J0QYzi
aPVBOjFlSW+C3gyCBb/hbs/jKDsRnJhvp+pL4hDQRcNmIedQebHobYI/cxOZas01
9Ko8yowaeUC4wM1xElXjRSug1FVxKqFYl7rm7+iwCS2/up+V0CJtBzex61qT4yOY
IcQfh78p73pFd6ABFyeir6q9fFo7M28k/KLXoi55Jjd4zxjaUXn2KQimozwtTsMP
KdkjfUIW0s/Ylo35r4ImvN9RSHqzkA8bMNmQ5u1Vu1HDowu52jXUJ5m59t9vQ2lr
SSMvuvRP/mJ+jFgOdFxALoIiQ9rYav2WCQGC6TRxUGLkVr1CS9A7l4CDoRt58R3j
vSmwaQ85PGpe+1VgvL/adwW7IuwiHJ4U3jlvYXngHIgaeq1gnqYZVBTYhkhvFly8
gOTABfl9XYx1YG6C8Wa+Vi0cmypaF72vx5rgmLEH/U9s79RQJa0h6Aa52IRvRayI
sMCDb0H/nwY5uP+lcdQyRjPpI4At9Fbsu9UMCMYIge3kB6e08enGnHmkEu21NmcS
kI7mSLPHTAFqlyMulwdn7bpGYeOTREtj+yjMwXlf2jIMJrpOty7B4EB+i2D2Jke6
e2H4p1nfnHln7rRC7Q53eGDpUM95iaJGEK050NLJYmOLEZJwMri2wUss6v3gklfi
38bm2XgCv79Hl8pbJ7B7Ijuq3qh8G+QGU4SOnqAAn02IQVJVrEjQwRaqUIprMl5A
+YC4FVKzbJNSIylpYZ18Kgg4jeC6r6wsDux/AMuMuZXMAeKM+Z9raMDHh7DVW0/+
nkKFSfVvtPrCWVSOFMvHxr5iLf9S8v7l+T99S8Vn5pF+RAiZgG345fpOTwYX0rx9
AsBdwTbDPdn9rGSlgYYPV7xq29SnVCIu/vk9E0SfccHzpst7yWY2HvqHfvoqDh9C
bxw9VPAwqfaOKRu5hV4Y3uGAyGdVd1/tMJYFzcbXT83leEkwB/NSpEV9iL+Rfwsb
qp70F8NV8bM7jAgT2+dVGl61EmWTpR+fdz47G7Jnz77tVs8MPrJswIsVUJG7B7qE
VUQATqxoo6n61tu4lBoZRUqJmnxC+s6DxtlwMyzyVUzJD3exHkil6U5GOD9MyZJZ
Cj7iAV/Td/+BLKWAjdDMWcPh5iqJ3YrOD/4u0vcYppgqmPoGjBTfuTiDvk6ckdko
bBXBBBYB1oPsCAv5YomrLIDjQYBVToVOes8jPehLJnUrN8tQsclWNnS8W8UG88FI
82Fp0x+sdyx8l5D1V2/uUnH96hQ+xB1Dv4g507oEuB97PncdfT/D2ckLI03ROq/w
xqv16r8hXm5T4+zQYZz2OJvm0vLcbs6nVHRjJn5qjNGCO33aXpx9izHlxHvioSWt
NN3iwlJyJeBkUfcvWiELy+mKARQEQ7oXRbnsBQUVSCcv038KJjWgqZGeYLwaLPVp
1OxHya2C6B+cBU99f4iKDoPfkneXz0UmYj2SsS5uHhmSsfrwHnOPaeGN+6tus5c1
wcs4I6zPmlf/W4qCD37P+xWBAjf9beIWTQZtVAD41yrGY+UZ2OYzDkqOtjlGt8AH
kNuwzQ9Z+aaguM6eRo9RA3PUX6F071Ke+YGTj0+plw8tN6rpJYnnFSHFmXRsL02j
U7HAOVh7eR/0xBj6taE8QvG3kGBhfszvI0MrgKxEN4GWL1j5UQke3KcV3KRTqJMd
d3exDuLZhtINPKRRe3mGV4AEsvRDrHcm/ToCyAv7AMtll/lGii1S2pHTy0v1P5Nb
nJdjupLatxnRnHEewqTtd1ZSD8jvZlPwoMOrGgnaE/Jp8iGbfrDZuBsyPTYQO/RO
3vBJD1daQh3K6IGrsiDnpqZfE5R/xKuEykXgVcvJptU2/HZA7hf/FSim5ZQSen3I
YyPmDfolL0t6gFwsls+98UQe5A8MKjuUooc3jM3BsdxPnmQsspoqAaGDG0g4j70T
2AYEbG8mRhGkVHSTbVjZwFPItxRJcmD/xHTU/QWmtvnzjplU0xlM2tt5Zk2oXPhT
BfUDJO2fFpg7W4Z3rh2INoekZAAn8MhfZ0mJsOi65z9cW61okgm1I61a2DnfNN6E
wUpv1xpPzZA/Az+4CgvFjpv1Lse6SiWp4f+cPVhOG8VLwlvaidX8+qa3BzPgqV8H
YKKhI4MNVAuq6inqgMI6EiXNETZE0x+JbfqA47znwumJPFCsBxlWrv30WkHQwURk
HMjOJow5lz6fxJX3RYeaDVdBnLP7jgWkg6cOCFe6JXUFDbomBgtuLBjAVVH8nug5
F+s9p7ZB128dzQ2/SU6biVrTZcAFiGcWbFmlAFtLtmTi5laB/a3x4C+8d2FnAWwE
fk8KJE/xvmyxqDw5OQ98ryhr/Zsw0YHESXU4NQ07ChoExBi77s6RU7JqBKZkvaNe
jnych0RsIS/o0kvLZWKzzc79OVB1S/q4k0sZN0n56ZlRWe/2h5bwh65aGJq/MT40
cLyO/yLKCkedSwUX4ksI33bT19wj/JtTf/l2hJNLgtts/VpdjmWXpiB9SXrMOtEa
pagQ0TdRA3mgkoFPgRMiWcrwsgDfq3Y7Sp8CgRgdG4v3VwBk8Q4XEhF0UJy08W+F
wJF2s81ZV74ZtlXZgvVH76bJYs1J3FhGXwTMcw0w4TATCvKxy0bU7seB8ktKfZM7
e4W8aWOe4vIZOQJHhDf2gLt+qukAmpVS1CroWGjs6SZBPb9+Z2EfWN9xtEsx2sIR
L36JEppqHQ9D8wbgDI9TOR9Hp4qXIrBlTF/aid6cZBEgdxt5Pa8wMzipdfR8+euL
wF1WLJx7/h7eQ6vBmrK9mrl8HNHYM3Zt5mJQXTEmk0Fwq4SJdpdZPruUtjPv0VM8
sLRLEwDVMbxiM+g6oJBflKM+MlJoGn60EIoq2bRfYgt4tcmhGT8BrS7i7NRnncKb
28q5Edrv531QfJKe4AxDzHfGF+M/PjnNIYoBM3lPG1kBUqzfjAbgi7a0vjhBJnNr
VnXgEX81g1RSubWp9l90lZ4VwWl/or9HLb6y7rXCComOnpPhhvbsMAI5D7BFTuc3
bB5cLuUhv/1rS6fZU4OlPcdnbJNbeTm4JQVbvw/Fx8JO8rfE9Bz3JfPRYyptasdk
MeJMHJEIxNOORhWGcnbELKTSmfmpcPqGydSKtxCKZjyCqa62Xq49JSBkDGy9tbEd
B4HcOJ0F9kyes8Q+Dd1xkXr6gerYQwnJ9aSu+rDBU20XCdkIlDCt3yLHbyrKb5wN
gOV1THDMMxcn8RX8KP2QIlHeOE6d8aGZ1MQGH/4F3v1E5zXLqFXsJJeUuSKIlsq3
KT2psPH1ecDrdBIcdnBCvkqfP2JcDuu005Wyi3BOxEXmOKKGaKTTPa/pf+ND2vgv
0XSZcv6xUNgSRYsHyjTAcL6Al6fZSyTo22zvrJzy6oo5s5FltgFAXUx9LPGsrl6X
M3FUEy5nTgUswhKd5yTxHk5rvcVfmDQ4wPkHoaYZT3tA8cj7B4vh9BwuCAIZlVHS
xSIIXptVwewoHuudnqzIxmDInLB0m3dJ09Lg3zCN1+uY0cad/4fMfWQwPfu5ZQSR
VMukWo3GYekcR23u0twUo6dEkrDte6aJz/pFWg/js7Pogca3C0lJXcxBfo4sjf7P
zGJHch3cR4C4/Lzr+/4Umlt3vp0lYoAwbUtISVX+I4hZT2EX8G+6DHKs/hKIW3nz
E63hpLoLcB5WyTGRSK7lGx2bq/0p3xkKXcxKnLnjS9wNLDNSU/rc8ZEoCOUrdfiP
picrdbKI6fHe2BGI9BJiEIV1fPqd+HvThEkWtY38Edbo65PZGt/OJ5jUO17AYhSL
eIE956pkr3OJ7Yli1svD8H895VrbR2WKivYAADUxKkHTyy3+XtProCemB6F6+iXW
dXUwCcV2AMRPPTkPvCkWg4XGbpqB3WG+QTcPWfWQT9AqweAwiLNLzLwQvXuE0H3e
ziUl6Etk54a+Hio1IqerswMXhMwaVoJ9S/BF+52cvI9TaR19xq0cGmN1xufnp2r5
SnK+LKCbph809/SzGoterLMsxygCFQl1hiLfY2BfRgssuTxFbc211UB5U44RLZ1R
kMh4NzhFZs7W2rfZ/Ok91KbfzuqEPDEvE6wecN2SsXNP90WVyPono900hYR4KOtt
PONwT5YSAshtmNn2YrwBMXWCTpveTzc/ypgnF1UfoWPN5jLHwOxFrOvEdmsH2fPE
a8RZBxfNxTMBkbJsaURrikfFdjINsFBP5p4S1ozKf+7vAet/FWIziHgk8F9jX1Qk
so5au2qCQpWEW6Mhe7ArW4EXQKafCe7KNh91F0PxVr0sRYiJbWTCewzcfVhH0Hl0
+9WGzymkBwMB0k5B3FrElO/QabChwkVFd0YWJMTyhEDW48CcZRfkN8b4seiO3D0q
mXHYxA62OWgGFHLiuRNBLzHIAIGryVp0vb/IKHGhJLSI5b5dpDyhuRiR5k3EkXWI
2V4+xpWjgIndVJen6zDn6CTCDcOi9/IV0o96Rsi2ulEEWnztbFkEtkGc5WtcsyH9
HHATkHDScS/7EwIcB/x7w89+7Zw4BMBwj/bazsCqOlNM2d/LgY6zxMTkXGN+/Ppi
nJXFmcneGonooAr8UKDLH0NhQi7MIRwydALMSiwGbFbjpcwoibKhaf8yLKxthFob
FWKRE8as+JjXUgzsR/H3vkiWmzUkM31FjgNtgNVCq7yj6lBiUh30OkImjqVtfaAP
hhabNekQ2UVvBeuW2qNNaNa1TtcSqD1Sn0/RokaHNxZ7MDbb/IWQr4HW/+w8dFi8
3NzRk54y0efglUO4Z7/bDQIvfbkonhq+9Oa89jq6MNeh78PyufUQ3wm2aznCzyST
AzR/UUtb3FdnnbSORYZEOkd/NLXD66e9WZXuqXidNDyt8QDbEYviUEAbEGm8O9Qx
X48dJq9P9icrZz+5lk/j/R/zpKFVaRg0Kg6NBR3cTLdjzC4vj/CD6EaZsMWWMTPp
cuC6ICVaBIaM477W2SI4Ybg9pi/Xxy4F3OGolbTx7i5JiGyeZDHbWY3t5jurS6uX
UlHgXU8BxRacVftPHl5NTYCAS+JgXaPl/g7PX70aSnN03BQI32vhNpwEfq64wGEA
zwa+OZz269f4KYSTn4JVNgJKc0mb9/uAIMBqGqi4qohJ6HBw2xff46IGYRazk0tr
3OeutIK1dvkOuJ7hG6jlYPcNIkbLtlY+JZUIlLGVvKwoYLC0VQ8mT4deiYsLTlJn
/+5gNaWu/bFalt9Iq+Uks8AdZ22L7hPJAnT5Qt8jWLntGetfSDvJXNUYuHInQvnI
WtRXNd1t/WefKPLXXDlxpjhZyAfZaDkV5ZVL1IZghMv7fcomI6zFnVmWOGMqRpVI
6jJvcJYtgq6k5JTQ8BGWzkvWGNl9vm3/lABXU0BASmNyyQ+zDncNWzexOSvZ4oSM
3bKsvc3ljJS4DLkYMzYyusrU6Zlq1Bwn6ag3VUmF02sQIc4Mc7lM3LJmACzhNf8o
nrW8PnT9M3v+RZBfFFuQGAT2CNoxbSlrlcqkLbPmgcG1r46FMdBzp28lqOG9BEM2
sNeCYAvl3doU4XQW++m1A/YxeJh40vlUogHZrkfNUsLvNHgY4r5W/HcHzfy2BdVr
xD96AevOJVx85+4vZH2Cqlf4pI8NsAzRbxnDP9v/8cWh6Rg+/n5ZmWD+X62ueW/n
GUq9+HoeIuu6QOmXP81MZZgVnXNPLB2J45JHuCHhy132HtKlDu064tQXEd+B63dJ
bwVSuMg/x4iaI0eOy/MlRVUySo8F7X/HiooQ/6CC5AQfKm+gVgedxE95xML5TeBJ
OCNe559Hjcxp5ycVHTAB9yX69ZPB/Mz7UE0ry/qv/s0wAjkkjQ5V6pb8szKqBuEz
J8TWrt5CvF0D0NIZ1uvWwTxu3vgRtE5GByd1IxbePJOImXUWzc7N5YSJsPsBvUFO
mtPZDG11XQIYekZexO7xwdtOGOayWo1GPQsANuqyUKD4T30smxkhpoLgf4ovrvSd
UqhCwuZwFITOeQfzyG6BlPtQv+SlmFn7HzwlHFs2wMdaZo5AQmTQupPUggkYrm8V
ZmfayqfgZbNufa/HgauzndmFbrfCTJ+CfmNke95IP23LCjMnuUPHrnO8i9GQn+ML
cVAeA02ykyLy+L2MAOqsXeEHAQl5O0ASJ5LJkjfXzwXjyVuq2ynE6JqgAssHwJg6
j4GYWtCSZXUVu299vz1hVt5ZFP9rUhWu7PvEk++tt1VqGz/CnyPJmfsbesD6Scb5
Lg8SCLAHj2BIi9s8UUbGEJBcu0gLnC6bin2WPViYvXWUfrh3uLFwobg6EwmO6LR/
oQVdxK0gx1j/yLtBZrOUimDBLrN7VnJSsI1Q/ta1MPe/nlkFqwaOrXa5TOAUkmC8
Onzr3saVtKdbsWYax4fcmc/5HbukyJ000+R7pWiDyL45MVJAWmnGX9r2YOOBH/f+
Br5TGA8iFVcwriPjr4zMbDnFUU42K0M0cob/Auk+jrG/LLk/R8k19BNtZAuLk4P4
9D5A3tsEk0psjvWa25gUpePU60EyMQipmoh0dbL/PP0c/COhvKbRHQ/JDY2qYSXO
6I9JyrqNYm7T4LnQvBO4wDAfHnBc1h/mGcVZf8wDSBf2nhMYLLLncoKi+W+dJdWW
yL2h4f3q09MgLF3DoLcrTc60w4qdC2zO/tFbNe9Yfw4LXcE6E1P1MEUSoLPQseo7
MJPn/jrr71NOCgGRWYBN/o/nIFqFauP5NphPQEF8pEQ8WK4KgRsfuF2Jd290OOoU
V4jWcv/ZRhwnWnsHAPLUDgp8k/2YpddGpZPgLg6Phzqsoh/X32VQW9S5Mus9CjsL
sxoSe8en81NXoBi3GBvU90q3k6JicJjxf5r0b0DwsiwY2i4nWAGwsKVoVelTUk1F
WxfJf08ruu6iNrNuzIcaKPCTMVYgnyGQrbAGHO/z4cyRGzOkZdWpoTDiPFq5sGrj
ZdUQ8HG2Ofl4vOIxnJzCM7kH2Bj7BDlWMvR4J7sZDTy5suFhhKqW6EUPT1Ce7XSa
3NzV/qzJALbkJKeJpkE9TOFNzUf1t7PXe2iiIzC7M6qkNbmhn+NbQ9XTpFBwdnEm
im7103JFdkq7WqlSP8I3G9tvOhhAs3TjDXBcW2Sc5G0XpumdcFFOZ+XbZT09R0+q
HtAUB2AQMAVR1YxETQvBcernl3aOrU4bYSk95WMrfA7RYJlWa06iy8WzA6GKQRuA
pASt3e1Gd6cPjpQKaTg9Qs1RqoKVgNRepZ0XiCCUhrAtHIjdvNUk+2akvEtXe6Rz
2RKvdkaDgdb0vAWpYfvGZiAWEQJ2QFd1fowklYnXQP8+gdBqq3u1RM2tZPh8IcSt
zR1jwgY3MO+K1d6npRfwa8SniVuCt2Lpno6AFc8F+q4bNGQgvWIWeQEp7m6CSsHz
BOS46lXEttmOsFYeE4rWmH2soQqYwn4UKkFdnuvIsrbSsFBUD6ZGLlglhZsv7Ujv
6imhV7kLhV4jhXPiKTZEuMvo5Jr/MXWKkWVxaLIbVnIkJIZCvu8IQ986QB2o74PR
J+pkFfAkjVOOfZU/obhuEHeGUw1ucTuCfKgOMt+lCpp5McGWvqtJg8A9UDYCum+n
QvhWDALJeXH3Phhn5HajSfS0nre2EUtF9gN4rzhhGBbfYr1mojKIbKCraeIHy0Xj
HzRKal6HHWKd0ffBvEsK/HJ1wpPIvJF79dnaJ3e29LVsSxqj6auiG5r0qvqDELH0
cVsQIMjvUpZ0TgE9aeOwNtF95rnoS9PHCn2fYn4Wo7wt6YXij6pY8SfUM4GCRsH9
basPVHB9cyoQmb41arxQrWIaMyLjQX50hhnxxHwlXWNIGNQtK6Ikffpe9wKftv/d
IN+vfqAhQN3J3n7Z1f5RtJWiwkpoYcARnLKtegtHh5ru4U0+AEr+bxyzhUqkK2De
qImZ/HuLmoXBSO631MOAsIb0bDQUtHtgC52bnH+z8RIMZqWxuhH/VW234R2+KBUs
t79WfSk3g8fBMyHd9xULREYG7k/iSQsu9j6avW89jxHNGhASRADVRiZ4oyEBE7Jc
RAeoh2PVpGWbvrHHHLpeVdGL2jjBOWPEKUQeu4D4DAJ7zHJyzGfAHDeAPmFwhNPj
ePU5V0vazVeYj5Z7uJiGhln+HvENXMue9QiX/tQWmamJ0TnQ16TuFP8L2QsOGVAE
XvnLwfSShwRQIWSfnVyCOmR+gfzujhkQgAoxfaDg5aHW6m14N5NzGHGuuj8VwFYQ
yRh08OygD6lrBvdqI+IqnPJN32PS9EMD35ulwwqf3G+l/ux/JuBFTGPJuLLHWw/I
Qb2mZxWqjrSTFBcmPV/bpqxo/1tJbLN9NeSRY0OKBSk4yOtXDeZxw7LiQ7zwgOIW
zch4tmhCXKOO0jjgmUP4CA1YRuRxfwocfTNB5mZsP2FBti1X9Xk5gp1aF5+cBTxD
6tHpqn8UXbocgmocJINFIrXuFztwzDKWZq5p5bQm/6In5SibdBc1Pih+pASZIIyr
GeUC+HqDOv6KezjqQwGWDZYPJWhgQL8JVdQ57X/4Nkxa7saNy/ChlhSmth+UBuuW
HwkYXdymS2ly/zOmblhQWzLvf/zAyJExL5D7cDG0FmMyz0BcyF6bPZHT+ax6be/a
wb1CpOvQ/h6ApAYqLhzaUNERN+9IcHDXVMNwJkVNhd40stWjBFL5q0q0kwAcR2XE
MkXDoaU4RmW8h24P6fD/KsQ7Rc96M8PdqfBAjNBuU+41SLRGJ3W9cdYrki7DiQhO
wJBNxZboFEVStm5PUcvXUPCUJt/L86zxXn3jhZtnrB6c2hf4EajNnhoH5eLT/lWa
G9grnnI6wKVg7nOdu4Zt93jlPZsBmNhWotldxL3T9Ke/7yYqMvbaDrdlGFxzfbxi
nbPyvKRkM5vr4x/N2fovXmAgoRbQjv2zxHpiKfhgzq3XxJNsORoRXABw+h2RGvag
r0FeP9mvuGNF55Xu1reOqyj9noFGeMWiLUoFJ7yKWetPP/zQ9qOsApyc8A8Yw6I7
OzJ3I/2XHFE9TMZhTVmO/exoWWSHEcr79aAO9I9tgEnMHt88STiWa0B3XRlgyqtp
s9hFsS/M3Kb8dZvFyhyiV0N0GNCyaV+GVTku/uKiK+ETLoaP8qs0QpYLiYBuQj76
TMDb7GdmQMvpCMt4TZ6VgavQYFGk34eKQzN+HFzxr0Kt0SG/qCj5mkzBVRWD9Nzn
WlyNKhcjzUDyBTre0PP8bqGpQtaT12/7dDt7KoNL57GGX6GzirYcsyvrS6esgLlA
Z0/nINrN5CWDjlgFWeKX6T7GtATubNvSNGn8meDs/+9DEYe3QWY9vDsKFOhTul9C
O5irpcyhMvnRhzdesOs6jivI1cR7OM1CRzMnEpWVcR0Fp87AawaiMxu6IYyArWht
Pfg2XB1yvCYSjUOcXjQIi7PqV4YkZtzcZ8xOvvRM9pELLRan3IbixQLwLJWikx4H
6pt2MBJvDetdT6EBRadMDnT+OTXlS7BhbHgnzXp82ImZyQhWvTaEi5HRDxNUKXQY
ig0r4AyMv+UhrdkuiUNJoq4RVbI3KzcVcR4rr3Yi4hYvgjKJZBarHdbszuTsmAVh
cq17VrKm9fuY99SjqaoB33LP+p/bo5RYkrMTd0EmQ+kjxu7EfxyRri8B5a0MCblJ
1knllktCzh0MlU6PJTCPoAB1jZb5egd5av483o1vt3dOYZ0kyheuROTNQ9oDzcJ+
xeUGgh1SYchFePOB4quaJCxh5/ZAC4bx//XQkcEZuPC6MyBi4Z94QyRhv5be1cQ4
SevT8KGxOR9hmBgXaCI0H7C+1pGENTUooxCPB0AHO9XoNs1gi5SWxifnFEQq19cS
BFIVUTyGjBkVq8wGQfaXD7QS2i5yoU+pdaLiH9PkEbiZsY29VWORUK8kG2MeyKff
BFPleKwWB18pyJcBOUS6PxEvJ+2uM23GADvIKEjF/hPS/V3H4uU4BtL3Vg7lIX3W
TCp5MEh/HTQLiWRX+QQJhzoog8wifnJDSRnyV+2DHBlgjcO8pZR8WrQiuj4ojyVc
RhbkNw/CEK6KdjwY24f1i2zXsDesYvB130XeVqZoSPnTVfJzQhF8Ssuvhx/QHoXw
ATvnhvgIwlNhjm6oYVtv2Vs8ujxKZ7uyHGHwXgcVo4bs+nDOPWGa5tVn1PMlTlKw
x/v0NOhJGSUfVNQe96IpRpqrL7AsPvlPRzdYEngMIen+JIoRRMSKG1R+zZ/x9PHb
njuwdDs7O9CCVys7jqNk3y1v53LRi8DkaIJX8GHol41Ix0bKN4KjfykiX/lzwIKi
paF+XFikz0zUvpnhJ0wG0EhUXyw0fE5ejt6e9nyL5XqEecquhN08xx2Inm6DQd4Q
BwCWTiyVZZLCcXkt5Xb79oXwlydVGSiaUdETfgfVf4hZo3Jpnplo0rEwxtUehDw6
P9iMVl0b7P3OkIVs6VPWc/NJYE2p9u9ctMq7lX1oXwquZUjEcMls2BV65jV0gx0g
+D/d+rwj6bZaSjxX4GjAwfNTFbWPejnULb32/tyhmFI0hygh0k8znlvOBMuPmE/M
Ak/Cl2UmHZqb2EgP+BYnHuMdaGq1ph3y6MNf7qjyFm23QLoFoyjaPOnQDFq//eA2
uPLsDM9ypfBnw6Gu3Iabti1rYxWWCunj2FqLUOybPdLqoekBcULQ8bdO6CCzivcm
AtHvB1RiGCh8R+Tx3i/7aJbfjxHjlewic2ydFluiXBo=
`pragma protect end_protected
