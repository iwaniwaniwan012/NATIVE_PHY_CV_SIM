`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
L4NE9IPpwo8gIbMVBcRED2WwAu8HlOKBgat3cd+G5CWcWNw3ZCODKxHLENAp+8xd
5QQ7gib3pZ9ZrTIBNp6kt9knKZXzq88EJMRYPJdy3bd9ZGqLf7mb82pvC/RfzEYm
hgnvkgh5g9M/bwFZ3uEHyt1SavGcIc1qGRFozfHqg04=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8272)
W0S3oXfAlErwd2QEutzIIAPC6mjlleJdnunzvgqNL6ZUe5sJTYTmDJ97v7FwR8L/
zKzDG2yHks4z1DYafVs+RH5WSPSVR83DaGfKa5DRg0/XsUu/Eq0INWKoxbOgykX3
YskTodWuKQwVgtmWw4ue62nb6I5CDVBd0TZdV9LvnNRWOXcHEt+K1tEmWlfFJQzk
Km8eoQUZ3daGHQ62gjbhFESswpEJH18utmMlmfbAfd6U2AKS2QW6KzuTeM0Em8bf
rZYrnbDKN8RHuFhVZq3KdJ8apvTZpfiaNVxqNV12cY5InrWFEW9oUiJqEQiVuh4t
+DX6P0Zy2LvHhuOUrWejxu1jzfS06a6vmNmL8R6pRmbUxUAzMaegQ+cwsBXN4O3w
e2HR1o5MFsm/buqCZRoC3f21LBOo30IrXiA4FMeqe8glJs2r7rJKfV7UjPAO+5NK
FFYy+lT1IklBpK6o89tH9p45zsN3FY5a2/3VRKn2GsCAmJOhlSZvAWyniU0aShgn
kJQBSv6rFsQvmbGqcpEFtwkpc1WYTl7VrLvQQhdv1Ug9YYGV3HnfEdWbFd4MuS3v
Ozu0q1f5Y1rm5kdxMI73R+5FzalMcZ6wXlB27pYod1wI/hmll+5Z+cDV/3MOOZyt
r44DBNAMtMOJaEi90GRs+kGKK/s8jFUR/GMblqAGzQLo3Zu3P+4xdBwid92v4agL
cmX/xO9YqnMWSs5Rr2kzbKvE7H3+zLCubeCTuzzjpStBqv4yU90A/Slq+D/1S+rT
8EkBzxdyPDriD+hxgXoxRfJ+sMuvQO8Qxt/sGf2ghC6d3iOziCNc5DjWMALRKDgr
rM2jiZ8UU70bWfUTuZd9XKIWzgFjk65JPcS7fkl4NeAlm+mO5tjn9j+HOUBFdgQn
t/3wCqJzk/FiMUox/TKuv0gUYUc5sRkSyl1H9x2Ext75RA2C3arAOErTzJv/pYPh
EolGJT8fp6QH3LLeFUhgviCDcPymFaJV2FGZ7C+iFUKamVb6LkU2zfDUS/LfTz3u
ndimVnr+m/+Q8VudJCdE2ZPKr0hP1K/I6REuxpmPrkzBJlzcCB7VYm/JmSuIInJX
fpCPiTRVqbU0ejbgxtAePKaLl3S/0aBftf9pBwPezBBnMCJx5PqkiketWiABuMjH
0VQA8fweRFIKptPnsSYYPB6mbwGvAN+S36/YxOSjWH7yoB0sI+NRZr51mJkHw0jA
jzKnTWrJBHWchRTzv26XsD0aC7qozhWkbAlFTMAKmOrwUQZASukHIXMnCMuBJVcw
ID+Tq8mvgRJuBUcjz/ayF+96Ly0w5mqSsPKUr0kxHR8KYjHi5ULhDIVblbqhfsK8
BbiAKDVuzu1nDIxCgqjGx3qsDCsCiQAp1Yy5qV7Goo+WfTbPZ3nl1OY+MtZjdO3w
3EWwiOZMmSIl7CkfUaHUJKmQ3h6PRX279b5q1Q5OQdkpkF+AdarhIASQ1ih74aAY
uQR14mwaoWOGiSYfR9YAUX3knOE08rmrsaML1fi5A4aLkRv5DuCmISo6KRK8MLun
/9I4OwwGoKerMT1xmbNhZIH+7UdQf21F4xitO4hz45s9QQOf/judYYvWJpnZNP1m
muydoFT8TVLjRHr7qGRrvv1VTCioiTpZ+rcMAO10vbzs2mC4+oIQ6Nhr0DHK80vv
F8B21005T663fGZ4PvOODhc1UiKWItZ/+pxaK238TLFVLjAwshXsA3mPz5DMkNEo
pcr18ZvymV97BFmO9A8QG1yBbtptH8M5bLvcKxboCPr7vAxw7H2pdx85HAsVeN44
6cCnLqGIdnG0Fx+1CvWqo8qxw6RbRypLcG13k1IDFEDysYopjr30guNUDmYWoith
5ig7TNf+W9hWceiIsCq3i/PJnCDcCsoOGRJxtU+q/ZR6uapSt6mjgwSVeekt9EaF
un5yoizhu0Sh1W/jb8cQtMEhpPd0T0LCfoMrA8o3+ucsziicn/7g8Hxw0b3B4C7l
x4iTxQ7HBLacY43sun+6ABRy3r0pkjjbqtvU/BfwQTnDHvIPqNXKSdMpB0+Ugn8t
P1uiafZdDZkKGDuWP9FJPbD/CQ41gjDTIUSwstu2ZR8p+dOfjN9gTETdVuPLSqWH
Qn1vYCEf5dxKRsza6ZMrubVA1MHp07M0Yf2Z7vAE7vcVCMCk3vZhCeAyIh6yGwBH
8ighpmIvukzR4HMTAW7yx5wWt/FAY8n2AcgA0lm9izkVgs9et5cFm0rgdGsSGJA+
sPViSFpptq2mr8NaKxolsfUxd3SoexZyYhS0IxaXhR1Q2krI3JdF26OTpouV5Rs5
YVJtActQ2+/sgcQ2P2bxpBbaivCzRcVBes+bwH3A7GgS+uKT1bUYhdIQ7Lt35IEQ
jg2+AKVLIJXqeLfXpr+9KkAhqyM1uIyeYft+Wuq9OsyTTVlBq/cbMCZUgVLzrKFp
MBE0varw7Q7NXdoYgR2iZ5x+hMFPMFyok6zyJYHMq114mzZv/RTA+BLFIxgkZyCy
8HSTEQgIdLkLlOMXRGPlifMk+rDn2OcMMhkr9ZMCMYjieiniWy2IUuMOdomH6KaN
6OaD5qkCySS4A1mobKsb+HDHIXF2rM71A5yfZ0g9ug4sFg+vqZjb8TJGKoM4EsP/
y9+HGVMN/CeqVg86KnynE3VXBkkQUncTLkpiyR+ZGs+zNi1P3cS1VUuFgxorWMWY
BgrhCKLWlPBzZtwpGlpmIgZvOLeVeVQqtD5Gg+ZHKSIndmeRgAaRCrgZ2ml+5K++
niqfnv2LtVXRpiUgMQzBWpgd5H2uasXQ92XckjxUTmotCjdBbJXLbiWd0Kxp4FPO
a+AvLtEgHYi/iqfhZZ5dT6Llt0d1eBhlanGXAW9ZAI6vv3GTsg/VoKs5TdSTAZqn
W8j1Hu4Ky1eFLpDgmt5V1esZjJWWrgChlw2Q55GVPoR3+zXoHphXfOGXHS7VmBem
Q/MXKgXh5mtTVVQe75BTC5bzBSiv0Oi2ZjW1O9RBRmb3Hq7G0xL5udFbolKlNwg/
lY9gKBhKCZeaRWrHeDj/Z/ZkKw4Cg0Xpbn4Ab81HGNXigOvQi+TANEZ4H3L+M6tK
/0s7Og66EBwzEMLqhbIxwE2V2+E2P1Z1P1mbmi8h0qGL+ecVrNJN8qJX2kTFTFOk
mwea5RspBvLRvihjqdXcE0pLHIrc0aMImw/ihCfKcOld4MjAOoe57gdHKwcRnMvz
JOtdVYFeak7K/jP9/DtWGU5X0rDzZAPJPaDJaQMUfdH15S+qFeduuAvGJQjLwmzL
h2aHf2xGFgy9lloYvrfOBr4zVaifbyEY8n2NtwL0bNPXj0i3IWruBcI/29NGxfUj
Qe5Yr3L4R/inZr/B2L5ErJvFgnwDWoKYb+OnUii16sBcHfdkTWlXLcFETvWy/L9g
YmAoqjA1YTYpnoc5ydhWlaPQIR5KJWLbBoGommoBgQLd+HuZ2QNuMFECXywazq1P
rJ54Uj2db8/diqQvB5Sugx45gvhRr1Ta33AzoYATxK5Sun8vkuL7H9O71dBCsFby
0KnjHyzjUcOD2wjt+TwsNIpGbkkiSjrPkHHK3yiB0QrHqknlfwtWYsat4e395+wl
KEiPHUtu2fSP9I7Zv2OF39a18Ls/LUA9fIywXsEA+mouKdazsypeH8TFLWBpm5PD
iwJbl1EX0q8suMvQUqxQaBXYbY9VwrWFMo40JzzuHx3IFy6HUhseFKVUQPNL0qco
es6X/n20n4WeSW/ZaHE0k9pqZMXI/EoYiDI/bLryIpleyC/tIZUM5cOopiFTF3un
1vQu9kExpK58RANFZSMJoSyQhZtMfesW+dW8HWQqOGMafeBF/bDfhte3+U8WgzHj
vDpoq5fcrqhNaaDSgTBLL6DS9ANTmB1FV8qXztxoX3dlnalsnRnyoVk9eKJ2AZgo
Auh03eO5hjZvbjTNWbH2XC1Efy5a3gb+dH5cE/F8XDy6YSbTe1+0kPI+l7wKykR4
iaBw+Me6eD04/e2iWR8JBADqEeUAJBOHbmypjSsMax+tZKaxdrhEQAJYkSRxGgZj
Rqrqkr5TUzH+ALkC4Sx+GunY3rRTUYAsxpVuLTZxH5wesxIbRs7mhoAa29t7ZE/o
SVCkxHuxSTIAB1Kp5Al9lV2PZBLBkVHWFiZDrspnd8XtUZHubxSxzsqigdlBa/MN
jGPtjqregwGYMNqMuNjVWHOeScBk6M/+HUOi37YWjzBvvoU7y++jDSCHDv7gMetH
FiR9I9F1Afmz4yTWIMGIX5mLwd/BScGqiOkqmwdELBc123bTCFI6SrxePBBVrkLQ
Vy5BVWFyQcAZEw9FggqRq582CTh0leAXwHxfGV4QCf+cQe251U9C6PX9mhYyBYgp
lkiA6jx/rI/j9ydyAtioe0P/17xDqyljAc8f5dsUEoMcVjgOVbGU1MVaeoyROjRG
fOvc+suTk6a0xaCynOBUBn0WTF4Wmaa8hF/Cm/70ZI6yIgesNDrRu9v8N9yg0O/j
V8E+XdMepVgCSA3pqKfpKHiT/0hkgC09rQ7/7REB+xrqZqCpl1X+x7ZJX0TUtevb
ze4Cwphvp481MvoovY4iKLs3NBn9XmeNVqiPT+7Rhpzpo/Mxk7FB2Cjvnr5FdkZ4
8Z4Vnut3fU6f9s575QcUONnb0k9lSuQzt9kB4AjGUu502DDezhcw4SZzKePNjqIn
lLRXi+rZsIVhvj4JuOmJBNGIY4oRVEZJ4KKjSIkPKJU8s2Awvd9WnoEDC/QDkZfI
0R+BxlH17DG1Eql5KQ74NvKuv8uEIE1pZO59KChTRDgjIbzDHbGZubauFDFAKfyb
iiLfZ7PhtBPTdeKKdjmSeDKEsUPZTZYEPaNpTM9inV4v4M0/WZ/ZhjrRndjG2pHf
PD++oT0OlGtY9RLJOkcHz+Qcwl0cW2GxNE3kTJEEHB5CaYs0LMkE6gpxaJgCtD20
JHeysytKZa6T4cSEeCpkUNfKbHWE3aSwghzt/uU5Db2bjTfWS7toP0iGqARAc5IR
RcpNUz6YJgjCmEhU+b42G20dGwuYL+AvMbggJnpyJRA55NfYo+Q810NNHnYK+LWj
p2MvadVUuFoV5vS2zv3VzGozQ91Nc957gO/aoNmP8yICaflixnrTQsH8ZUfey7kj
re32WrtXUMlGN+VK90jHrJcibJhHWJmxLYkW3rWWpzCFXtuuuLM2nmvfXsE8qWfm
FPLD8sYpuVpygpuSY5AKyRtweA27E5jCxq/SsCCEARgSQ/h+OIso2BfEm2g8pIfN
cU8njF4LK/Y70zWAlSQrrw1Q2RslhWPGbuzv2nP+aL58ZY+7dGJjAox1rxIV7K8v
lV5/gxqDzbQdpvqCnUlUIyby8/+7VoiF0RQiG691icwQZOOBzCKeqEdvH+7RzMhI
/tgFfECdvsX9ZFbLu0Y7tIKm+yyQ9C2dbJr79myDyR6mzRX6jtBskkY3xgCf4LNU
1yxYKPWH8HiRzbBlUgK3RfbKQMipSCCJzSE7f6m0N8KvwISEFn2NVUZMMw9nhH5l
WwwDa1HqKIpM8VHIgzq2hISXJbaX8Xhkg6z38EH617CebHtBZBLrYuhSOP0/MUZj
nFh33F4mDeArd7dFxX0cJWyBHlGc5ueeTJde4nJ+T9wopVa/b1LB5E/3+LiyhtUG
vBhoaLjrlGCu/4Mhtt8tkR8OZZiqTYyYt7Xr2SHL7wbmPEWMir09Lc3yBrbyZ2bv
9lpdQkdxqMil01rvLk/YYjHz4C93pirPTplOn/8y2gcJ/DI7vrOimKeckFqvRfUq
QFO74E9cESeZwGJZj7RhUq2++dMGCMn6uYbCS6mLP/EFnBhimOPwG5UdHLbZ5oAy
naYoNE5X8OT42MEQUSHMqKhXtjIuqObSDt5aVKi+Zx+o/YmmWeq9QAVoBcjeIEom
BjzbbZeYK4tQxcMu6uRbs8KWPc115gLKGr/ZirwZTVkCnDFN39/tUFhnrrCL6I2u
crYW5M3jXyxyJ5pFysyHrPJI6RP6p+0Z2sJJom/vS60x5Jr8mgqbWRqVGD85YHOF
IeCiu35qV7TfRe5aawpbg4JvQntfdcxXd1d5yMvV6hunTjS3P8ZGP8cW7YTjMCSf
P0Xcr1bCI5oy1zlVf0K7yhxmHs7qflnkkNU1sk48fCB6G+pFlRlSP69A4+T4f1y6
A+3GA2rDyrx1flLdt8WcfI8ipI8ZX8fqmWCe9mKxf08zirTkci6IYh18nRNpJ9jp
YzNiKonBEaJi8rFNyp9+4plle+DWUckV5EgvE7Vlo7t2B/g+Rc2m90l9fx/oxpZS
xB9789M9HTEz40hRJXXj7T/L9MnEMOT1EoLnz6vDhTUgNYkVo3AvTYh4pMv9Sc6s
4EoMv/bkV9Ow8RAUks82LQN10bL3CsJVlQgtWZTgoOMVX75v7JHVT0p16b455mwR
5PKP9iEWrGX969A1luTdPP72OM3RUu03W7/xXI0zbUVwZ+e2bqZ/3kwP17F4TpRh
30wDgEaEKRmXREWmXqzdHJCN53+ZQEnmCnNrwYthv4Rh+JJ1ODCgorSwaL1OD6Gc
2h/X0Xt2ubCxRfq/Ef8vEHJSGclQM4ewio4Sg9xm+K0/XR+QuQs+pkHsWAJ+vKyu
I8O7V59qgxBv/aA1xthRebv+EW2kRyCT9Ngx3Q7Y3wgh9ky9lKewsNeEMFpOb2uB
/oMVLE/pVEtZKqyHsW9Fv3NrAJix3UNdqmJhHk9iUCjl035YfnbO4YdIY64nEaZ1
ph59WSJtKZBmE0prEmqJEIXthI6n1QiRSwUlpIg1dWURdHZ+RLEsir5TRb1OII/x
yCgAbljdlgWffYkC6V2n/vWsJmRSp8lhZdPhIT76HqhL1KTW43cAEDFLRUDA0UB4
afrwiWTIbvldtS5X8lELB+UOMHKY2b6U9nxiBtZa1WgokHgbKYpFb6HENcChMSdq
VcYqXkeN8Rok89mh9MOIt8OJ6qd53AVdz8mi+CFS7uLT+bIQ5Bp5jykbKW/Keikg
gNXF7DpaGub4ptQ2zez5hmMMrr6wehrv1gdNBRgl1+brD6KqKvAD854atUEi4xT1
usEHOUdN0kku8VQUD3nOzR4xJz/UFYViVgwCi5mw5sN/LuQsRcMc9XOMkOdFotmt
glHZnYYYzUVtYYmvIQ5esFRA5MytkoHmRgTrbOOE5hLaWLQO6ryz9hx8CT/tgbUD
yKLCPgW/ZNzs6r0oqhhy9EwLfoVJuuwqen9yhVfRNHo0z+WWMtBXl0ECJWY4Mi/J
Cfoq8OSLkfidi4h8V/Ld5yVsenzVm3ptYpJnPyGJx/FqezmvfXSHXH43sSp27rr9
7m1yhlLyGnovZfIWZox/EHl+k1DIoi4PGoYi+e3e6HK6e0mL3lw5m94kezDuXNGM
fdjs1DWGETqvemb05fGfE6cw0kd4TneEo7bEr2qujBejFUgVl0hz6zL7VPoGxj6W
9lD9VRnB//RXWRWWCjP0b7mVQnV73Zj9WeXYdrAXv2f4VC+qmedQVYEfqUA+RDDr
khb2OoMMX/nTK3mqwgIc0toRe7Elm1Cy8ssGrI72hqClfsFPuU173rxKo+4WaJPE
6NfxzCTuCSncoYR3x4Rhau04vPAiqLEYXkPHPk5rkVtk4DnZkAlMLYqbC7mR94IT
wS5YxMeKCQwsEtdYihLvpHfPUnYNiBQCVo+nJJuJkkzicO+t/pfC+G4m1rSmRNud
Hk3Yn4NeVIA1MPR9FGVEO7EzC1urq8v9ZyPL+WtihQm0SfKVMyqqnktrFWoGqSqK
xgmvLeB63/OzWlhlZbm1+3eFhd/vIefmdbHfltQ3UFLBle4ePNL1wo0szh3iZlYi
qKPFZYdF3QQyaqK892gC3NuUs48LzvU6Kf7AI0YRoW3dCqLwYNMj2wYGX6e33BEQ
xmmiw4YiydC2zp3NXAUADMMMyYH1U75GYOgllTRlfshAdnjDlUyBPTYZZVxf5BoB
+XkkTvFVA43us5Qj4Djy5zbfdYAE2ANIjwCZRk8r4k9hPO5EK1Im8mZyQvA5iSsd
cMlV1MkFdYObeOpZy559TYlFwJ+3OX2c/CNdlbFuhOAx51imO0AFpsEilkT6LkYh
UenwgPukm03El2r2BQS7ey2cS01rk3oTbwrs/9FTPLlxgUcqWVrHQh0WyMUt1fWZ
gXJml71MFCPbFQl4exK5VVzJtleujvifMVcXOvr/WOvq+EDyMLWEjem3pKW9B2Gs
i2T/Vvj16xA8CB017UuaTwMZONhNyq9BlB6uXy5dVO2DYvF1HG3PKHXxJFTLbAO+
fUbfL7Zo2p+PP58Iceir/pUXvZP7FtbElWrW7QgFFAGOwYzs6oWyvH0z9ZdplFIv
nO8B5VEPDkpGoG1iacpCk9yGJ/aiaCeSbm4UN9mlUKniCjLwrykaiE1Vir3c487f
jmw+PqKwWD+hRNQugsiQi2v2EUROgtMUHI14mReIe6i/Tb6+yrj/bHpJf9qOEnOC
AlnnFnDAGARNgN6GIwcyRXiIgNiXTGR7Si/7h/LdsFFBaWKyOnCXPUY+y0HVvOh3
zxYhevzMbJe+wkOsZG4XWIsJlPeQ+CrqX0y8vDhswR2qCT8BNNBQoZEtmuXk85Cq
g5o30wqLYFpPqPhSJPt3kvAwbxlOEy4bDRaUUtWoe9X1nKiPGrDedaT+gUr02ADq
FEX3Is1a/H5TceZhm5Z6WpNDcIJ92vKypZFJvuEToyFGzcfBBOK6izp8+N2TosLA
BiLcBa2xCWq3nS0ReufWTGP8B+J114fD4OAjAkwVVh2aBeG0Q83ODHSLSrS0p4G+
D7Yg4BNdosx5zOdDFFkJwKxXxIJIAjOgwN+i5hj4Vbzb6B5vHgTBEfAWpFi1lE4M
VaxacxzLc9vH8MWzx0teHv+j3Vg6g3/L/oUjEmlAuoBORAczus9WSQ4zUjnEWdX5
cdbatLTX84P0/02UNgxNGLmjoevt6hW3EQzWOGRSUgAJmYNy7j3fvJ9La18zPOg5
+mo2TvuBtja/Pao5Wm5LpDro8ufb0Xq1lcGIGS8pM3JU6kc6qW3NKfyuUylAUrgl
H/mg8UEuz1lP2hz+OFBs06SqBDG32vywoPaD1Wtdl2W8nAXxCMnI/6/ywM4BfGAn
SpYkl+lRGZMhQ0lkE1++4EBYoc1zHtDbg6ChYBQNOcYGm05pD7nUMhy6bk65eES4
DttuCl+JxNLMpppQ9N1Ip1r14lS+g328O1MH5xz+FnDf+LpfXPegSplBRzYmhDNA
8RkN/CuFZIYIG4uUUbI7DDIyiCaKIfQWMpkcsuYyGC8xy1E8/mMRRzE/EmzZID9J
5/klNcYHk2mhnQTSn2z7q+e5WO0lXTjh8r9RXFjL+mBEp5PwhfSZk/akVu4ET5Ja
NF/6piBzEnczN8joGs37Ur0OMNCI5OmU+HsFbqTSlbLm4TJoXXfCJqKa6Pj3b5XO
oVAaQsaNOTn/mzhqVzTIQDCakFoldH1KVOLWCCe1ODo3h3ZEGVRAsL4b98H/5a9E
8mNTRJrnDC9rkkxcQNAQUqPU9JFITC5liThOHk2Q8S2kbJaZ8+7JD053jkPdcigA
6cd3A7t/uWCo//KF4AhMD8/HpVGbDGn/LZBKEsBdjEutptFCwYutGYfa6hNqPaQw
QFy/5czHEhMvIXfkz08AWNwo/Xo8Nh58DDryjtWCq5RSvKUxXrR+LNJ0J7WW8gEe
UlfCkLcxH9eRxyP/fgOg4LhnvOPfjrdldqDyTcq84ych5Z5IZAcUDCjPQ0TaWFiE
wioQBdz2/9agwfeieeN7ZSgr0twDcVHPYMuYBAM7pLOZRUDhLfbIIOkYCpCzNGtR
8h21NeoZaSTZVgVnkXSJCCHsx0hHlVEsLSYSh+ri0A/w3WBw6km5Jaz4mtsRU0xa
IxqIosAbEfRZW3xUuL1tVv6SUjNWTk3hzeD0DDKccnS1qQvPqNFW4/9xmxWq1vnk
EG7irqnDzmw8K9Ri3xi6y/7/oTikB5Z7heKLJO6IePL8BDtkFpFub7HtZE/ve1Ii
IunkcbbyMZ7lgajbjIfyTAPWNZlZdC9LbYcRa938NrfZVWL8xaGgn8V/jkcjHzQv
MOydL+005u5qZe1AjSL6K8IarocdoeAktEOioXMXRuLkRDMVJNmpcp1p5vdOugeH
Lvlc4DpHSQyMH7aKpddSw8cDmj4RD2UeMZasmiTWbchxV1F3odDz8D/oafFNlcqq
iyXBfh+LKha8OvoVXNFbT8iaPZtDZrUdIBuzDhk/VzoSFBU7XopljZVRg0BLKItt
aRV8nMMZAfyDEH1o0xKm/zxaqZ+YO7cRiZHAd3Zas4aZNjMD6SIfX1NYN61goP4E
ftLL674H4Uo4bns668OrPatatNId9ZMWxZBjFQ+go+2uPBV3ntnNMj9euPsZmjqF
PFcQ8VMt2zQW0hxpm+vQIQvquVumN6kAui52p5LlvJpaVZqoTbfRz1lE6KnkySB/
P4qyo2SAXwxNCV4Gr9IkZEkTa9JY66PGSu3m8pvxIFI5itEbWZw/k3Z63anqj5C+
wvxFxYMoyq5cJRYYZNF99YLWI7NNqXxv0B2MIV+PelV+z7m30VEHJV6pxmRTZUlf
FFM0vZh0xlJSoHo6oJVcocAF2uBEZ8Z2gJsKw5mWIaRTv00yEPv4l0RxoMHecfeN
LJNX10knuXMTRio3K+ngS0KopDJZckNEaO8xGxC6fVF1Aoo8mc4oYKxk5scsWgrO
/8J/r91D/Q9q1TNwUQ24CO9PMMpPrqvLFfg4U3c7f6ay7T1rVL0nNpSmVhouYMzA
JU7LkDX1ldSt73EMsxPbdwrG4OP+DMH8yLzmmJgM62q7nAZPwfr3FIt63kAwzdrl
CHFICGnniIYRrgqV1A2ds6VowHOB+hT4BDyYMDoRSDFzSuFDMybUDQNfgHkLvPaX
GT+JHzSDOHCC4pGpIy9Lmv1wz4m6pofnn8D6BT7/9UfU50STSw6B+Wroe45krklW
NJczQWuT7bXIYMIhDcP9wii/6t7DOjKXXSRpwiM7Ypw1m2obUpYKWpgTO++pgqeF
G3MJpT5q/1Kqa2QEVOcIyw==
`pragma protect end_protected
