`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eexVztt/duIMnM3a6s95t69ShxgZiButyCDsUYnbhqvQ9iMEvULTK7i7y6Sj2CY6
vQ/34ttm/+mXCAYA8GIQSZuYpuOXL/MzifZCKVBsw35oCinarxjPfcvIE2t+S9tN
zSz8fPKJbs1a87xOwMCLCDLl8OnSgh4QxRtXqp++XEA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3472)
Sp8tUeCQJ7QlIp6uLiBu3qH5KPMi5CETx5PXIPKRmvEq4s1ra0m2rv5QghIsk2sW
1hh8D6ydRxdEjptbxPCE9cWcOTXBBLOk73Wq9j//nl+UeG3FZjxai3IXduUzMINc
l3xL51fWODhJ3cOlSlsuTp0xkFv+8mIdimoIRNYyyolJpHbYjd2LXrgZonIloaGt
9KqK0JTQUcBcOJIo9QiDAWe5NFSBjafFWNB3zJSMVkPiP7T8kxGzagkgXS843jsU
R6tFGSSi/1FyNBQYxEt5w6gTwCL4k6wzH8ARNYsVipaphdg/pZmKmaOTzgExvWrP
b0eiVC79Ge2ncNDG1ULp4bvRHsAhQ64WmPoy+joFT+sGS9yjQ2YRcEWP5M3PCK44
K9gU7TfXG2c3T+WKrIINLlZcDLx7KQBgV3KnlaGrVfQZOockvlRQd+dg5Sp7c4jn
kzT8XL1TZtkaqDXtSScBTSSk2hfQyW8w2fz835vNwbjqHkWFeLzfWU6IXZV8X2gj
2eUd7mXt+4zxdsqbF84KTWy0J2iGG2fZJiU9aN1B4mySqKykIXxvBL/5lGaX7gI1
wNeHF0VHktjhxBpPZlQpisRB+uMfqA/0wDyz9LN9MuMDBNazZWYEt7I7SftyeHd2
3+/+0YeciXXZDSF+BPw9JVilouJIy8Goni9o8x8CtNmhm3Xb1AQU8R2XtYe6Wcf3
oRCNPbo268NglgYVSYKbORq9KwvBYELhlUANdcELed3OyRVaoobZOs/Gaq/BtJ8P
KBpL9hxieVVvf0jZJqYuhr6M52YfuPMS7ZDuLxkboUL5RtBNFqiCHMeGYrjKDJno
yVyR9N+Bjo1N4V8SJfMxtFWdibcWgiJFzgSZja5AC2WqI+ZPS0GDjjt8X75AAeTi
9NOvSocas2tHzl66hqEuMUb0g84rv3+XGepg418UCxz7PC0Q/W8/J+Jfz97bAJDr
3Me5K6g+EtaUFfgTUzXmRf+oOcYlosa5nJHxyYivtFdiuNGSnYhRYUy1FFwkj0Oa
MbSQ+74edT4ydO6tDMYY9hPrGjQOVdvenIMjGK9lqxIgNVgOeSz7MpkviDjE07Kr
j/dgDxvCx9H83MAFoyM27TtBo9MlemxqJKg0BSbfYzeHBbw2YOD/4Mr6tzIG71h+
C5Xp7THhRpK9XssY1x+PA2jOTFuuHmvNqPn3oNibNUjUj9COC7/mnhJoEMQ8zE/k
89jcvf2tid1khMgGeLipJ+tw9heynlYk04s7YJgcWmJoM/34S0qNiFvzj/MH4VRc
aaeditAuJ3rQqN5G19PjlQhwTT7ETCYDbCbSfx7/TOxrW1Tr/qJZVrYtJXQZCAyL
RS7Mm6CwBqshvHcS0mOWzi6sJS7FaOUWZnsRc7aldo0KtVn1NrGHjmlu57q0zNsu
RhKR0P+XecxHIDQpodUMEuKVRfMDCJ/3htprnXQx9cBBRZAShZgbVSLHzOZFhnC6
6ZYp0PxYsW7OH22w35g9cfux/iyOQArvvbMGzIwiq30qiSPVq8JdrV7NVudlR3yY
6HyV5pgLtdwVEZCytWiz1S2wnZf7Hwb+h4uRZgin4GEJr7hdFgUdEsD2YhB+CLTD
xbWtl+KTozvxi/u0mYnezGTlyeoR6QM47vLgO612eB1ykYrVsKlEm4Aw787LmrPz
194Myd5xhZNF0SkFnm0fS0Z7UGA+UQ5yz6SH5RnQJZs4NXR1E9rWbzI+nNMxBJ6l
KCJyPtsZH7NXwdpU6BIy/gHFYaWyg9lWzGCl2zVfIVqFIkCuT0IE6c2xtN4GJDMP
SH8HZK8fN9+ciOOaxETZEOC7hgZLK7Zn0WNnnUOahFUZZrrNkMssvI4wLm0z1qJe
5g/QLoFISwlYh6xF8SXp96IA8RzN0UOFd9G/1dzXTXof9tlLpDAfaW38op6DuMe2
N19+sJrwWCo+tyOjdU9kgR+AaLwgCnO6HzEojlFATbcOQ9eYxL0GJq/XM3/aYBrR
eKKZdnAcORROekQb1lfH1TV66O4hEx5XWrQ6g+91SVhmbnbs5h2fpd318iyupE08
ewm/Qu/A9JDBPeLUbKjoBOyG/CSPCwWO1wJ8GJUcDf972C8z/7lnHEdEUuI7P6C8
ybCrlRe3Gv8DpRzNkEx9Gtzave/zKVi/jN0C04R9lGeCiLv0BQBjpUMjIOzvfqkX
aYcKwkjLMh3tjXQ4/J9np8gckR1++xEh0kSUkQlcLunEzN58rlfxK52el7UNT/T8
j/yb6cnfz1Yb+AGkAn7GLfvUpdQE1fT8Ku0JtbMyW1HGGgrcmf7ZmrtO4mB+14lg
ZcoYNpXhyqcW8cdYgVjYFADRloopa56zawfI04pvwCdrRwVkE0rUQvyFWzZxBFdJ
r4T8NhNY2P+mJVM8Tae4Q/i2Z8Yx6nYxjnbF7EaJy7IsqLH9xqtPui07F3XeG02o
DcLWsI8rQeIJvTIVSgL+4jvzd/v29TnyXokQzsJIDbScwVvA/t/0L8LzbCb+AkGY
EHR+aXNOEb9qBdOOg37h4QjJh7fhSiiayRdLn7FkWxsIgYkzGAH5cv3c8VjBbLwY
SCtPl5nJqb90U1NuLIJp2M8XJUffHGpsBkTRZAXwP9e/JCHeHHxUDmNLyBfKp39M
PE68fVB/nnvOd8i9iOKuvrcrOZmL/7DLk2PE4TFJE6DRWdJIvgua55KiJWP3vJBA
wH5ixvKE49kl3Q501mUwiXYdkiluXRkZnf0K/74WeNbtdRNQjSiZmsolgdNC/lwL
HqDIXICyNEg+DsXMBOFyTU4hI5FhffGEJme/fdiZgKYG/6HLy/+McYr7Q0czACZY
io4VCnuRRxv0ovCcYsDC0bQmyDCbkyjNKbuXFlYhVxCf2DkZzWxVpO7Zud+uQZMu
bKLm3M4LSnkfqSbEtoyDwIY9jR+L+4+4MJkJTUfh5k9MyqmImk7tNs5bhBkmRSnR
NAGOZzWMEonsIZtBs08hHbxQPVEalUDsxOniEaL6B+onNh1mq7M+HpKNZSDaauvx
pCOecisakdSGUMc34UCwe3RhAhtBl7CL5M89CC6hkH+YWhHNvPCMPcuUD6vFRqsE
Yxy4JQaN1JnNQnhD21MFfg/+idEVplNqhv5oeQzIehC4PLdk5qGGAXHVKBXaVtiP
wqiTeDhoRVZEppZOFlfWEl1gpdUgQWsHi/mp5eyIDARX5wCvp9WXD2UIiWy0MNcA
rFIyDUVhkj+DjfCpjIp4+SSBFr3B/LzbaD1AGM+cHTUbLC8KAYRJEDkmpNPNcU49
FgYtsv3H2IWQimwImsP/DQger1tUbWjNwEptMpChFQYWwm8IuBP7cKFKE7/OjRtf
cqVZ6KwFUAoOOjVT9JpiRDQ2iNFRCKEAXpHDVuW7mVhBA03XU+K95uT+HrZzdD7g
wg8IuqzUhM787jj9t9v3GIj8iJarXS67VoIC0K1d5fT8X242lJfAAkwlTlkdVroM
Ze5J4O5KLwMiSCN8ipNYSVUG7WCLN+ZSm2zrcLeUaAlp0aQGylKCs0rJH+0fUuIK
WB6NGnhOPo2OnyE0dSxQdkGLLHfPbCf/5pn/iwfB4RLs0uHZw4zhzoXEoMbeuubL
vw0ic8iH+g/baLoqWerTtzGRCGPa3MhMcjUBPD5Bhh8Ci8tNqCP52Is6cjhjTHBE
/LU02WtvMNpPhLsCixY4WN5YFrZDef+BRHtfx70Ck8ZA82cpOjhRIdaI0KkMjteQ
oNx6h1jwdfueoUP/fh58wadcRNwFWyJ+43zwmLQ2TGOVqcQ5N9pv3yjKGQtPuPL8
hhQ3hxcLLW//hzxxwJeoC9jFOiWUhpu9Halw6fDxb/TilH0yVLtoLFANuzudI22m
g7FPsQu1RH6FiDMTeWQnyF7G3kBY0b1twEXaihoZaFQPTgrcai0xi16rEPexpjJg
y6PZIpdOiqdZN6YzJQBYwIplisWNTi0R0MgEsg1mbND8HbC3yOSe+mRAFctcbRHx
tcrylXLWR+DBJxHinQeypiaEbkUoRBqESzQkh6HGWkrJn+YgsiAzFADTHCEtQOXC
tO8GVR1UAI/Rta1r57nLCsrXWHD4N2A8QB1Mymvi+jvV1KmmUIOH5zUrbL/j4B/l
crXAOryquPtylzZ1vCHb31I1uAvSvFkH2Bs1OhC1A8HWHyOD0Sj0cvpbqL30VBnp
X8dib/B9Q1d21l7FBco0WWUGkBy1bYW1s2d0rANx0MjDGlxbvvzY51b/8wyrlAP2
KEDQsbLXgh/ZvJcKzDPir9jAyUkPUn7aOhGzFQNV8QiD2dFfjpQ/RDCJn0DivQ+e
AKdINvYv/lq1wbje2kaacSn97MAmEOQe7dalGPktyCctbaT+OtAkeVCOoDIFs5+o
cqCLYDUoWhMK1yfvODf+SKR3GdBhXr+OSwZeLZw3CDx27Ec6+r3LqdrS4H+4GDy1
kz2NA0NoTLm2/QZhnDiZBG6UGwNW+0qn4X0c8m6Qk2kEZZIt2+WaasbsxU3q8ThA
Q03BBEPlJTXdrSGsChDCuyK5kdSFjt4+uTwj8l9WvykVooOuF/V52laXqbXaBuvZ
VvG8s5wB/Mr4G5k6nFbLgn4/A3LG+sspz+lt88u157JKVkaMl5V6O8IBPbrXehf2
ceR57mDNUZVocM22rewc6w==
`pragma protect end_protected
