`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NtFfz21j9WSpxS2qC/o18KK1t26RNYh6/VVuvI5BRy0zijQsIJRbW/B/ZRMYAqwW
+0OziCMpQdoIsyymuPP7yV/mBKDCa04B7p+t9zAxzTIpRNSoSGRNH5oFdWGd4NHR
mitCGa0AlC5kO+2tv9LzJhMLOWlZAauJsuvSkdgKOBA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18000)
PJLUKhGb533inGVTJ4m1JLjWdZtkh51aU9SssOUy9U2gUtl8E2cleLONW/npHgNU
Ppd91cFAwZOy1cB3DPfKN2KpVmmK6aH897IewYi87dVXCVhyKt360bCZLeXJ3M9k
Faq3RyM79Wy5805F2YLjembN4WaWkEBuIG+Nvct+fU1a/Q8ops80vo+VQJ+Ktuj2
TnLNJLlA0ymyJjoRyocvt7VATTeVOycOxHkAlYoVRNnjcdGUrWc4aMlMMAXuC4VO
QGR4y8F9BFum5VfrZEmk2QW5cdDzL0/IM5Yw6sM0Xo3QWKjC68O52nFPt0iX2011
50ky7c7Hz/G/uF0gliMJSrMa6qHyT6DhMUf4X+x2uxY/Nq3aJODr74Gge6CTSbuU
5oEqiaVYnhzK/2E6+GUFiN/GYX4fUSu76m+mCkCrXB1Lsz+sQ4ZiEWL97eEyFQId
6Txr8rExiekfER9JgGwcrcqnUhaj3dxnYR1/Dsi4U8k9rTNJWMZ64Dm3JjRPz6en
HVS4p5H/wCU2pFugJrlzmBcP/IQAWzwaL+opAlAMq9K4403V08GTSQS+sEsmyQvd
dV9KGhTHnTrsdu7anwP7NHkywtbdZ1trSVKxSSpFy2lVb7f2aJ4RdCUT3qXg5S/8
r2tnp3ikgpVAV4cyOntYzRTN5Gi1BYo8J7cG7fzog8mwpATCXtuchvOPbXaTNFMG
2t5Z6LXaTHITuUBaauhdYAx/4PLpQDti3QSlE8jotAhzamLoiaJbSzgBptpbT6Mx
JjCYvLkg+Qdj+Zskv3udOWRd3CIh6OySFk8yMIpo38Nlg0tDwp/4JeRrOaGPPP/9
CG3qoa8Ey+eYQhj3oCzF2qm2f8VH1SwvRzr20IS1bYthunz+a3W6mwRzt4vmMB08
y4XTuvCBUeRmpRyZa++DTxBcRlDw3/SK+PyiHMzgI/4durLPuN53zlCFFxjClgbx
IfrPek2D60k0gH++FQpkn9D9jw54BI0jNROifJekzysJTmD7WSDr2mCv89UuR2mf
EBghUTrc7my26vpJiJWjPbj/6vom7MN3oCHCItYTJ6ydfl0r6cXzjj1WG7O9V28I
CNleJevH3Hc2w0A71MmvnqzUaLCJTOW9T9pVKaSYl517W+ZV65avnSQUK8J8JwJq
McPx5I8J2/QJPEjO86xWJ8iio8VGYjwQSh78+dt0piMfpfq3aeg7YFDyvf/35Euf
EpXDAJHyKTzxQcz4DCfoXzLclRlDPExhuGvL4yMHuFMsk7lEWUOnQLo9wh98aWOL
RH5VGry42y2RYvf1SnPf4Jhcg6oNn3Ak/cRle5Nuqb24V2KgpKfyIjwU/ZmE+0z6
AEbChdOuKX/U8sc9ShUh3X6w7gbGWO6eUfLJZTGhP5IHaY6B+a94C3ivz1DlFa9y
o8teizEsUDGOaxNjkqmD/rtCIWRR3hr+fmGOFbKy6AGKOtFof1ns2G4ClNnlB/LE
Q+ReQ9rhS0pr4gsx7F8Mubpk/UzbSnWm+X733jicFZOojiAjYoCTtSVYy69BR4Ya
qQcWtTGf3azGkA+g75A1x0k806fq+kUFFOcImuwFivPxMy5jZ3Xfdfcs2U2dzWT2
oaV1PQAtSU0rMbmjvnSJ7nKycCBU5Vi6oWOraVgORhen8f9BoTQCxsVe0IycXYH1
fTNOMuPDbxQy7n17CUNmkamzpbM3EKsNjWnU0DlqJTFAkQTX+SLIXZNpImvYxoAR
3YjvUN/7//uARHUfHlZLSdn86XL2Dv+6bokyBvr7CS3CO+n71Uhs03e2sHxm59FV
XnJjlJJb8v/r0HmA9a8udU/14VsBW/M9Sqy7ctdr09aLIbV3t2T/BKJFoPh16PIO
aSgxw7MzvWAvQxSPx4nzzL71xZicz3l9IUGFfhwYXJHaL7Ol6ga8DutugQQFAtUc
VMplG8FCr8B9yUjjz6z+4fyURaUNwPygmHM7lAXF/lTl7EeOf+O6FGFiWa30k4NQ
trhJh5FsPeD/b4wKCdzPi18qtnM5TyEWI4djc1Fr/J2K1G4XK38xzcKJdC63exwU
9CdyohExK0Wtv1D83jMKItUpZ80L1DaFVB8XSd6pLBW4Mq/BMP1RLbkEWevsVaDb
E/MQfhPXhEk97abT80u82nO0P6vovVmpweknO/hNan07LrI2wtqOdBSfXcMstUHl
c4utJRGPQvejRJqh/080I5EB9TtC29cBXwOUHOBOt6lhr402cj9pUjGQuhqUtTN0
DYVNaS2jBTzeqwk2IYAinPneMNOuSLIEFQK0Rv1S98PubJq8OjeyqQJmJ0NsZJYD
6jhffIrhSlSDbBnM+dBoUSgBIBi15fD0Kk0RP4rqeRWnUgyhWyLu2DHcYFVoHJ53
b88qDnW+BmZImxhfhjshQWvLiD9mWKDhB+1P6k/cQLinWjtae/D8EEaZjdRd4R8Z
KZBDCo71PEnZwOnHt6zA9z+W8+/9oezd/tSY9U4lJBq+kuUJ+nAJ0zT3RxkNUubG
ZztrlIv2Xh9bpXaLm27M/zZuSdTIomipIu2jXgfHBSvpi9qHw8vYHPh2c4Rl/zb0
/6wrpa0mfwc2W2U+4f3OGxTIxa8ho8AYljT98e6uUePUpRHT0z1pB1Kensagzlni
6p2++nH4SrrOR1lsha1ClHhJkQuKFr9emiq3j/x2l4AQucBEp+m4uJ8hFAS4TcET
M91k/FUwmm6Mh9p8iEfG0NlUiCVXsoP447HvsBsfFGk5kIf7WYg99etN0bjC2OiR
PNEpmNy7O88RNxcZt4UF09nQ0D7o/BL45egVn/CToxsbMOmsnrvKNvjvWe5dqEIW
7wS7LbpLfQ3vawj8Z135+fXt5YN+ANvZVUfMab3XfnWnIwR03SEUAs/nVrctTBCe
o0Aq/HBzfZcMPUbMdpGOttOpkR/Rve8Myvo7ceVgOPgypFNnLuNdU2PM5DssS8rm
Au5QsWowACTXZZUuKQQhmJaj7k/Z1j8W6VpV4BvDCJQSNPJ86nbNy3yuFrByyEMt
ZH9h+MSURDwrnbeuFOYw19ugoSr0GnDJaPrM7qI7wQjWGdnhZDEHGFGqxpmXQr+d
n/5RmAvK8U2z6vduXTA2B/gqN6kxdTL9KOH3Nb96NYrVmr4LUIcxc23FbU0dzUr8
NfI+I2AIB6olrORB3NDkAVLaFQFKZc1rfSVT+8+bKJiRKQ6Nc56v1n3PH28WL1cL
9puo5syVFF4970ZtlsPjsK+FddJuubvXBKdHa/SgFwAB+DR+0t4Ancv1rkPcDaIS
ocr4CYM1VKWt22DOmqou+uobzg4XuDg+VVBJ+8IKiFenZLn7/pTWS9D7/aV1q1+V
SXGHi2CKoVSeagtHM2qnY60v199z+rhIbaocnqQueQ4m3AlWLH9iVX5RNOhATbB+
EUDqnBQeAVQVRXB4UnIXxeOsgQ2j2Bw/8yeBprqghJKYcWvXeeuG1b5DPSMJXR7I
bE9G6HCQYWIAxvzwCaSB4eV16dnc9KF4vXIodVKnLyzw3XayFMiDVW777E8M2WQe
M+WquD4x9+3rQKuIGqoIc4FHlYa+jv/pgYBuwBCc1TXoZwC7VgAzfWVHcS30EcaJ
voLWJfCOYwMyBfiJ4h4OftQqEWsDAvLL9P7g4Egfh9TMFBuHnMj0JSxPuXXqonPQ
0UqI32Qs+ABGr1xEsqyvKSmDJHOz7BZDTIEnybOOkHW4SdI2io/QA8v0hw93pAIC
5hrHvOkVrS4WbUPkMmU+Z91SF6r61+yTcZUwGqW++qUm/HBVQ18lfpdakI8zlFE1
4TENnYjQHWZCcmvA9YoJaE/KaMDY2lRmwEmXizLCVqX50Z6LgbMSZRpWZCBUz5s4
fayMWDBeDNRAs8H9m95j558DuUcfgJmCc8qc7fXyxN3O6rUJSTO84t70dWlsQ7dm
Vs8docBKHzL4G01ZKIG5V1tFhB51MHZpA4bjoT5eNrMMB+Tgu6tjsVgRcLmUcxw1
wtqCI1lS41qAn0Tv0sYEcyDc1/zE0FM68BPGvo/iEHq2k0fXWh/xzIfXi14nJEBD
J/1oa+8Y21SWeVZmXVlQGoYLsn0tc0b4YXTY+7jclDwuIdhfEAIeKAD7MFO91+nS
hP1Sc6j3/m0EXERUN6BKAsfEKx2/RAICikEgkWCT+CkWUYlbMyucDVSiW2euS/Fa
zvl5epc3dEodZm31nCMjwz2QafC5tNcJWHaYRqcGidj1fkAZazbE7H5OlF7EpyBB
0AFneENUiFxVUCezAsKyOFjXAz4nSKV27vUCSKmrrjkhXo8cQYcDLkFjhTIcNjnY
WywZ3yQUNVOovX7FSsnEaZ3EsozmKVUzHi/OfI271+9d0cnEDQB+E2Ih8CRgH1nC
U6RGcwiPXKgo6ZPkQv8w/npU5OyJjz+a1iv0d3I+gtuUGARHocewp0hT6caDwGfx
dh7jdHeJ6a1tHJ0JtnbQq8Qk+mbJz2rPrmfEMIOid1opxn7MKbaQBXa3SnGZw/hL
YWsdfsi0Ed/eafu6Hvu9SNGfUDBCXg9J4uvvOLv45hNr4jlfP9JA58suVFy1yl+p
8YLtA1HbHLi2TDS6u0tBO99v1Le75kRR0euXHdLyDJ1aQjM1GqEYOVr+vMegbVS4
+7NamENkB2Ae4+19CQY6bG/ypZ4SJD8k9n7y3hHNyfnXX1PcdaLZfDNcsLCVMcWl
LBTRSayFcQRWILoh9YjPSBrIAZW/97+ocDhl6efFGTyCBG1GBurfGzTmnpgqt3Pu
jfFDF7/8ap5naDmlSCXF7CYIv/e7G0kpioe3hrZ1UUZ63jR08RZZe28GeFYre/lm
fx4wfem8R+Txi2N27PUpi68577Dp02S6nl6FZo6plFUCnftq/BNQVqvt2X/FDCMz
B1vYZtQZfKOfkIBapWGZkoikkIsjD4dlxxCU5DuHxkWKZ8TA3YmUcibJOOa5A7sM
irNHQXQLJFmijhr4qgxRQUMg53f6Rh105UVmfb9YHLUPmLCgua/ufJQzkMEZ/4BK
jTg8W/898cH2NqHhWjXykGPZ3ts4XpRcFAFi4CtbRAG5A/ZF8RtJISaZHAV7T6GQ
H4qDikQtTouB3M8FWRNN6b5GY8aieG8KUQZdUwORa9sPMaSCCr1EFpbVmeugXIgE
Q8WnmcziOYbB8BOmPm7El15WbYAy/F9+pQ9iPQwn5ND+XNwaXhRnl7I4gK76YyAO
AoyKY0ix5nuricJlBizz4OeI+YZmZKFu1aqNBRePpnANoaX38cvjnt2hEUjFD+/x
Dpgrf8B+BgSZV+uXx1Td0WR2yvMf4dpj6S86yNugJ4kwgIlxX/5IGEzHkS2hMZTQ
132p5ES9Sz4eatfNHM9+QwmQX+rKRrhQSe53CK8MlFIgXtwXCsYwHt9qUI5fi9dl
WNLlfh/G3X1H2zuTYzyPrsvGrM0VhN+dDJOQXaNXhYyZwSaa2nI9R48XEhZLZmsl
4xC/jipAz+Aun4V2auiSkZneq1ZCNPbJGsW9DDlTLCibqzoET8qbqZ/BO/jrXb+a
IT2Ksr3MZw3r2QENY4NT7XfoUmherhyW4IRrhlZE3+zAj2QDdzJ3H7/hZjlPKErO
4cdSxVVAgnntIsyI4mxJ0K2kJkG4lD6hFIOaRpdBdsKRvPejLvjC0g4zqCwFY8+n
8klrBoBCnRLorElKRdzjEdfLahaDJlErVhT/6gBXcr6YV2WFTMIDQv8qHsdpyWoM
6LvVlUmJJP/NQtBeW7/nPYEmxhwmfsuOsVVOkxGPRQS2q5FanY2QdFj/lPw9yUAN
sBKelQ9mB59w3hy/TB5T/74p2mvhGPNnWUSlEQSyetkmp+cgBNvI8xEgR99kT+Pw
VaA9GUIpBhPTo8vhPQGzmNdCk7roUe5PP5r875wFjI7qtgG/llTVbZPSriB+6eVe
uCYs5C+6pKfSPhxG4hiwsRnb8mjhFIc+ts3JLrXV7WjiURJOQ5+o6IMgLgOQDWcw
TTkXl/bvsR5Cyb03BIQsnT14gy8EfYakLdsR889MiigqJUl05ViEKoKBkP1JjOvA
ZzdEHdgRWwjwwJFBi2w5YZu0ZfWXM+Me6aUvjdBChfE9tmH0Wxb0Vl32qYzxDnJ+
i595jjwSoGRfWcEJ4FbqIGg37wyU8gTBgiWgKMrdx3BB2MV0XvT4hX8Xm88TOEyq
RSCPV4a9Rfv4XMBLFinIq2JQEWwK84c3v4XHUQhj83duhkeyJJDQOE+4XBQGZRzD
viR0miD5yyC0SaQr2HPuc7Ya7RAGphqPsMrDEl/d3N4+nLY+XIbSzhcetxJCPFLU
vNwdbfo5jiKDBDoHNA1vZ+hE4nMIg1CSWhv7IqZZQEVv4cnLK8uLUbeJI4OwsRr4
aBfesRAmPlgVVD+eAxED7GxrQg/ZAL4mzs0Xx/WE0Zoy8O302qruRgoQn7JOz0RL
FSD4bTIpFBOK8e2ExyQqMEnE8b0jNte5VEzhgz/sohOxGppTZMlh9nIdiy4tVCZA
tGZ/7pkZRdtVGnPgpvDtFSG3S4XXRpI2C5efOVo9ILnMhOI6fxUDgRL/8oU8fEOq
G4UT9eygK9l0qudqGq/WVzMpBT2SV43KsK4G4D0xmmKd+IZ3xfnodOWCwvJhLKyx
oyQqQ/HwOgge+BhLYSXBDZr8yGb+2ztgXTRYyVR4ue8NS40NSgXlyjiRRAA6SygP
vGDj5R5abs/3S0J7NPt36Vm8R3S8a5gO+55KPCC5Ek0oTmuxY6t9hdsQe8xTTKhW
cIXW7mi4havu1uLUCJPQh0I4wuzX4CD8fmxh/z5Gt0nad+efDQX0PXk1+GgGJ+nP
mSfQ5jW7QgTBqR1qKicupHurPC/NvzDyti8R2tts82UYWssQzSrAHm/DDljoN/Qo
6Jkt5Zyh+KcieSR4soW0HYzL9g5IS14pnPudlZnvm72On5q76g0OeF4wERNkccaM
VCn6gvg4Cji7jkDjFZPCfm8cZLH32RNzvDvV/LHNSUnTAe1UwHPoozlbyPDHpdsN
7dgnVMhqI8dJonT/cCN4fb+HpNPr7hnZALaoGUj5MEOOA07vRFFJOWaf3KkEwYwa
8YbYinT2Y0K757LL03YaGzm0f8FqNH8+pXeddIY5HQmBfHsa0wVQGeGZrIvK9Flg
4FMhSKvNw3AYsPpdkaSS5gI8QlnkGcUNilKzssblrUutNKPgtSkaVhROnwdUBoTO
2oAw5hqGfeRAjagZsOPRwaVYBWvHoNy8EQisIGca9nQKGNobSFZ8QN/4LgPlkfJ7
DXX0UPjJHqAR9KHmUSQWjSOqNH2yaTfvpMId0w0OsQHVOfVy/pr27+YlDT/3Yi57
sAa0nD3398YZgPQAFUMz6ES9HA7w22rbSLp76TZsTx+VHG9c1y5YwNmxCyWeg8LA
1lw/2xpAaN5/3l9FXEcycmomsBi3JlFdrR2XJcwM5366JPssjfiv1lmC72Oas+W2
7ufOImhxkjPu1vlJaPc2nWw53RRjUnqdaqhV9Z2Q/2TzKjlttEG128quJKwiHFnm
YltE5mSNCrs/nRC/XwLGhgozn5f40B5gLZeWfB9Z2kNH8PApz2502aLSiJ5ylR6d
uB/9I+yAMLDiv+TD8yi/wGVBNfvcl+gQjxIIYAdy0l3+2l68o4qxhHaCyzBS8UcG
icL8NOwQxF7e7ULzoaQqF/cUs/HtX+5dlT4Fx8Do4K8uekKovGvkzupfl75ax8Gp
VgHdHbgK0nIdgITndHBN5kFU6pChaSJHnyTIjqXZ6WAhh3PobAOe5T7hJfZimNr7
JMyklODJNhsKsgMBfaH9dxMpbqeLpXbSzX08kmvQp8ad4HF2rMLz2f7OnuYEp+kT
wTAFEKK/GHA2/flmi/WZs5oreYfTN0/KeNb32FHpnu5r6dwB+f7kChnF5a6JX9qE
tc/EP1R9whYa5WRuw407wyECZfo1Mm5gqLzlEV26F4SbU2O7kPoX2L3+X6hUW06o
fE6jzk35GXGJGsGJtYgHrWfvfPqn9ntWa9F66zuTtpU8r9Ol0KD7X29QDwZE+465
dh+crZwo+Yfx66mRD/9/TbaFMUwLYV1Tr6l5gu89mVg9C8wbLsL9AFnCWO6NW2s9
6gBE5LNDywQJTKj7vNbztvxL3tTpwyKsRBH5Z5ER7iaBsT1dgXFLsMSfYYgbY4WW
csSCkuLK6u9rGANMKX6NixRK1zU6GzKRBzaKvFy1c18cJYUSdNry2sJuaFnlTqku
BAnq5/iNBz0V7k+OMRyEF1kYKCeaTL2plBeLglWdHKSB09vuEGwak0X50uzmg4j8
NuAWZZJTdmlypFXOP7ETu7lsfWB5kQ2kPeAZwi2aOaMqyXF86ZeH7NHt5encAxOO
FJZzi+edJGLUALHIdHVCGnA7I8RkF5sR5e4tsVPZkuTfIacgPA3/fgYDzyZdMx3r
hgK2uz8gVr2iXWjkAzG1HJzrC5kd0p/UiqxcBO6bqXX6EwquUnmhn+RK1k0FSzb5
3u0vQ8pTcjNUHfXpr+mdF/A/hDD7Qs1Hv0ZLsmMAVfEJKywJvVW0Sb75QEeNOfv0
5Ih+HRMlEUNSyvCpOECfwB2Rx0TdSfxpV7HJRcnn3mx2EwTd8zEddKyUv36CbGDQ
jEZn0JXctGwaLccozE9zopxdNmEXCleeac+43BpCATgSeSbcV6KGgxePseiLCiBZ
dA6GEKKZp7SUOLPWKpN9YnLxRL8U9Bwn5IelOXz3wf/le6AomCdjQXPkXvGe5scb
siX7yN2u0L4bLyqmcw+W0AePv8/RTIEFu4mLoaT61ZU1SsqgZ8ku9oCeROGZJghe
EjuMeH9s9FN4PgcS1gvloYtoGkDwxfInusmKqhGSQfoByVhImRZc9gGfv6Rs+ViV
86PE5zdcaY5ik9dyuM79MWdBoEICrWfS6C+1ZnuZ+ua6FxjYWpbPBbWGRMoEoj+8
sX04yheRkFMh/wrlExIebktoYV2iQ4k6GKPQSCr2QVvXS2vfuMqHf6o7+zLmQV5s
5TriRTL4VB0xpzwj1pdXZXHuftPN2456zdzWZPA/x7ZdVd3zLWS0AaPbRHL3w+Xr
C52EVD7jFheXInA/FChvPqxzlL4REqdwzNfhJFeRjSAwd0lvVRKtJF2neTzjEmrv
vpGeMarSB38SRz3CCprmgIcRY9iLM1xhD8XneUmWbMUPGX4OMKQRGTyqvGm0tXzM
iXl1Sy+zb1Rl1x+jeY1Zu9L4WPB4KbFFCGI5DA0HG4ne/ZUQ4OfLZ4zoQLrcjiL4
eDEkQIneFomdFohdu9OIW4JasF6cFds4XYfVMuCFa01PuWQIziRNPcHvhA4Z+NdH
r5moGYKU7XHHWmJwid1t5YkspdVOdhf46/5bvLMgXvc3kMT/F2uMJn/iiZ2xJddh
5uF3NKuNI5U64TngupoOZIUWw53ENXkDuFlNCNZGbiuR1FXZ7Y+kJ1MibqelQNzS
71nzgIscjnDHimOfR7kJXemXnoSFnm8Oxn03OcQLaMIdAx08x8G7dXFrlKS1MFM7
VO/X9RbHf1kDoiETEgSPIXT5/nrZhkR11f4ZeIlh3NeE2QAyqoFNoBQ/U7pFMJc+
4jrQHqGelGc/pVy6b3o3j0OOMka8ULDnLJkoMXDLQv3EEsZp+/099NNUfhdfiVBu
SQ6PWMVAHneb+GV9CM00IQ0liuEESluS2RCrpZFtCrIbNWtosugYMiffOZXIei4w
Fz3S84PeNaA9RVLWy+wXvL4nc2+u4VlgJQzjPFkw4qvgvtVsYdZc94686GzYZCIZ
py1ntaXhCpN9fBV1LThaVSvRWARBhBbcPJchKufKg4zk5ssct52pf70aJKrsVwpJ
7DtSiPxxvuaAVmnzR8HDsy6Yc6yUSdgH0gg1qiUH5D8ARddlfezJiRHDWLVKkXkE
B3JQdvbpj4DtZptiQ60Pmdlz2HNQvrf3/rEiYaXdZDSb5sx+5seSrXY/kHECOAJ8
FjWvP+E4OdjaMe/VDsCdHDsLz6dXTLKlZxWzi31METvap23ozAVZnRhQBRhC1qgW
8L7SHvPo2KZlohfQxp0+kRAgiSEOLZg9aKJX2CLHtvRi8JrsZxdyjPrkd/syjhJ2
6x8t9WcxdQEMSK7y8j2DYhR//7UuiDUkQzfNt37hwSmwQV1mYiMz4N3yK2A1SZiC
s1/CZsmC99xJn/eu8AFC3Xpo/V0754Z3+++opKtPyRTRs0tGdqnbPlqzCJEO2+h7
cA0vHKb/TiWbI0KBx5tjuWZv14cxiQeJzd6RWa8EqmcJMt9mX3fPX61q52JCOUVJ
Yojz2pK13ZwSDfxWLH0E/vr3ZWEXbO9Fj+6dKzhTZFCR7K+i9Cn44+7NNk2FnCki
0TiUUVsI3hQFWLYbPaIld9/Zmbh80Iynlq1pBPAeVgwyKO8uGxYngfqzwXdRlefX
XwfrqcUce3IjsqUoUyO7lGHETQPbeLzhP1iiZFyLODKklWDEM0cIvROmlqj10Xe5
TCZ+Ya41zJNWpI26rAHe1Z0dVSmFrqkct4USGynlylLI5EEEyLiVzkhrl0igap6g
bHc0gWRg10iSLvRsueeSJQW1Q/hChEx8fDSrwFzZkaVcdWQ77j7u1ysSyGhHZxap
7m/nDUuEwvpiIC3DytVTRQgwE24K8Emq7rtXmpGeIJLSaVKy7OiKg8H2us4doLDs
dWy6osQDKTe9riFm86IB5NoCgbWsbz2yvs7H1HRohg6Lu/4sMKAZKQ7TxSNl0tZt
HsySXNExSp196reHiJ6tE0mgGmwMBtGOTLAfCjim2i12sNwGiGUxvBK83jdwkZn6
yGWoXWGhTo13NzcnXbRgPbeyxnPQ0/Y1l01IDQim4/MmQwt1pzotp+0/KC5kKLN+
ebMJlPrMgI9jhrNyz1sf909wg05UDNzh6dhT3nYIAMIcht5bCH/oWjjp9z1YwLwL
pARF3oMhlygEUXEA2ZOLOeK2atHrkFslmAhS0RJJqK3tmxQ8P3id0Sdhv7jO69jZ
mprlxPXcm8o6HrbxgRPZjRVsrFjZ/D/y6tPaVTQJpw9j/ZxESomdWYwQXRvQ7nys
TTnprIOky5a3zkMQL05zuM2Oju9cuuGkl6E2CsV2f6xfeH/+IQe35i4JVYhJmp52
f6HDyu/hTKHEn7qxmq1bOqqUZ6Zvub5hWtgVU9K/adaMwxu2Fu5H2WEyFf4TrqpO
mZsnCMXKfferhVf/2qop4MGucdbI17/buQRNAtlh8BtIGD6zGTI+gBdKQaP9GGzl
4w7D5KrTypvDhNDfD6kSZYqwo8x/vQDSonSv546WKsCsa9PFoPCaomXUkLj9fJkw
qEf2w9DqYOpIRYIptJum0mUyMglACzWMtsw4J15Lp/lAL9X9atsgSZQTjCpZEnW7
hB0L8fulKdYexFA7MUYqwLDWBgB37DYdq+7NWjMiDEzY0wHs4bKze+ueuSBaV76b
+1gDLDTI2b1COrUcZNAAs+eqUofxlBW3WZqVPwev98iQXGZsZkXM9U4pLlIF9se8
WQulgQV476nD4KknVmUbdJ+O+z0619+i7epyJEiSKSoVAI67lquIncMgWv4qO6Zu
jF4ANQ88cIB9UQdG4r9Ptni3JUQ1r5LiXb0adUhfTcs9zvV9u3BRFFbV7p1AFrmM
fPTGk1rZBPO3JdGLf8LkMYsdv+Nvp/ZrwSsF1vdpil+fdgvBvukyjPx9yW2Xfqw9
Rp3H0vcghGtfz9NYN2hPDfxAt4nDeLpTYRv0UPq4WBOLWS6gFAz1n2xRkU/x3O5t
/64qOdg2MZQ+mghbPnwB+9537jGOzZcFqUeflU1N/WMvagObhui1iw2RkCSlUTC6
zghVKcVeiHPqMyRUFVe/XiH1LR6TI1LcLX4cMpwYu2QzjerJ454JI4kXjYxFK5YV
iO/kdKtYIq/sAiKJcFlVV+RRWjIeLGbswT10Y5b68vUivUJpXQAb+JIfpxgUtL7l
/p525cPlYuEWwwPLfALZkC5rXmgTDz7dkfFP9mAuHEW+KWH/dAsLEQp2VUQGBaNW
IYmoobLdPJgopWhGH9Pj7cm9s6WrFOdsyYdPK7fCRiTnWF1Eof8BzEMukjTB3t+P
+lOO/mL3WfiGtVzyDwdAK/VF1ytIR9g2q3k1r6JFPxTS8yL+iWwOoGnmkunObLwk
+sM7kKn90TeUqtGCxJB5bmEof8ViauxATMbA1c1kCttzgUOLiXWc5PzipYo2LoDm
QnTZkvrQhzMCGrlK4fqjGqDL/ixXI1gnhw8DVFJ0hBoGvvQ1AlphxSBASz9GCZml
6KpjZ1GCXye1NVJN/iqmZUNNsf7Kn8TNkzwrbIunFmA8QjETxqLmhNuok6vULR38
6jg2HgKXHz4GW8IBG6VcKg9Ie2PjLhMTFJObrlVAPid2bKIc8uHpDi9l4oezBYaH
4hXOxUSNEuQ0JlIW/HZELupdT23nZvxiee8RmH75bSuqeMUxcIuszLTph4OvdIP2
KN8uuduoQf+wlxWrvIU91MSWP9oakkzeOTH0jeOBR+/G1bRlzA9cpgxa+i5B9aty
PfI/hSPpg4ARbY0/deqZ8J7aX03sZ4n99ghmsDBL7FTAo7xVfWRpxjjbvm05C/3w
IqeJvSrTturQEXXld9bnEd0i4oZ3EjVaDXnYzZIJnrG3TpEZ2HbiXeNNAmFnqUy0
wbQ/1pB5VGWUF27rHCvBqrfO7e5mO+PbRaL9enUhf6tv1IDanReGQiT7BMvvbYG2
t5dHUONvmH1OmDf6pdEt+wCgKIf44N1Wh0mkz01PyZKhsh/fIjJUlsJbvJIx7vuO
f9+LZNoOBIRMAjNjUDMBlN7IgQa7ix40+ACcnoW8+FVeIEvdvuVdFrH1HRyCKdDg
+dYVYowVghFe7orcC89CRxHg8oaove1y5fOnhvL2uceWoWnRZ4Bnt8PDm3vuLi0S
nUxjc/NSO8xZs71fEqGe6OfjSdBVy3tl9raHNaUUenBwMaYnnMYQzWot9Z8Ibqyu
qepp5kdb5wWmVi8NsEH0/vdQQbTKWpXvMVasty8lmqDwb18oWt+B7vmXhhwFoyc8
zUCpuiRLKb99dYmaqCoYfdg6WQWL5FXzFZpSzywp7KVOK+1ndK7MPkEhyM7cobDP
Cv1AavcjQa7q7ZBXT2iYpsoancJeo3fj7KcwtrcQCStuCDKGU/VI93AldRTmcoiV
XwLs0m0rPhqEMMmbOELrb6IWzKAwsr+aup6m/aWo/UA9ABmQH5UwwKmOCjkWbknM
MQSB9kJcV6FNFlkrUnTC4qIBehQghaA7LOo7jMz2siDP7JCRRuveR/4wF+fsAU4v
UgEDiv4BeKqXT1O3oIadxU4LVTYQh9n0AvUOqaNPu0qHQ7CMXehSHACUHV3CgIsn
etXR0eT8FDXYZwLeZMzPpvojlCcrS08XdhNi+QmrNqEnSzeDwzQKwU9A1QiS/FpV
Zkgfann5kfLzV7OJrT660PLA2GsCtP3zGqBhdzcIM5vItx9wHI7Usx4SseEdy8Aw
IEK1rdIl87qP9Z2J0NpOwilCg7KO9xv6pCl9k81bPONnzRB/vBvqC4CVK53mfWxX
btY/37cq3ZkRhBzRNIvNBmYaKYT5+P+d1b9Pfrlr5SJbBWGpQbejWSsK/HhoUJkd
eH9CMWPDcmnCVmBBrWQrlJinPzN9z8GNyrgNq//+OZV4Qs0dxQftHjYAaXES+vZK
HV0vh0Nl9VfsHixAvqxp8WEY/G2M2Kc2RU6Y787IxxnJMoM55Z2Qz2LGEyZdTICU
10m0/QWy4oGumKsMD1c//plSWLY3vgvJpE/CovYa45Z2HuHvp1hQigEItqxmwPYq
AFV9Yx3nHd2UCzRJf0hujscqhsYJvO/E6VURrSdKKwWXy30h/uoeRJdfQM6T1ocj
uROFGu9MHo77uMQliiHFE230s1dXD1QdiPBki5Og2+9Akg75kxPZBC1z1uXA7+3Y
yjdTaiExJuxyu96wGlqAo8TBazAqLocdQQY4rLQJIsvCvCf/cuy8UtloFuapudXX
BQEX1n+9OHqVL6W923iyuvUXoTtTVxtQ0k2N4h0xjgx8Prn92BZMAYZox5zQylTJ
Dmxq+G/pv1+7NcJDY5LsX/5UEe6v4wlvNyMWP2DbB4YI0FvT22xiLLa1XIPPjD1h
BCAEIDEaRHSs7Z/qJSIW6ySZa4GsCYtlIULNBLaTtY7Adv2igirxFaYlwccX+90q
OpZie5zGXSn2y5zpFFHlsEytM2C2eM7JEpRkrCmJL2quyWhdpAS0BT39PXJeWCXj
oHTrOFuDFYp/lH0Se/6WNFBv1APB/N+XhX0TqVy1FunkhHNatWFZW/vMjw59llr6
FuMX/XX/RMYyG7DT/HX8+MePcdFzPgn0DFnPF/2kr6H0iEYCIDDRIhcBcIglMl5C
A3nm967jBueYGoAk1jrPjduqyTlcK5c5pgmrnOk3BwdaVAFCdh7Db3+B+TmjdHlU
6oT2n3rDyl9RY7GWaF9LyS51/ro3EBc3Wt25g7c+A0XJ1j069+rLqikfFA+rEZP8
qdu93BBgBKEMl+ABAvC1R2I2hlX1005J159gOndzm5OktyZVtQ/tN2eQvafTKDIL
FvBcp7uMwN9/7Zi8nYzcLxY/Ia1eDLQVM6awjVJVgtD8oMNBWmokuqf6GQ2qgXXJ
2kR4I/OuKoLs3PNo/ZfIDXyGCYrUQ8cWlLsSpSqGdr4aRfInsNbmWiAZFgvnNf2B
n7UkucQ2wKaCCoUPKN98l2n+FmL7IkgLbBqhMBaYVGneb6PIsN+JbEGVWn4fAcz3
WnW9FSTu93i47Awx8LZer45jVRgvIw1AaKWhRPVhQXVwdiA9IYlhNrEFBWkJeMIa
E3nhiDkJm7IDwKQkUKZ9CPSVB6pQHqQWQcYfgDcN+RrhjgmGm5jpDZRQmmlYZzny
Qg0HpBkthJitioIEzBy/aG7dvzFdjxWP6s+8HAtYj+fKYR5PV4ikc0CqyMxyLCLS
ZBnOteGG4/mSaqhvruvZj4WsTZJvrfccBgWEg+neemzx7zmn/gXGOaAxAI3NUIGx
pBoiifWjckzYnxooVh7+Jhn2qSmxyg/10cQI9IqYyFJ2DXezraTvUR/GcTrTcPRA
5kEC+0i+Gb9kAG9V4WsD5GEETfw6zeFB+VGxf2RrHLw9KjCiOBrYb5kq85fJth7z
STy3QrdWE40i+q94IpGRXLYz+ByP1HBMajNklL4+SqbbYEIHm9RB3ifcKlAYx4ts
glsw+/K+nSRkcV7WD5fajL7/q1ChOWhJGifgCWo+THIo7S5HmUT5NnckM5qUJGqK
9BKVfpIHyVzk/WC5iBddziWCA9S+QpG3B0yCpcsI+sISeaRJVsu/gxH7A42vm//D
x+Ha1x770jW/bkmWRO2CSUr84fqtcSMnh3IkX0Q1vFw2LxuXllFaHbHs0On4No8P
7EVa/j/d2AGSHENGPBrg7DSxtK1rF/DMsVD4e1ZLyuYH1n91m5RlpvcSgTwBTHYI
XWShB/hnJgaD7I1HUyiO2sAfgsADmt2yz29xD8jnKWBHWewD6H4tv8IO5kfkpSNy
9myTAzU6qT2uHw3Iv9anBjNZDdwgho96p9Du89ql513TFQItM9a4gC+aH4A9571s
zs7dHsxBHHlbN/URBEv1FYauStWL4cw39200KTV2BO6Qlnj1jNOJAbLW4pucDfY/
k+6xGKx68m60l9U9jjvVs45uhhNdBAhZZukPZYuzD9Jo/ey+L9SD2Qs4PmZhD60G
Ft0mTnhNlopSiZwxOpQ8F2QXQ6PrbOcrci8TbNMISlflQNmdiTnA6znoCLqqqpqz
CHNNjDpNq4jzdvD9DYDrqdcWbPU67pp+0yzojqCD7M3uZqu9527kVwQfTCOb+Xjv
EyQwxs/qd6IOzJiQYrCW0cqLbp78+n3w0R6pG5g2TyD6YgQGIXVmncPkQENvj+LC
ZsgBHwr0PY62w9ZAbptglzA9RT31FYoOG1L9eC1waFLjjxu/70gZVG4avR4VunAj
YeN3jvmNGr3DB1rTYg+2xUzaWpGrM9xCcZQdUWEAvBJjN6/zplQ4Spubg4aH5GR4
uGpDx3V8ijQVdMIaX9B7vgwNpuo5e4P+Fl/ZY0/CLvlwLo36qBdYsrp1uTOQH+jZ
yVKDr86M+fwMGwVX3YOi31rJJJ3iCwqk97KsgLJlcZ2rMoJS52DQgTbEaCqz7EJ0
RH6MlzSPb3m+K/j/4uu9gKi/E5i9hSzdXB2/8IDv5m4ZrMvWL/8F11fG+qaZo7Sw
IdxEwmrQInQ88NrJ9grAYaMmBiUIWvn8qhbSPt0JQE6bKQ2Pp3vQVE2gnMXaN9fH
T02x1KLNNBqQixAud0S10Jyvq3k36H5s/H5eqZlXGMG8T/VM3OqLMr88HDYSTdWu
6nwXQnYwp+31eNZ7iu9tlRwy7TzQlucVjQagBYRBVwOSalFnClvKV6V1vw5o0J5A
AfXqIByimA8JzbUx2bvN2n5pvtHX2n6t5KCQbkVtLyTPK67qvZJn/aqyZ0UCfp4b
7bUskfAfzXyX8nhFtyaHZLEU4EV8ICmorl0tHSxwcRwzYNp2lNlvJuZfqBiwWdxY
HBcpSfqwEdXZz0ejMmNsmD8oppTW7cGPT4/SWICCLQ0psoQorFe0nmLzBcIujTGD
+eQowtbPW1KQfjhYUPJtKLPeveyumot/16+M7Owjn6m77VDLYAm+B2Vxg9ZA3Y37
DzRObKLQ1ERDe3b2W/vy6Sx/UoUFevwHshZvxM2ok/vo2FEc7kA5GQHWApOSmo15
64AVYa38c2XulapvhwSw/cgoP8QHFNo2qY4/Q499e8vPR2LRlfvkYnS56J22qKpa
co/jMuFlGL4IFVVcTG8LnEKooSgZ6p6WrbPFIN6HAmlXMIr3lu3/SQ93HHe7Icmo
5E8yDOe6wyVXsEiS+6w5xLww3wVoNM8p6oZjaBCj53qqQN9uYYEzZ8UMok4rsjiL
3FN60fol0byUmwa2HnlzjHRpz2aPGYWPxS7OqPuHNOBOJWLlfVqvXKG6yOwgeieo
CoEyZHtlzjXwDDCmiaD6ASW7czzfz64KgwPOwzP98lJc96HJDZqujrLzqqK52pkp
OEBJYUECJFw69EhK7IAGLhlHkj1xxQ4/VK+IA1Qpuj/94sG8N1Qh8f/9aZuFbTJ4
o9PyPuMvi5EB3+/2T0BHnXHr5rsngORPhcTpPyfY3VFBkyQxSC0Q9arqm43Ldn1a
u1nmsCvTBVgRJWM3Uhv1xG8niLtV8OkomhwdgKK3xD53e6v3pJMbPtrnL7HZjCRM
avaq3w5/43ZdPwZfd3ubUQPjPsu24XjeZCaLe8/i1KwMSn7FVsFfoe4tbYPqOCI6
kihtALwvyCb3411mR+2WyxvjXzPaHKsPOFOZZxdCwkssBBifxqk67M6HhlpryyTn
dE3Cb0Vuf1xWwITFUQMEifXllujUMWEorgVu5iCqpKw0NYeXPVWWMTaxP7PlJoB4
bOp2oaa3ozJAeiVkOwLEKPmKePiJMiDr+SndySalVDEyjiW+8WkwRRdTGrE62YLt
h8tg5OG+1GrVjYLoRSYjJaOns44ZKyvyrHmPiUvh/f2ScAJTaYkDry6Z2mHmLufj
SpLUydv1qqf4kbvParmIt6sWUYmu6Tq4xhXIctOcVt9Cssu9srk51YLmqZxGergS
GYc+mOqaOND2pUD2R3p0zxCrPKWaqELK2XpiY5Aigosa48kI3Z+6ideqjfhfFB0h
N4qTaQL5DsQBYrsAblzLEh6jzja/uWibv15uk3wWy136UV7AN/SVnZcGZinEP57f
SneIXlDukJqRC2tq4tgJcmcp/UkS26F0eRIXjcu1USZ7NULvbTJKylPiR1bVdYxO
kFj4JiUPZUt4RBRklVl5D/FzDofm0ff6PrhAre6YutCwQD0hTfCu+synFc1vdrt5
IOnuE3PDplaCroA2zrMjxEvMXHcSIH4zjBiQVh3RkWCzAaZxwK7Tv3MU4J661gGK
KrspFDOoM+In1wZ5jZVRwyQxogddy1nqRi5rTvy8kiFN9MF9Tfmi1OyaAjQOFrCC
f40e62iwwZBW+tvYcexcf5TJZy602ROzT85kHvD27BhTnIkioQhIYcA0jctW983y
0WCFs2/MUG2LqeA/rYGKzg0vnWq+jL1nqkHCWN8ui4qGdA030jX01yxPF58CodGI
6aTYRrZsOAhH5VAd+CV1ZWyhtXdEcxSsAsubBsmqpCByVJQvA2a6CNU4tJ7il2C4
X0ka7eN4g/5uX/8HIsjn8TQzWfjLnnqX50CyI8TGLFKs+gzZntRMxb/StbFQs5ea
UusnIjWmPEHzc6Y+7ONPEfs48OFZMwe+346yTLEonVBBUFkmt0EkVfeiRKtqiKf0
UOd0WnsXdqStgezQ+CVMXQcTFDH/nnhwo8ZESb26qp4i9hwJ0qvLMR8BZ5k6EyhF
oKtBPvT79cNKy4xAOzI9N0WgVmMqhBcDvA8Fem56orv3F71yGbn7C/KSQK20xioa
nVawQNWDAnmgjbzTb0Tu5aWI4SJUbZt6iTxyGAKZNF0bXNgwQ1SaVPM3seSFdL69
3bCLbl2vxnOiX0NcycfczH8DlxLj6pu4WiPvZS6Yv6XKeevwvX7P5cZYJTvJq5vz
OvPcHFBniV6idTkaEtZeGrzOCg9qNrouoVQyiV+es90A2vFklpqmwk71QVLykoY+
HT292HQN3EjZyFR8f6JeAWq0j++3IevZrx++nMynf7Ug/w8PDMxYaUdntrlS2p5S
cLVbQQF9NWGK/2nQ+RJqc14wQiMCb8T54A6MAeu8O8nwig/8NHXqd5JwusIlgUeH
QHwaAeBzIiDVyJCr7B9sDEmG+XsdBn5IAQNrkcDmaJVmOI4AdT3U3pGVGd15FjqT
66YDkttgzacWvnhCYLqQRmL9QgMxp0HQKYE39zrIGYZsMjxEEDfjzP9/omasdGJd
wzlO97wh+BuJpMJWCyWdNinyd9EEE/c5lh700YAPLy4LpknDV6mbLECTkvJ0WuAZ
lGSQSil5gFY8E5LD3aypLotOOMifi0E0csdtBLzXQNfOpzfoxoDbVYRyryYE0fXm
IDcjzUisk1sHZFWpsJJBK70oAAJeQvBqTgbJcnvOxIo4iYLU/Pm2LcENkBkzDtRF
SQXxTLDt+ZxUSpiccJBoGePxuLD5uW6VxAcGkZaKDBh/bf1LacwSgajn0yx/tuji
JazXa1f5hPZk5R5Mh4sLNp48wM2pXFDHT1nUnbWau2rgMqsN9LCFdjySWHL1FkiA
JpXedO3zGDPMMLzuKd/Flwu2tUXcVGV1JA/xHPb+MCiaoJbocNlS82Q8MRxtSxCb
0QOolJXT2K5WS7Bdpg3J4pqF/ptv2aCsVtekfYFvrVISCLOUY1XnTnnugSheMg35
r14NckIHL/QPA2xIBT7jwlNwFkGEYHGL1sIj0izBuWgMsbfZtWN2YBu663VUWD5s
6Fc0vHdArns2YuU3x8mnwb+NrUcuN3Blgr6SLW8bmkmSpuCmmDr2gDlaJFopLs8S
y3mA4Wvf1jKnDlcInmUpOhK0DOymU9URSwuEpDdyLmJT/dj2hkQxWyta0sfB+F3m
3D68EksMYR/940ZCZNA43d96wJsjoTICkw0cd6Z5wM1uXWUuse+uf3caI/9HBBSn
LSUeOXeg74DQSars2/jQNJW4cL+/wRKTN5bUNz4J1JsiiqCv+xMiClLFqV6t2bAu
1M2vbewjftHwVX74y2UBRyW7UtQdKDofWLQMfpFKi/kFIb3aj56WbXmCNPdUewjk
9E9P6yHxAKuyVOEio30xughO2jXpcrMhdxtxoTe/I/xTJE+wE30XRXmorVpT+qM6
+xMLXbuek7uXKQt/p0cNYEvE48OY98XOzlSLqLpnl+qqAO4PgDuj17RWHr/tUiWU
UAr5fVUOGHzHHWOp3QEZrfPYvg5R6dmV0c2KwkuWN0PHq0FwHJxoGhcKowXFODXt
cpGQ7X5iLoanM5gQjnn5HQ6mLlGVugGokCVaAiaV3n4A6O+qZGvab9sjU1uDsOAW
URaiF3rYuJLV0DPmrqexaH4SBw9DRYN8dv1z4ZUUM/OlSi4aJ4Iiz0cpWsXVPWzQ
lJ53Q0713cm7Ll1xq55fcqhOlo5qyFeVz0Mj3ljOB1bK8wqMolqTpCi+b9G0Tly8
Pe08HKssD9KUVLtv1I7v7gfhaWkT3ttPkOOk4ldW2CWAyRRD81cZhJO87/Ph/XCb
zLhQgQRKGO62K13HKwec2XbS3QdDaOu9+NM+cFgtVCm+o34q4HV0WUSqU3h75Aek
L8tvaLYsAbL9Ijfr37V/I3SLAS+psNCPU3w+i4rKwanLC/ybd26nObpoluAYm9fJ
A7hN7K7joW93fmWNxCWs+jMhem6peyVZDva8TeCmh/xRm99byKQSxIpUNQRXTNbJ
rEKJxhAFSQ47AN+irdbIPdYAc95iu1CY4+lp1sdQ2AJ8s+8PyS2kTyBCC9WSrVrV
hyiDiTI/zD1uDLmgpbRc99GBjq8wMYZ78UsFaV43RjA5shhWMGGHO9QicRcQze+J
gP3vbv4oK++Vc+t66w36YKBWWaOZc7bcLCFpU+YmmZQikYfgpEtLER3tzxaSbsOo
O5BTm/N1gBupwA8ItQkZ7I++3CqqWD4BMZJa/GvuXEzFjq7pwukaE3o3EV9TSW8y
loOcVHY0T2ubMiLa1wZU3aChWNYpI1ZRYlksBvFslatDSFpDdX2yFkxU+YMcr4uh
hRJSBZFKZ6qdUCoYUgLmcyGu9EQNC012oaJOQMC8AdY4bDycw/yy+9lJlccgX9xf
ZCUj2gmGEwm5U3ng58c15OCoo4yZChofgAxq5HPOp/9dHWlwhp2TtMPrGYkzUC3x
Zv2ZgdEsM4gUTrTcNLAUPW5KxoxIstR/+qAILmCjHIWiqbSaI4uE4NWcxL0hkzMJ
sVzKJlabMfAar8ZXt3LxA3OoyZPgRo9GH1xfrMmnaGeR+RySahqhcg3R0Hy58PWs
7UrOtxt2s7m9DjK950vUP9VG5GMzWX6bh2VIzfOYFsYzT8ukuLDE+QmldBVmuldO
HQZ5zqKV23sDcf1K3JTqOnWjENdW/zuhT2U/69QWsC+kQ5FpEBladcAFmTNdnie4
dM5Tdk/593KEKcG3GFkPMQpvjPhnTr18lYnvTyL3cgQ+ir+hyEHD/ft1pvnhEksg
c7bfLXzSVI5AFx0Iwgp1foNPCGBMmDR9nOmLXU0aPHfDXvItw75nDlmY6+9zW+nh
YF+MYJquFapl40Uro31Qyy+gXZHdSB2CyLMzt8j6AnZaEtWIyMLw8w0ebKwL14Vk
/cOLUs6UjuFSTuycEfP9DDnrDfzHlGx2l76zXoNDxyqFu7S/2DRmwNeeslJ0P4qA
+crPfu5J1t/Nz5KTLoF8sZ5rMBn8s1EwwK9p4b/0ByhwW58bkdyXkFlU0dK+tHqx
1Qd4Qeysx0KmUUZbhIvbAWVkoJ2W/vZGCAgkzuo/hU8UzTOJrWk2C4DREznVXYUm
HW2LLE63L/Jie0984odDk2ElrllcvmxR4NxXBjFKzHztAeHnH6ViqVj22innc1q6
QQq09xWqeF/aV7NVXtpFDGlKBp919PevauOSyuCCctZ12aNcGpWMYeJMCQuL2fmo
X4qeughPrMafZJ5BykTF62ntyEpGLYxwX+ct9E2QpAw5mTYo6WdhLwHaMmss9diS
sPh57W7x0hLUmIM2gmucXgJRTcp+VnY6Ch7Z9QDxR6cjLNfVDnENHSKiWhFHpI+k
17To+1DSUt3aMYo/8LCdeGAnSgSxUslYBCbhcfFg9uNN6rZtxwNX5FBAgrpmcSC7
KbqGacldCBK4j3kdBn02rP2b2wlJGy11cJ2smPmk1wrm9t+h9z4SKkzI/d0zQySk
KkVA3bofsJ+TeFMAxU022NVPzpj1b1uyVMVmhGrJBDbXroRclr8F2/v2O6W47MUW
Acqn9kjydHMu4a/KIRVHFnZGGuSrYtAxf9yH7yjNt9/Jt+JDhR4rAAKe3Bmq6377
+3woYvS9twKXQAPr++sAhYirArNI7pQGowPgsejlFKb435sDEpqjqm95i3X3ygu6
narsgoB1JLtPqfH0momNvOOnZfmHOJtgQmzmWbC+orYzjvhT5M6bDoY6G7YJAIQY
dDEtcvAw7msi/9cLUzkuJhFAuwu8SZ1fvyihloMPjMJ3UrKqrIxPvGeHjvOmGYx1
UBhJgv836aP+ZFBGAZXBdJeBEex4QVxDsMbZoeGCQOEcw59xYFESBJEXbiNj5f/a
aOpxb04k9Uxg4AQV3acRC75e8CmSDPomshPG8ZfjHzqqTu6RCFOcDn/FYXXSdby4
8HG6XSUjpLMc5qByyth/UxT4j0hXs7PuZy+c8n1qqqCmSo0vIR+0xJsL1oFMlMwZ
YbyOz/GMdahIHjo8tSEfMorG9BRb4PsocTJOQOUVxx2Qv7jCM3JO4mxRtsJOMH3D
/6U0+CLr27Retdwcl3osB4bMBhH+XL4I5wMK2pKr9MCaJZ5tkrDtWMlBlJ3ak4dq
z4A+SgMUj6ydZOAkrwB2ZlMex357KN6cYmAcEfdkM91rKe0KvCJNJGr1aBHSSLBx
xC9BDpzeFDx8MA9NfJoDLUUrbooCe/RcmszFsV8Nzd7xPvevCLYLx45EdbD3algv
CrjnFWgR6skYR60s4Tqf1hSNVx0a16CQk0xav6erCoZsm9pRnOZHwj1lKqJXNqaH
eftGO/f1r90mGFLRZ/2gsVYHODaerjWL2e3rhElNNx4pnDhXGYqnHXAdm48HCtl+
sliPEJwDt582I3Imsh3/t3g7DdbvlUA6FCkIx18OYbjbR/deAtAwZo8Y9veCrWfF
3UqWwM0YVce3jBiy4H2JYT01WAuYS2XogudVj6IVYjf23QSC5E11dpSjoueQFtoH
uNpT8qPZcx9Hyyh/cp1Vt1LD4Y0uPgpLDptCMLt5POOxH31eLKdZFw8lMLtLrT3V
s5hFhUg9F5Jp2MJD+cJgQCkKIk5ey0pCI5PRZiEcI6Aw+wE0yOjxMMl6qR/8bqgS
NjlW8eQzljsuAyTF7nWXBl5R+PvsWA1Myr/uJdpsuckw0esir6/MIEWvFOWkEBbh
LbVIw7IFf9T4kNxVjxWCKfuKDTPTr/jufJgzhjNu8XYr8Lse9NZSFWNzcYIA55EW
4IMPN9t2yb568Co+gvVPHJPsgitlhAI+soxDJMQm1qHfIrlGcoUaINjZLgjVapRi
+fHHgt5B45jNKKsWDJ1aEc8lULXqE1ZO+VWs0UNz+04znNNOvDPE7nm4Xktmw7pO
g9Aa82upe+6W63eE7Kfpr+721sCztm4T48D3xu3lJ3ExPNnlNUCnMFGQghnpkOsy
bvi07VeEM8cbiEEE1Z3jm/8N0zFieZFPoSO2e+zpZ/lty9v+4kNJOVRTdGtfHcSZ
nmm2mKwfnBkMChHMFasDlBBO7IkxAHM/Mx6AtSy8166nUGBLGacRP6s6s8ecpwnP
CzDjtSd485qrk7qyPPX4IaE0R0NyaAdkVZGFUcm+rmyjFO5P8ZqV2zsr5MJ/10HO
PK5zZrcxf6B/N1FCij3eJtrDx/SxSsy4C86kHxOWAR3HO9V+l+VcjU2nXDbcY0Jq
DpFUDcX1Dpn7bkl6T4G2i2HzP6ki/l62vbcxUPMTdleIEAhYVqphjQciT/SSWRy2
iH3MQfR+FB+0apijCr/hI4BcqK5waYD3h2XHsndUj8JyvY0MHCoP+S+CvanU1BlT
xe0LoiviUqGEDTpv5KR46cJxK95MOCCzw662T1LUYVoiDQzm4icNd3bgIW8wLn5R
AxhIbbIAJr3iRdmLFuLw0vzbZvCE7pRjLgSfclG28X4KYBHDab0q5LzO2Zv0AaCH
yZZzHhQXUG7c0vkaQ2TefmyMNa69L/MP8Ll71pwu1C1i/nosioTxA4XTnqYR/IJI
DU26uW9U9LQsEO7+7ki1/TelnU7MR9tq5VD0000EDiVS1cr8isGwEzh8ClBrhq0W
7roAwMi+LPD6m3aOEuO4gjhXWbKiAbhQyoO4qaGJyZE6SUi7vkbOxx1ImvtPmEIe
`pragma protect end_protected
