`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QwnIY7FKPsQxIVdhVOJiePYlbexfLZY7AiM5V/N5nF0uxSG1W9KXviXfROQrN/pi
6Rs70DSg/xKR+e2LT+5BzgtkPxYlH/gionpxdonmypHjVuAjwC/WHcrm393ZAUAr
q7DYhwkBZsNVFF41725i3w48/GtuWsKY700iRUkBigI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5312)
PnRDv3gJFMWzGxL0Sl0WecKBzLq0xuCKP2ek9HnQM1TlNBRK3rYC9aPvHnvSmOiw
TqpTes1BN74E3XqHzdlZV5CwS1tjz7vDicUlJZOzP2Bt9g+6IIbIPU4gvxJEwQqI
1f6A7CyctHRGLSG7AThAWDTV0Eem4ZYl02QOQkW/ppHCNPhPtrdMtZUNH6VoG7C3
RAfXsn8Z1Dxv915NiipEJs3gwXjyhzCPqVdK7tCQweOk3K7/LEzLB4kWABN9x60Y
Io2tL1PzA4D+gBKgTZ0y9hJgZFCu92+aWX0kDXGjZAaSTvlVOSmF1IMPqnezJ6Dr
6xlfl0FQsgWQShR1seGY0vwBGjpVlFb1N6K8d5p6/473yWnvb85Kv/VpIeiWkls7
87J+7IXky01rS8Y2krmbPq5dxNCEBMhPkE/YaTKWhHE5g4vUjWAce7wDLF/UgIks
+tvFRfL61aVLUcEVmykXI8c1V54OcGsKqVsNQVrG42TY07dHvNfsi6VrEhLUmAu0
RcLxEmRf3day3PsWVSS5BX5zFwYdYE9UEZxy8J8e2e5IrhiY4rB5pRiOjd02EayE
TiVZMmzIMfkcQBqApN7T0q5ESEaaNZH3HOvhUNPQuxBIfZ3PqDh2R7Yh/iGwdWJK
71iyXMYayXAD0ihss1FkW4Vyq0Wb3h23qTSnCoyuhdxdLU2C9sKHdJ3+ezQJo5QU
PxekvgZBklPsTSp+fhpiQJWWNLYYcx0sw/QdZvcuQzTi2l4Ie1pPdCr07Ym9W2TD
ccg3YWa9rtZyXbJSSh3avTbUHkVpnsXXaE+NNRySO80E/HkiJ10QmOJ+rgQl/zxx
3pd8GMs9OtxhNyzjQsUy4IUdOtCVYhZBDPVFlNY5cg1u/iLvYGXicbIzddESy8mw
blOwx+mId96l2ejnvQh0C9xUBDZM/j8pYAo9vXAIBgcQ0hcLrzRZdNf7v61oAvMd
ufL0hvy96pu2Ymb9eThfdZk5M5aW9ONCOzR9iakGpRlixU/DpuXpR6ZquLNcgdF3
zt5jm4dCvf/Vk4Vzr8Hnhv4Zzg8tdANUYvK12JyfXQD+Ulpqsz2aiq+wOKi2XIOw
UYzgL4DSBkOCCwbhfXgQQg3OeFrKdjH+FoXihYchRb+x2l+aqpqSYFfibiqzJVGk
XbqJTReVQU8Lkl2IbnNIHLwMBeCc3mzUxSm/ji2O3dFEcNninJ78w6f2CRLz2Kqg
WR7RfH41sZpnG7/Em8A8il0Htq4/uyoeQf1/yfy6vjrKNg4a/CC7IhboL+gY3rza
Tcu3kdv1ZythpupDyRQe504DpRMkfyKS6/BFDdCuOijUedi9bxKdfITF/qtVMLr6
l/htV4avQVREodfh0vD8jfHiZTGLvCYddj3rX733ujzyMaPlVVqWKzxU+obGAzD8
SMkCyTbdZR1Qb9Ibetq+ZauqOT5Jhi+dreHymAk2PnhvsTdkHVlJQQ2K5qpP+9vp
L8a7Bh+U08Y56TCd2E4jW8hEsF8MiXPIVngKZg1daIha7sFdc73c8eywFBTbJPBg
OBEIA2urv3Iy/v3ZsYMChQrW1ha98ThspnTObtQPEJdfJaCNdF05vAMNrU8iOf6k
efjTucPalrVsoFaBFNV0DW/iHUQT1S2dCqDdkXKdaysXjXPGydF+VTXFd2/7BPLF
BZbuZYxDm9xXh+6DHxHL6GNJU1VQL348WKJ0XRPHjTE22F2THEbdZ/TDZbuGO1dM
+9SIh3Uw+cY1OIUeBJZsmkSIRz6HgF/Kw0cOXpnlqDPiPhvkkaY0m0ShfMFSMh6a
1w/jppeOlue+MvEIbrysu/pePHymGdGuTOwR2m48oC5vuStqlfDXlO9FKXGIPZzs
F2uxCCElNFnk3B28BQrf7rM4l+d2vZDSOsPaJcqjWvdzqLwrTGYjINa7DY+unFM1
oJqWFuyMcLC7KbG/0ldc4juuBP8uoYZA2iItSqQQefu2gVrrbJzqsuW4e3SOBthj
WGzA2KlU+7OovYMwyMzP953aDdrJr2mfoBkuiAPcSdfkEq5qWfRTkr3jkttEJCJZ
1aO3IDlts3/lKLVJf0f2Qup+x1WaVd8QPa8VtOMqosXhThI+VCfVOLsS6gU86ZIx
iY9nR7fWM+JW1pBsZOJ/4fr68Dh5RfOeolNepbSzM4TeHPY/NSG427dEr+1SqJa2
ICF793L8KzgKjBnlYGhn/ZBPYEeY5ys0bWSkBYIQeW9RbYu/4UzlayOIGyIFqmTd
EZlzMZUH74iQAPGp3nclLp9K1SR9NFAeVaLwi9cSPoo/+yj/z8i1YptWJajUVd5O
yC/2KSVEHpbu65vo1cPjtft3wXZcvc/Wx/8l3pGrdte2psBRNEtDDya1RtNrKHqP
34C35uufVE+O5XIQRjH/oftch/YM+78QH3sk5tYXiywb/wVU4CKNycFM2fMeiD7I
PKyWvj02ux8VfC9dKawgfHSfKfVu0s9oIlPgdLuxQAyCJFyqrlVLIUki4br9H41z
Ry43LCnqpg0BPV8Jydp83b2gLyrqvQwTHVFnGRNDu6EnPtFp0PmfvQ7JaesAP+3J
W+uqeqjweTktU1DuZRYiMaqtzZZjHMPWcaUD5vC1Brf+Pk4heDDiePYagKzM2OBl
kTlCmlLTLDIQQHGj32j6+I19/T7YAnav4h8PDba5Os6TLiAFN1ybaP1kt0ZGl5OU
1Tr4Xw4hjTJNJpSe1GkoAjEbmbrDSh8Rq5QsYwRUYoq1+oXplEe3FOLDPomowI7T
7QQHD5TyVU8cgOcvub8W5kJmA1XVOyE1+k8+oqkSmJBDNJ22ddfCy4fJdVu8d7cY
ChvMU+iyEUhEreyfEp31mZplRFNjlcEimF8HmZfIM+8dO7bbRzp55HGgF+XfWIJU
i99TaBUMViSwZTPV4ZceGKG6e2m3GV0+CpAtn3tzxpXYOiVRyphZ2hSTMPRuvC7/
+Crvr11XVgNKE97HH9TSdRXpVBqUYsq0tgpream/ZBR5ddAmnvecNsT2xIExoXIM
5R53ur/rwWPKFzVLR+i0sbC+hYKOJWf2t3hc7Isj5G6pi3WTeQwBL2V977POiSfb
5ZT1qEnwbxmEXv8MOe5kf4WOOcO5i7rr083X1t+VKwtYIQRfaKDiCqMbwF380Y2B
WL1lMeavrmsTmuI3gUOqTfcVpwAer8kg+SxFGEhrC2Br1RSMShGvTnAFQwnpkk5N
uZHqpvYkhlX0QrkhWmrPmTvr3HWLXCMc1j5Jv3Zac0szbPBjzde0rJg4gN40JdCH
8FpZFkorgkUznVtVUYMMcg+BYyklJ4ZA7eHFWJy+AbP4xfMvBmxZffB9ZlL5QM6p
kwWrpBH4NE2vcgagLye9OwYVXf/umlhM8D6B0vTTfSg69l+gywoPdJE4ieF7oBOO
ZH+ccl3BL45TU30x2Nf++rJHYXjefbEtzxWNuay3W7Yzf0lFayvzQVREg8y7OgF+
7KAoOsvQQWROpt6F0yTBvv66YLDMI8k46bEZByGiPuLdjEu2Aw7GglLMCp6MZ4K0
eAxUd5NXzWeQZJsv5DqiqI76zVddsEDDpU2weQnSaVqHMsHw5X+DX8HwR9AuN73v
BqT2i9gAmHxw40SeSmyvGrp4jN1sH/0wLxPLBL61YzUuinB3mm6duP7NW+LMxM7I
I/Ob4yughWlKPgygmg6PXcHnBtOpiOsG6ChWGQT1Y3FsRNnf5IQO8jR5JuisaOEg
PeSvsH3vVoTWESG8GpHD32/n0jVWWcM2Fy8dcFS8sN4Uy9pi/EYvZTYujFvo1O8y
30JspbrhyRfmf9nqBfsrkiWwQ83BvdUcmJu40VU4eE/JnIBsQw8pVt0f7MkMGJz9
Q4kP+20MzY+YL5+BtSFZaPluKVfJFhPXkVP4hcXkmpB3eo+hxAbUdG0eNAdLkUSv
wJJBsOwrk7WMrqHZfj7NJEAB4G/DLrvctQb2Mwu45CQaGOIU64X5FvJE/ACYBSii
JMIUKE4D4v693XcZP6Djm6aHn6ZC9KZljNZHe/CHord54h1z8vyCyoD+gBkpee9V
h6tkGvK5tOj/V8vQe3W5jD0TcFwbaiC1RmeKlNAebSiGIMAaNY/+QWqljGSujmaq
jcYOkMQMU/uzvspTaUldbofdQvX2X/ofZCJGvs1pKhQB/wrQQGMQWEhdt6LdIHjy
VDwBCn6UsHdezN+eSe01j3aCg/gU8epY/Z8R/5KrBhM24dm15HU6XIuiOk6UH7YR
0c69fNOOANgAtn6keB+g0Hf2oaK6BCjJMK2NnMQVaIYUzGoWeZ2tBnsY6rNMfjvs
oGUS410tjW24qbdm/Yv9MY+ccNYhZb84Se+yV8r/gLgA4R/fkiLwM0QjR+HOz8yK
w/87HkAuogqHkm5pcFV2xllb0LZMCoLrOTuCajIeK2KP6p1XOlrSW7g2XrGHsfN6
yjrA/i/kygpMNwOB6p4Dw0qNWhc+lUbOaLVapSWMSdzOHwAMD4oSojj9vvOdHNBe
qco+YYQIFCi+o3DbyTxVtEF01tQg0zKka0cBfRnw3kH2QBtmONEEX3GuhFEyvQ1L
YQQRuaTcd0Z1XBGgRWNZyJp8sBi6tzEsq92+RVi8mAnbrZJLGINHi/YJjZjTozxD
fjUsfhk0ncufCW6HYXSQ510+1qh4IpFWqHc/piswWuFT7Sqk+ifbi8NFDK2sfnuf
X8USA7ReJBElxOpggGY7EoywpNs3XpPqjnzVIdyZgZzPkl6SPZwIHYml/TbI9AGY
PFLMtUYU3Qf74xv9U9FI/7vL3qKcr4p9fN2LjrMoI2Z6JJpLdWt1OaNIy7s6B5KN
+6LVf4GbTxoma48JUXtK7fIO+MfhwMxp/wqgLYf6TFahBdrOBIY49l7Ya8FxRLfg
FtjXJ8m9BtX5pzQ5f+E+HBW/3Y0rZvMCuru6nQ8m3DX5Nuiu4ifenBjtiuZrKTM0
Y0wDc4KUWwwuaXnay1/buG7G3XtTMOexHFUzEquqLQGMkwPIwMg9HD+5xY+TLC2k
J+RFKLmgJ+ZHcpviO4GtPA8UBzcj6rT3pYHHzpKk7hm/XnW55x+Pa8QXr+DLYh19
UX+XItPVNq0YpPz1iB9otcymTJFtPina89Pz9RgZWi3iD/4nG6uHUdqmaEEEIQwX
ey4g915+yAThI4MPYb5Oz84CQuehE8Wc3eEp8X1+3iegnURWlGOyXHZC7Ain6Vpa
Qdi4RmDPOsIlCgtER5Zr6kwla8qa4d8C1oMrZZJ1Bi2oXB7axrcx5uVBHd9E47r5
Y0aCf2toPlXpkoJlJWCthtnb6AXs0TNWicEYZOFy4z5zmmlI2lY9vwOzz1BBeJWF
EplSmg7rdvtIHUUKwLkoL+zcLPCCU3j4Uz4XMEeJv4WHKKxSX8a/I5j6m9s+mqGF
jklY/PX75vOBCmnE8l4ivBuRuB1bHSQ9D7zJY8JJPkSJud+Q8vQRw/3Eh9x/UP9u
QgoKJpT0582q04KGpOMxMJNmMLDYKeoGQpDN0+1cqS5hAI1+O49mIBgmEh7B/KPJ
W/J8dJglTCUMdV9uKNYMJ6y1ML5BwPzmR5N+jql1XQO3jvUU/2/zelwt+IVjXw/Y
A16+3w/C/nU/hcelNgUua099yDXdsoATGPlCLj4fmgoybOZjAj788Ah+GyYnCLKJ
mt7ErEpZU0eNPHAVWPoAmRUu0gnaP9Annvabw4TeGM6AvT1oh+v+zJXZWe7sowRo
pEIEKS/SporG0DjzCIg7p0ZLJXiHRmtXasO089IWeAEu/SsbtSs/HX1YPySOMOhR
Ai5kjdiCjeklpjIrOl42MWOgcx/desdWo12viIVA0q4nsySFjTb1NDL1rOMP2G7d
+paIYieRAG+ffWr/jPCTYtBLl6gcK28dI+5c+9U9pz1/3R6kkkP2WrzLRD5iiu63
WzwZTp+RzvcrVjmoHBggZ/oHr2mmE0FKAPeQo/KCD5fV/jv4WbU2KL0g64wgFZ7T
2Wy4t99WsbOribEJGMAmZJb98B7UP5ZTc3NsvLw0kNE03QMZQ6UGiWO4bB6NDh13
UnkJkB7ZP3WQUoFq4dOsuGiTCA0hWmXsFXtxIXz4Cm4NkACYcXD1MH2spjGOqO5a
IFujFG2VjPk/iR2WJsx6E6fSyBlIMnHkQ6vRVa9gbkZoD+0W7vBCuWCAu9OiHUSa
4+XlT7aegOcd9WkGxe2AEsd7xgZR4VwVCJC5JB0tukc2zmHWRFsmAUWt9+0rSfU4
M2WIhtKwsqOkgwRZ5tk5X8IgApK6fCIWoJ0QfvjXMWqUAgnUrDMEkS4xFBuxuLhz
BwgzBfO0VchpzIC14F+iMWdrbzYJ7JA5+/b+eKq/TK/rd6Pq3viWfYgndjaNKHfZ
iMCUDH9WfKkvwwHg2T0f1hBzkisEZdDHmgRxzSpDUxFkKOeV7HfEIEKTmGzWyHw4
tRdY1nqQB2eQPJ/+swdpD7ZCCqAAJjPiqU0lekEr0JUeZ91/qLy4dKFh3jejYtnH
OluqQMFpA+VsKGMh4iLmHSE6lO5dOybcXg9rRsoVV7BfuXWSfwITRGfainX8P2ZB
7xTKiWYQAbSQuskTkUhu1NqMBDGBmDF8A06h59DCrjGSUA1ofm4EC9ht45fFGDA3
Fswkf+txBr+hlco9rFMrjqcVc84iPPmCNOVj951ysQ6Ux+KWk4LrLNNyBavJzRD2
3w1AKPzjPNHEcG1I2Iq1I/0NCF2xQ4DFIISVxukhrTyU8saRSJHaodJiK4XGxu7B
EDKwi3JUE4SV9lc1PZ5TM+mZ0mAWJvu5VGtXenyR9pQbmHxenW7AKUsuBFq90s2W
lesx1MjirceSNZc4XXwyIlS+lud7TH0ZkeU1NhPeUiRumr21RlWC3G/10q2G0gzy
Kj0+W0aGsRrWctoMv+qUg4B8uJKHJcmXNOA33fF03o48mEYBFkltypKemTLcXdrE
6PPYwK7Nwk9w2omm8waIdPltcW+kZFYpvKzmY59CF+Vm4z/qp1hrFaAiO7KaKP8P
A/FiF1KXivfkHFwbtL9gmVWXM015AWZ+d5CXXbv0Em3mAys6c9CUuZZsuGT4rIM2
rIFhj/Oi1gvxUaTb5Zr9Tm/IiSzan7uRvTmy2B9tFa0=
`pragma protect end_protected
