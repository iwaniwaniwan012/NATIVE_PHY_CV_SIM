`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CJYAHiXJ94RBm79G5UB7uXwDwV8mvHmtADqY8h3h8+wfw00ibhRxkE65gAZ0QP+n
i6zaVy3mPcs/rPPRwYM/Gz+rFPr876UJ1XFRTyqvP4lppEV3AzwD1EXGUmulIcSo
2nVVvM+r7TBrq9Q6pkJL4Yc8yB8nCybb24RGbj/nsyk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5456)
bmuYkoQL6Uln0/vAjBmtGMxv1i4COHvRrHNh/68mEjeO2pDeL8eoys11odw3b+yV
WWMakmZZMG8ASvVOgHNmL2m31Mp3txSv6obU1kHJe9TuFtapcdlDwhX78AccGu37
2ElIhsFbuIEN+ccTkHd+kVm7rgnzsxZomqpyVUCoKg6eMorrdk/8+fkjrInchBXI
77UvchcY677hZ4la7U57a2gtNPpwYBLMs+y22Z3o0oQTaWfUJS9yPOfo/6Lpo3fo
biS9hNNOwhpyl/BYgG5H0I+kcYCfxoYjnowsNxDvwIWojO3HPjg1dYmloUYKv8tY
++EYbNxyJaPYjIgUSxvDCOTTBaci1WXhHLz471zLuYQtKR/Vn8/DawO8Aq3GvX3p
ReMPxfj/ZVP15L58queFYuTf8Y3OE2ggUkp0kLHsIURJWZxkKqG94TPOfwBgDCRv
+prZrwyIuY/C1LwLGJPgj2zScpsthqa3KckOoLloze8Qe9A0nTdkRAVb4MGV4SJz
3ohpW/Xusnha8kFBfhP/x88TR4sFySzzUn/FKLWz2+uRF7/l4X0AbG724f5AQ8pt
Ed3BZ3dSzh/vnaMbwyoaMyxLs6CcMLTNputBT6an70FqKn263jRS/7cOmVgIZH2C
QH7PFxjGt3NioSV2r/kNAN/Nm7LtfoY3onxopsDcHQ+a6S1VgGwQvvOsHNvIUsvH
pcHR/0ao5i4IpnvNnzBf4VS/R5hz2fitlP1v+bro3ZI11EFwJbEohwoXj44Q5RyQ
VfrCIfmvEHhK8hgMesSVjG6HlmBWFlMDkPS6XufkbsfAwGOEFB7Juguiht1EeevM
TsD7llD4jfQ5nF9AWJzXHDA14JsCtDgl1szk0EmFoDt7oiL+hmUL39aJkEq15o4G
K1+l+xBMVqoPoIdWL42ZU7YS9G6FG6GIx/UKNt6Sb5zDFu7u+SDd3DaZdfxWgw/6
b6ggvxX9PK/f1dyMH7UibbmAcfTyPTLk31NDe1+E0wfaPUdl0+FJ4JgjEzySuvF3
6zZ9Uw643HJYGGZUQDM/tElY9ltyymFRjQMCXD3YphBK5AOc/wp3T6g0oCZiQY9t
mohDzvUm5DUt/Km0ABQa+5envhKRErwvNxhTt6yMwQvFkR9L1pIFU+wkQqOl+DhB
tXk8BeiuKkaGDeblrvO9YYRowzRFbqY+1E58VAnJrZl5ZD8y8BLHZ3HFcUkPMzdV
m0JZxU5cjXEbryPUohlfwxV6MQo8skywksagl+RN05ZfyJXhdA94QNTVJexDVSDt
YfcYBF3nqZK8Nn9CHEWw4sA+he4I+OOVC3Sf2RSH+1B5mj3aPeIEH5U1pyBp+FlP
DQk8IpNiv+Zoespou1wk8ufMXh+V3i1Wj26wTuHV1Poo2FgVXNRYYCAEIWkQJTzH
XQ6T1UJrdSBsxU3iHS3j4awjeYDhBXdeImc1zfKqV71COvexMj5FfxMawpl3iVTD
v7yD/5Y5JLuhW0jOmd9QLUmAjkvqpDukJ0YSF9LTUC5+Kayman88f0a3MlFK7dc7
lia2JmPw6wbdtK4+753D7FvzcSgOQ5Vnz0GcWlLV7QLi+Bgc8Qd31O/ctaGSOhnM
EyfFMZTWnolsSwftlOU5+hnYgs5yy4WOw+U/U8Kvwae8ZFrfxmWu3Y0/09ECr0Fk
ljzy4nI7d93niWxJDKKkXDo+9ce5V7wgzbipHTAtKHZJFcuc+xvTvvIsef553QbL
Y/UlQEjl+NvMsNq3wqo3NO5J5HUmrz2aotGLoel8t4PRNa7EVj7fdFYJM7Qj7JAx
U/sDzDuyWq7hf+l5R3NNptvJe4zzxgXXE56LMELW4UseqBUa1/6leW0ZSglflwrB
33otvm8LvAraid2VyJZvyUGUxRlglshwEL2+AcQYJSWGsv89h08e31/dFyoFc+S+
Z6xzNonrrK6r0u5jxee/g25V7HeSMO5qFtVC4vuSn6JZh7LPz8y7O02SmXwepv6w
+r85y6WKzz/li4HfaOFPHIYzQpyco2EHhPm2WM+PuwBICSqjz8U+Boh30o0MATZ+
yvaFJuI/P5Sk0H4eejsEO7lq9ebgm5N8c5XbQhOFs5f8NX1uf/Ps56lU3q6SNoan
zAiyk/RehTtxhVQ0r/l1uky+GtIhwLv2hmPC/3Bprc4sLKmRhLBtmeCR3+Hwu0is
moGFyFD91bim37VVR+RZmRazIwAAK7+IPN55RB/48/wg8VZWBrS4T6k+Jur9Ypw5
iGCa57P9iebhm6f0Osqb5fFi23vQKfnODPovqX3ItU1TLHSGNB3IjgV+gIzYDa5D
4NC7g0cRCTfSkfsiKPPVmnIV01aCh5DuxEZXjFy3MVC/kogDimdmUwuYv0NVS7io
Fn6YH0UXHfIt/dRj1d5L1tYHMaGKhmCdLDlbUQe9DF4h0IcWt2hlgNmPlLvW+VU/
PPZfvKe8042LUAyhhFC6kun9Wp2U0HjubaM85vOgAASz3D3svkbucd2Km9yr94ul
E+V1X8gfWZLPeulBM+tCdZBA7PT32XkuaK+nmJyzHzBCGSxunKWg8ztrePr6fEtw
h2ZDbbpwoVwkQmWUuysPkzr5I9ikA7t8Pb6Z0yAad2sOHoyiI9UobchfbyhiOcLU
KLgSwBbVw6oPaobh413rMlDrFB0kSJmdmgj310go/dXHk0nGQTX9kdn5egFIa5uK
cTRkrAykZWSriJufhy4+Yp5BwpmdH0oB6uM1WhPxhW0khMJbW/j28bXBhdrsWzkh
TYmidXlWsSz4f4vu4YgZMoyD8ZgR0dH3OjcftTdKLvgIR5OKefVZG3jPXAVplsYS
J5d9+if6skLc1EmxCpfUzQmnFL++jqCa/ED6GEp7MEENwgF8mlVht2JglsAh0pHY
Lyyjn5GqPe0b9Xp/rQN8TwiMFxGDek/ArX5Vu0yAuf8QuRp9Tdhir/TWEHOLepmn
BEHj3bv92OfazB68wouGcA2/D2ls+OCbfQGUHtMMbbAp8La2NzsvSdtuJIVUiLR5
vAf5ibKARcevg5kUaqWp8PQkBb/XxwkH3LyZTqJgbZ+19rCDtzrNbSOC9ns8GiPm
5g0V54z5xPpG17HhLOSx2k5Z6VoTTIcNqL2vK1CqUZxzpPCO+kQpggec3rvE9jBI
W/X+E9sENodjZtzYw6UbMxQRyaYKEhelsM7KRKUzAYC6mHN2UwDaodJiCE1HHGrq
oPy9Xv/F9T2nuuYoBvIIE5LuLAoMgbe96NhVUhe2fqaLawjsZwTxMEvGbUAT3RxG
P1H1c8DodFxbutgN5XmbMwwdzrMe512v+SPtwxYOUIaiYuP9xmr9LC2CjYC29ypK
xUAYl+Mw+8tsMN5GEgyPX16VIAi45pOAu9LqmRcmVQTdNcZL8zZWkcI81h3D4oLx
/Ht0EuYyPmFvKcb68z8AiFXA035V+dIEKQCZHfJGryz2ZUM1tLkCgsYJELPGyb6B
+ZCcA5pdI5Wx1gZtGL4nMxTJLCWSFKQsn6XlzV8PcUeuQ/o9O7lNof8id2LyHpoR
CSj7kYhIUO4Vl1kS6Wcp5pF+orGMZwYUY0KtDwlCVdozqX5K4xf0H7K0qM/artMF
zuxnglqmcpwY8H5SE5CgOT8pJjRi9AEyJpEpy2kkfyBv4uvZRZkxeSzfWjiulYxZ
pBJB3jCoWYNF5VGfHuKO5y+QTpKwj2cuSipgzSE5WhsI+/04btUyuLhTyXyyjyrr
adeOt30w3pijIvA0DCAolYMvvSgJyIZSzrmFHwO3oNYqENTEO5uVjEWUq5BrPNh4
QBtdK9XwIVtcG84SzYrJvexLx08yOusLnnMwClAClT6SusNMh7xnfvsjxcgF3Hjr
sZb/bnF2fNrfcx7s7ibTPXwO8fz7lN2VMCfC11EdPKWB+2e3E12gGbFarOdOF347
HnURuDYxnBEqco4kFrJ3MFYAvPcwzSwAnZHNhJLSGDd+oLyLg77iKx3eJXebSnbt
QUQWw/BWfgAxoQZj75NltwJXSp2jYHG1Z+z2t9Vj1FkTssjsBXDehVv1Mvu4EnqC
VTwoPzQMz6uoS/fbX3j1EuSzjTqFAw/nfw6F1lVL7JvXAeAB6jumOMApyp4Kqa42
3jdZ706lwiAavWs+e7w4Ez0oi9RiZg6kEqVAIFd4WUu20sPa8VWBJ2yN+35PSJxP
uoizrws/o5biPRZziG5Y6FW46qQ2gOuFzVUz+boB4T8NtFoym+UYQfmksUgdHM4l
KRGMu/s5zSP2aRYmQVzl5Md2c/APvbLhqFlAn+eVXf6PUy0oOsEGMlUMvfWB7jRb
hcE6IbzvoCr7jpepRyCFO7q/8iek4eMBV7nCFiRpa4Ezzrwydw12W1t5k1JYhvNR
Fp8F/wsxYPN1j+DE7RPWyiLj5KAA1NmWKw5y+LOKjIu8v5s8CuyWTUwrvKLu4zDx
+Q394WTUHyKoRvPnxxPTkFeX0peZFVLedjv7iaR1Yl5O5iDaJ/3SZtjFXNk9M2aL
yzT7fl8B0qumpdRP48+fkz8kR47e6MD4SVaNs7xh2KvE9UQIqEnfSEHPt5BChn/w
kvQHIKA4UF7qC2TY4wAIBUaFO+L3ik8ohDJzFA9dJogVRtywO/cjxspPmL/2uaqE
W/7i0bALVAMYXDHij23uRg/69o6m3SAXR9QghPglDln2s9uwPsQxK7n687SnlQWa
2EBi6mW8sI4HtkLnwGymS2EWfTycJdu0ebc5cU6gODVixaaXUI2vjqj2AxEi0X6l
I1sK+RGskiELPcY27e5SroNTY8oIxB/aWfVMsE5HjiG64LKOdLtYjFk0Bvz0MEMb
HfJj8Z4GQadvdJyHfpOM1jRSXeZK+/exQ7DDbB5KwCEI08t1tSWpuHvVcINQg5WV
GldRkTbq1XUMacZulyGNjHQGCDk/dIpc3NeQQvTmv79bXTCpTrNQ2Dra5QGPXcx4
XVA0zJni/o3cL+CGdj7crA5bWV409ASVtfQHukt4t62MW18A0XO5x3r8FGWmNdCQ
M57y0KuLsqne4n15wnR7IYSqEHeFscidNAtit8iNyZNtkBy3rT49N6asyhIiq3aA
GWv0yYEu7j3l8O92EKr/jSt2miJ/WyoAbBZlsJFxo9QXf4qkC4AeHtPKb7SNXUh7
AQ8bH02Jx7TDF7SMjodVnZJSoiM4DAkCCQHVh1fyVWKOa4792eJUQFSmhqkjVxhK
0QUYpS0Fw/eGVWWGlnA9jHP4x6aD84CtCa9RaeuLDcHnrGg5oBMir3e5Kvp+ZZo5
aMEbOYvzo8BHIN6Pj4jaST3MPnlJjgIjDW9kbfN2L/rWv2YLJN1Fgc1O697LyURA
TuApdUr2iu3AboR8JW+eU/2HYPXVKNwxj36Z/g9f820N8oyN4eIc0WwwicZ01nVe
hMw05VbJ4bEWNTHBiebmt4MpJ/EWVuX5mwMD+L11wqXVdxw3/rhw3RJLGabG0vf0
1xuNZq2yTjWsZxJhlesdVrqo37K9EVo79Fq+XH73SdKO7hgrTe/HUFVMTQxV8wB4
x3iTAj6HWaWjK+PRFtd9Z6Jb3fpYrbz951LVOIXnudddKJOEoxCaR1tmA2frBr1P
EYtuWfEwcmDuSjvLSria/tdBM86Ds9Fe86MZF7XH5GLcXx/s2Z9MqchQC50O4pBO
pgYqnlLO+SW+rnqeBcDDOY7P3bxxf3PHxIBE4OXhDDyT+L5ZPNu6ncnYWv0SscPT
5PsUaN9ppQFlITqtqN8lBA7wEbGPD0BSTnu4MWe4vUgZMGCEmN1u5rLN0LvW1coW
UrIAxMTJ7RhC9F9Px6upWYZoCfEbR1bwkOJO2AUIhym6dTeIihbuFYwe9BYI6lF9
MWA2qD5c/6uQLipQRpP5XWfTXcT+vCfgtyLKK97HMgrb9xNY9oireB2gvR5YaAAn
csKZmd99ZoggNWFagvjIIYYL6okVP/+WbZXBpqENKwctdZ27Seit8P36zkaiuG4F
l7vND8x4ucVF20wzTKqqF2yJuW3Efd1Km8NP8TFi56RaNKgeObNhTG8FYvLIuupW
z67VD9r1GIj/6HU49189yxGydj+W6N6/SWf09CiDoupwS9jwgLjqaNoI3Nh2l2i0
SpNH2EHdjqUFj/z3OGfKcTp02aG5s/sFJ85r/huF0KQ1DCeqQgBD0y1D3w2Uc7YW
mgTZ1OnUu9VAKuf7bJ3cp0Gu+kV6rH0k7n9Z303xJRXkOkR8o4An9WBDoyZFzGTD
f4ov2LRXYZ8K8yBKyicMCwW+9rOXHQ9TOQjRtl5HbGEQ6/T+wSANsCI96O1yEwQk
CbHnF3Pj10Q5xVB/Zk78Meb+ATD6ozW3tsQVXPoub6UhziXR+PYSKXN19iYxheu6
/RB82jwKhwZ3ueVixjONjgwgl8tRy5idP6kV1qS9M2gQh0J7gobPhJyciJr+LhbH
YjBLgdTF0I9FLMPpitNh3HWndVwsk0XEZwRXQfYwxQu1O0W5rt1rgHP+979xAf4P
Hj2EmZ4bu5wNNc590gU7zv1wmO80XgIYA91HfcUswfHjJmP1f1bw9we0WtmGD4Er
ZC5+59Q2JsTCVbKmfxgbpD73s9t4OaVm+nvA1vAb+Kpc1Cn/an3Citwe2MdL2Fo7
YxUBtX7O/sh2DFOOYKJhwRXSC+qjlAGr1QsvzGF1XxU4BkFaGjqeWntDUSQI0l5s
FRYIZS1FnjppLgliJt88uIwOqSG8q3wg4j7DPCzZehiw9kvJETIcMNMFqIjaq3i8
N7pzP5RpGw6zxi0YeX/6/Zs5erlHBgPsxM2fr3vvAFRcaFkRQq/3p02YM5JQusM8
6+oYyj0Ji07aN2fcGkZsfPes8K9Giieqe9sY5ncPAvgt2zRfqJQz1LHMPs6WlQlL
fVJkTNYaaLn+0hOEoVzxCLcav1y/zJA4nI1lO+4UsnYONtu7qqzgidXZBPk+uxTB
ix0AkLyZDSD6Ij9XkjK7RKWcN443V3eQcJY775HFto3kQYo0VCuPd5ytThzGI0TM
wUDG1d/Vo7QHzXbtU1y/Tr+tSmFoTnOTPfm25r+qrgx/V9QX3Q4nq1RacF9xMy4Z
4NvA6ME2W/n3RyDbgS+s4K3jGJtrqSYY1AeWXwgvq6ndWsVpgh877N+UAjoElrUM
ECAXgmHDYlokvzy8snn8Ie6DDbE+cNGbsdQDObLoXJEWqsU+EUcLa7zHdKJ9EKTW
XlQR1IQFf9GQRCWwr0t6LaGvHgJ4JuDOEAeKcJz8Cmrpp22UElfHZJX0rpCQGfa2
rK6XAo6eyBYwPcbmAe+PfhyeVAXg5dyQaab56IyS7IE=
`pragma protect end_protected
