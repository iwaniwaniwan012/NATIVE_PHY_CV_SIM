`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
l/+8UY3SSrB6wmW87zad+7XOgy7augVY/GZtBVpYG7OMQsoidzG2GRoocf+J8NG4
QiFpc3gmXulBkNjR/PUScVDh9B4RZDHCwtp0JRY3o8ZhmCL1bnXbSvLtFMq3TNLA
FduS2ITpjd/rbtu9mrNiNrmvbJoK1+WwbxgFh1OmskQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12000)
C7p0/gsVICwW4zrCNe/QiqOYcZkWNTA6dgepBO+EZ2+Sbbu++Ph7ramKPmTUN7gJ
xDWEaWl2qg7tuqs4enmDasyXRkec/Ku6cOK+GfAKXTIJLAztIb8IuRLk1eQ7vWOY
l8Wdxj6qDB/ts8byBIaSV5DLaD9WywtyNuJaqdbND8tsWsXr4zLSgGGZF7h5Qt4J
YNWvuiqixci4+YW/9hil09xy+M9Xch6anGd80udus90hqZ3WunuHdZj0fZ9ZcPzA
oH/u9lBkv9lZWDSp5TmmqmBuR736anNpKB1Ge1djTHC9vLEYupiuQaMK71UOzzLH
UyPr/ze46RRkN8M21gG9iDbIl08jRG9hZY0DpgVUEeqaQ0Q6+gdAhs9PY5lxSncs
fBGC08qO3NVAWmflciRjMA261XWoA85pK2xX0Jsj86XM68xN0jkoNzmXiRdPDFkd
HIquNUZqtQJ33uur5CPXgQuSytp/9xNFdF/HXuXTddWt3dTqcFnjXFdx4+2sL9Nq
RlHlV80jn+bs5WW8V+v5Z4yqBap+qsjCl8hFzqgtPkZwJoq4dP/1hVx8IS7g+D0p
VIVmBT3D+YXJJleV4N5KilWSSpfDSw1JQPL+yjX+mm0h0vBQZcfsx8ttp14lT8Aj
IOBz5FcwtQjRtGYPu6mlP3gLNXxun6PJ+MQYAtd0jWolDKXJeyd48DoRwfkMYFE0
lEqKzRBZTrQIqHOSvCB8bu5OwI+AvKZafn7N3iZ6rhqpcKtFugjJ06ahQBNrD5pB
1o6L02t7TucVPao6UCflifBcFf/s4mSShYbwXjjmu263CM20zVmBI2kmd13odT8a
w7MHAzjmcHqSLCcYHi7DxC2UPsUBl0qDXG1OwUxj88ScVKMpqAIbIpt2F/MI6/CE
jnPvRv90H8xkyDQcCCl6zk7oIKK3b5ocUc/kGMgSsWOz3b/4zMVaJDwRYGVkHQdQ
l9XfZrUrFTcFN4TmRdI0UCzkVXBdepr9u3joWYMLZkUiwZ8X48iLOymHnNq/vG8+
bsNCYlsWN1Mv1LgvOuajj+oOopyN0iCfndUCRXJPHG+Vtd2Sl9kw5+ICJ/kGjcdU
aO0bLSo6Vuv+JYgivAFFfcrhYj9WRUdPJAhOFyAFaroZAijl6oMhEIg1S00+vo7Z
XVZTcgG3LneuxUrSJeYigB6uGybCTgaw/56gosdWnQvn0eZOyJscLu6D08WgZh5q
d1QrQVgYfVgMpx98WHrHWm1E1VitwfXKLO1eMetcWpFm2t7wCx7zd8q12wWl7afP
jTxCVUDl4RgfTkVJM6yrnHUnhHQ+ITu5utpjQ0XXWYoQfJiWLMqLBtXNKScvCj3/
fpV5SFL91IGHpgdRh1j1HoyK1IpYhLBBCIJnzUB3Ek+atfl+yN5ICho423JV0FRS
kH8ThbcK6iDaX3uPTT2XhZVHE+j0DMqQMCMCk6/K1dL/oH2IUrSVdr1aTT5UyGIT
Qi3px3njpAlcCK0MwiSuFD3ckBNaSAQygEqzI5sn/i2Xe91a0wgWaRMvUY/sGyRa
BJHF5FRfqcOBnVXfaYdlOK43DoTgcsaO4OVJyR0Fkg/QBw1d89+ioHXZntR3azsx
KUgQAAr1PD8cZOieqIIc7M71UxGtWnLfbyB0vwq80clZ4goiq3giKxDFJ/aJDjg4
VxrNplgHFu86gXhRBwvMV0RD1SfgjNMiAJSW/I3ormc2cGmX8bWzZld0CUXEAtJ2
Esugq1U23Cyf5AceXuvRcpKw0+s9Noa3W6MdT+EorP54+uszK/gQzOIbeoDmNb8b
HWXjExEh9TpyWCWByKjnOxPtBS7MN52GhoEb2hghvGiPr7Xz2Bwql9qHCDT6goLa
7aaqJVP5ecDWD7JyP3Hmr0Q3Tbk/AnvhwzxjqN9C+aGniE4WMsKgASwlHrVPWpAu
w8AdwMONJyVXVt2l/aP0qDw96WJHRqOruJm0+ORaDC7pdMqY8B1rSgtC5V/h0Vab
mgi7zgdv0eu/cSz9Lvg53qY8MUmMl13UAxl5Edn/zZU5rE9ozHO37+5n3peWwB3m
9Fkdv8Vhd07RAmD2OJ5or65iKGmgEzznfKOO2STS7JCI9p9uMH0i+Ct4QLB0gJci
mDBK05AM1D2qC5S58lOIhETOLGPnNaevbe57kJZty80fgHzIEnkKKspc9FS2Qxm2
Ey1Ty35YQbZoc4yFYsIky4POrXXBAiDBW0Ml/CHnhJu48XwNgsEP8j2EGmbX/iZW
PFxrX+oiRvdzr3Wpk0MEhZUa5blIpQLX69eO4S0LxdcOTMx8Fv54ugbOxGq1+Xg0
LAfMlFG172zovI4KJPmMgCdHNfg3uaFJyT3LQWL8B9v/CENXZv0i0355+vmum4sB
GyS+PGgq3Thsf1Z9eiy1+4iCXC00X4HJglqTNg7tXgE2XDnJF4VhxAGxahhrR2IV
3J0QzUg56Xwn83FhbaUTVJi1FYEdxqZTpU6Hz04Vs77QXhosIKiR8eCzLZyHPdBn
DDnyE2+m+uv5gLQqPJz8Pnj5iXyiiKC1+6vWEdchxtiWRzqIcuRwruivUT/m+abF
NdhLRVbX8ZfRoyYTOS9wQav009hDadDsTSTLhQ0vxVMj3qnIOSYS03Pyg6uMZxvf
9KhVCNqF3pipZpN74p47eA7JWzxcWJuqGCe2gmX+B0Ibi2GOfRqhOcoa6E6/iTuo
lMBIb+5N9Gx73lY2NEHE5nwYmwhFli4BKYEDrkwbre4k5RqoMIeZojvaa8ugg07/
QOUGgwsfqpJTPsYxNti9utdNiR7Y7mJpIBRdICLdfQTdkVyh5iHSqpH0ITFpmJCO
gvlspAMsNj5bvy8+e3SFoNZP4P583KFFUKdzcoiq5kFCSlNtQgIIA9hl2zTzf99K
d3LPBjK8oH5bLoq3Rro20bepL0IH993ixs8+g4Re20S5A3S9f4f3eormQJeXlbUN
7NzhgNwuKEhgXi5iVJGmMTOEATbJQ8FZNx472L3JFZbGe7WmGLoRVhctAnQKvWkE
k6DYZ8TwTISgy6ltnLbfEQBMOeoID+XqhrO0aW/VbjEqpG6Muai8CTkuNuwimsLl
/bXGG+FFrrUUtJAgTKhblTNRQz1QNQWR7YrtrxKrkREhoN2jptLFyP/VRHorpxcj
cNP3aKSvHcef+5R23Q3oY1SG74NgOTsOLFjLkJIGC8fyGhD/j/3Y4wfgP+/MHoEq
FACnr8UuXk0TdCq+FzYGqFJiFxP7PVufoiIfSFXUiRJrYlkUJ2r3f+O8VCoHXuwg
/oW7bjRw88ulgP8ZU3nZmaxRh+dwD3wscvsm2wEc4o+ZUjVJIshBV0hI5NUNBnrf
zKnpyEcVKxoBK9tL4EVJJblK5J6Y8jBIOfYxqhvnq12WiAoK2uOFK42zRuPVtOkT
3ISYvbIoKJ4hy/BcwAyf+iaZWaldp/VZVw00FiP+uLpJpV3qYESOGf8Gyq2xGlYW
nYBrEzti+zkOhYz/eZaweyWWx+23cbtTldGP4cfKd3xlrKLANYdVR4GrrTYCa8Ie
FZRcSmquVQqz9kr2zDUNQfLBzVZKnPEVzfxudAz3UVLNHaUgBpzm4y2XNKD858XX
CzJJiQPwnD0f52amxuHeK3C80Qn7Y+9JY707LSo+SAO3iPorN+QfgzaqvBwUANWm
hX6pwmqsSZU5w2Hctqzcu4h+dTMRWs4+4x0pCqsGbjpqgSKWJwuNm4FE5zxTuaG8
jntgi25U74Ke23OjLVPAGdTd4V1w+9UYZDREYPh36lx+RY8xG33rF5i59BoI9wiK
j9N9W1etgYvrx5cA8LbX/27ss/NxtAdEZiO3TQTWZ175w3JKyrI9x/SymK0c3Ehi
ZBXN8FGkWU338+8iOzA4+uIxQFmNITOO+MoCpJugm8KqTm6nVHdMfgUIumdZS3hB
jfO+Iyr7lQY/61a3rOeZVJ4PkWH3IydjOI2snjMeAVMCPsF6yC2tsgITJrXtArtN
4t512J8nrlObBeo60N7Gg4JqCrLvHgQbaRIBI/OpGJASwLGoz/z41gR/S4hA5e4I
XjLCti+e/wz8oFs47EAVW68DHlpwzb38c1E2JfIiafm+P4QXBFtcys4LznZKE0us
rBVu7sw95RHheTbUfDIRLSJQEw0o+3z2NY199J0kT+NKLUiOuJ5BaYf/AyIb5tk9
FLB7fIKeCqcrkV74gZAVlK5Yw2dacfmdwFvN0NsTsW/jWie2h2I88w/F/3Izr/lZ
Cvn7ZjUCdsdvizS/K6p0+rWaqxfcWKDa0L/Rq9nUUl1JyWfXEY5J1rsTke+6fxF+
bSEJWhjpbxt/XJWCjSuFwtw01C6xe3HGgmQFD0qDz0UDKrTj+h1b98LsrSutjJ9L
6soBB1ZIJ+bWl1pTsQujQ3pCmDCwgA73grT24oikEzQJ/FY0BSt+gv9uq8TEbXJK
M6pXcxY3Jbcj8Fh3luZDEhHYCCWtftVUKU1tQPgFLm+sqpRWzr4t3joXIUDgeqUK
Y+x710cLF/+dwnihScPEPafj/vvw3cuOLHA7FC8drfCzV3eAMvyhpgn/yH+p51QY
Q4DdurTsMRKKtEiRc1+YHgJsvedn1RvGntMif04Irq4+iBoa+HN5G05nkHmFGiVG
mw6Hycb9NZUShQBpbi+z5ya3rMyOxHl5y57DyuhyRwtWM1VBC++xeRs5vEHKUzMj
nCkZqZj+3KlQCE44Pcp8bDnFZxRgmEwnJW9Q2cUzue1zJT9w+ZJaNynErNzEXOax
UCU6/5W32YW/vToLSnHP7/NB0s4QvfM4dCPGTMwgMENx2tLVw9NWQS+i5NxBYfXp
XUu2sFPm/sn06uFklN0PQpQzh4zuPRLHGV0zNToZeJR1dEUJlsv4KS/Cy9Ns8LTC
79iSy0r4/59DE2LQX0cKJ3QEepBpJgQVBcDSK8LdVZgcaXJ18Pd23ZEamhEhGwej
kyn7cmN8hw6daKLN6j0qTZ1KFwZ+fjSFknaT3dNgii/pQk8xbXFnuD5fld+iASDY
b4fFpi5E7/agNXg3hXjaujwm14Aly0zLW3ILiA4ekRex1xYlqckBkS9xHC1UXAMo
+M1nr0yi09Z+8U8PYDZe8jVULIhJjXiZoLfU4PPeImmy9sDzmiRLuluPD7v4W8Zk
Gb/xH6jHeCK2vR7NcV/OlBfNPrtGPYvaN5k0iA4mvJbsAP5bxgtknJSIFs+CalFk
9hdpgcrdZ2fRJOa7guMXHX/PHLOp6sDenxv4jah+MdxTscCiq+zfR0Yy3D68mtxd
CW6wVxFWYyr0JhrasiY6ZuDSyvltXHQVp5wvzKk1gbYn+tvR+DYBSVQuwmHhRczX
FCGjHZlTDz+U7cXrb0KlJWo5TvcEWf3JiGIYDIfpYK+J5lz9aGt6WoIHmpQS5LgG
N10OMKZy2Sm8pWjePhsS9wyXV8yrDERf6XRFElyHdw7UKqYsGkb3y8Wk5YqmjEnJ
a2rx+PqB0E6jzwpU+XybuJPQTPdLi8pne442I1fAwGu+bKX99ZCZTu0/SVxvWo01
Diavz61cBFxNDxuNqj3S4bgG3uG5q6RisTTKU83nwdvZ9qLug4tbpG6jhe1AxOaf
LoK48E5y+P7WUF3y8IjO+IcW151Wfwi37M1KEi435/VN1EFy7svxOg2x2WwOtDlp
xB+smwixbAK1Cpp7Hzuqv/3zEFRqdoiE69DOSdjYa1MXTLdkR8hgQ82RxJwvxKzG
sXHLV9caCw9rC3P9nB6Wfeuk1hWnh0kv9wPV1N9m1LgwExWFxgCsVXvAhTnRe6Dz
aFMxGLdfGWsqRvftAGleP3YB0CIhW9e0N6njQTssevYfdPsex4cEQtdFfWxu1Eqy
R/Np7LnFqlmlIs7479FXU/tsBeqKqXbnAMYv7G7OlPhLW/nhnQhgwZT3KT1Hdcme
b8Yt4Rm2F+dbCDVosLXTDMpde7wIe81i3FXVwvpIN1UlUbiVZxpTILc95+xDnBdD
vz+2eq8DNvuWIK9rAjsoIT/sPMGWJUqQQUnhJ/qBuozE41UOULd5vyKuKZmRA7Fj
cZGvwRf9eOeFXvEYNTh6pjW87llEL1d5ETDWVfpNa45fKJabANfTVG+Y9m/SJcby
xtQ3yasCX+ArJxenFmUnqtCUS1ewWO8sltXZBWPjlL69G4mzSLx7wmmrA/0CggCl
DJFLjWT/Oio9mjxKPiYHfPAKPQrJucIYWl4xLIs2zClN6a6XoFdrF3BXiTy3m1dE
B3il8/B+zSR/WwdUNLFFmeeinELuhA7sNXNZhTNzx8Z0qm0+5DfqQ/IXx1pS6gF2
Fi7DMKq5PI+QdCUyy61TVLLUZyOYXnqz0zoQP1guQZ9dSgErbwb8dNXJi1FjnKu/
yagxyp0GjD7wFrb9HIwjKWq08DKPL9MvikIzx+WlElibhKGeHErsvGLrSrwPD1Nk
+e3bXbtDpBf+YIJH1f59VisiFAaCoYY3m5uGQNc2u/CMKS7SFCpvFM5TJYhAt1WB
mNkoPbRRUrLCFsbrwbYdZcmfqOlNntPAX/4ErSQRfu9yf+vmhTfLdYoa8QCSi+wK
aEDcwZhTzwhNf9K9kNSPH0+mRK+aehWs8/5wlmJVOdm7n8Thf3l2pBSNNsXNHVtW
c8wIcNvIk6J+fHrFQ11geCYJDxTaQnCZ8Hn/qexSOZ7Bm6sNOeE9XECNfcjOnCEn
92MkSQXxY9fuFkunKhU5z9VudLpNORfoNpVZCH71As7CKo4HzF8wjZczIppgrX1T
M7kblP8zRX2d3mLUOkCYpumkKL1HuamX5EM1rHSwJYg3Tk5ksHVsaadFOBv5CXF0
R5Uy/hjDswQU/C/KRMBXvBx3kPy0LXkHphHO+NUcJ/KllHIHletEgv/j7z+b1lr7
2gjFJ01HqFHuLB4M3IieNnL7BkAsuO7avn0GR19s1GBHqoL6RpT2TTplNHBCSznK
KGG3EQqUtUbTIfLRGK/8j3Q//UoD4lnZpYRpncPy6jDUTFvo6KOVBqkeXjxhsDMO
k+nFixTZKQzqtQq6eaJOiO28Rqy7ycZbe818xFITTw02nEpEE7/L0UQuEzr0i7Y/
XDzFCLpUWeik8k7RV4SxxXZlM2PfI6BUoHVf6DzBUbju1AC5dZJgCMB7/4ztElma
tNHewYeC2+ES6uIN/1ptgGHtNiMgkbdvfPkuORh0PQgLx2O6L4wmpj1nX+1BddSz
AhKvUkOEjYOll9WfoQI86y+Vq/Ur130kp2zHerWchdRrqHdjCrGvJdeII+i6E8Z3
SZ2VXabYzzGHSe+dxri+TFg9sYyr6pALAva7hM1LeZS5398mg53Z2RwIfCpIHB7O
2CL/tL7vGdrrxoYFEBwgbE1k/p2rXQEGKDi9St4uavGDbL3dElQyWQhktRngYdXS
ppFqEzRhKvYd64BaQ399XyOvEJHeFEBK3GKjftYfgbKUx39WuPwcNuDxmct+eGGB
wwjKOas2lZF/bmAPDK8EhdCmuOJRvR3eATX2KtZQFfmpuRitN8nl07iPqWkNXRzy
bWgPF5eTZQiFlSAbnLfSPJOjXeoNWEMLQkMHh/IAxQ1ynRQaaF7+QXNJoLZrgx00
2N4GiicwqR17mL6AWlA8fMgqXuZWVfjHswK6y0kAtOQt/JSettlGo1hhuVEzAYS2
duKm4Q1kcKkBcJVIx9u1PXR2Ll/s7plUWeqinvLwSm9eX7v5sDHHFCBuWwhz0ov4
7aF0bKnob/Fo7DqIaD/3kAFDjBfqAkrxYfhGCYTIYzrmmZE+E3Ynrn6/iZ9JBBEC
J87VUxuF8m38zcoqlRVpKsve4S+cQ0qk/plat+XVVUI8KZn6URN9EWCnkv4v9cu4
ZH1/ZvhcXMq1Q0h6kLUL6QMSG1Zsmk5P9HpB7PPuHtJ0JWDtnLOn9wMkAupW+2AA
YEF/qSbpoEqV6BcOaQzdxQSb4fw3kb1im/y5ICy0LlbXhfD7GB0s4BVyMmdPPINc
cNT+AiORsA8cQUsW6+cBVjjeq5sBxvi7154pSvvsLtPi8ciCCBw9+NzZYKN+qXBN
p4L2JkX5x/Gr4NoZoq/PxiVLxSsrvIYGP7QQBkMh7CjJCxOup/+Qy97U64pCnMgk
NuKlOW9uJeYvRpg1Te72NfUF/ueqJQTMXB5hwuYw2HsPBgE+do5RwgZJk01MgYcq
1SS48rwXNo23+fSTl99CjKWrTctwiu/e40Z1IsWcaN/TPl3QetgXlLKiaZRTkBJn
CMph5ybxOYYUrdnhkQyNy5eZgx09y3r0xrrmKubE+T4AOrfYUBXGbhiwQIlkYHeP
6r1oc7uQDzzA26WjKZ4BdKsu/1wSOGJkL6swMiAyXJdMdb9GvN34RaIspsRH3srU
xGceV2CuGtyBECK0dp1gwYmEtDUI7Kh13Q/6nzsnbUr2hoIXO0LAhzIRufDKKOBc
5vfWRLPyGtzla8XVZqazaWsZBkVqArk7YmwwGSCrrvLfB8W1NrH6aKVkDt/u1hUX
GvJcEuXr/zKVfN+xDP0vYkZxobX4Q8nII8fe/XijfRc4k/PF6GgTrLFEde/yEIhR
mBG0U8/2Oam31oem9BvmQEmfmMFqg+5zq+jI2eVZAitNaI3lTSTGddHNQP4gMBzW
uvtv8+4zIP2D/bijnU73+D6ZCWhs0u27cnFJ6Vm2wmrexnJstg9EoFemDMOsFyXB
+xVx8UL56N8Um68Z/AEmjXyr9J6AFO0+mjoiM28GgXoouJ6B8925V7Apr2BsE0gL
yocVNBad3N3WDkGa+Cr0F5IJa5exT/fsyTy0JKcDQwrYQFO0ztvLXusXLMu91/oT
pLdCc3JJ38jZmo5Ymgh98YZKrRdpdIOLcYz9UU9NcD8X7lzNb9oVvIHjy6d7zKfB
j5kEL2oA3at8YGa4TuC44KitTOPlygwRvOJd3at15mlMCg0GyinkMIP0R+qGE0eZ
6ewoZd/xKT6A/BBxFUPVWMnHIipwwik6Eyf6e2SxyJNOlNcj54xI44cYWaIh0jlE
bjG5oVqV22RNOBVgVbUNcQMFNC6RITLsxQBEWJWZr6z9mvrXoklZ1bUNdrjFhEM+
eUtG6RNvkWuwBLRtYG6vEwLFY15vbhk9+uQHZsj19qWXQ7SHGFP2YpPHmTwknzIp
f0gLpFDlyHk13JJp63bHkIc2vHRntViWxBJksdd39Cu5UfHaW3Pk1wPyQoLvcyG9
gmcDTeg0+LkCCWMtuTrfk+NDLco3dD6j/NiYWLr8bkWLerMISUQ9DhRg/z62WK31
NjR7z3eyWW786NTDspeTBWI8XQwv+sDmsYzBUg5TKm+1XAutr5rUcPQHHwWwR4Jc
YQEbV5zHzfY9XtakqfWaUOODnYd4zYM/1dzf8TkephtT8zws2WLq8CXomkR3Au62
tHkXxlJPs+2IvRzX6BHWxmkTfj7OUDWtmqw8y/WJyoDn7tKjLDiLZPYmezYLxGci
vyQRCktgwKb++8I/+fdm0Z3sLl3ftlfCfbIFjnVVE9/4h/SvNYabo/TS81pg8ncW
1AWa7De35EBFHxXYGJr7/+JfdbiS7pjT7bBSV/FxtIGWwft2tzaSq0U576HYU1IU
rDK/oWFf1W88grfT3UOYhUQkrp+qYwqfY9fcidAXkPtqor1eMt8IgwZRtwweI9eY
8o12xgvwkhGpmAcoOe4yeC3vS5u4v4thsLRg7wTT4pLOi9VQZAmCnmzZBqzPs7Gt
EZrFprfFp9q/p0dVAPk0bjMRyTUcZNkKLlrrOemnUtJWg8UsRc9oYpgXsy7ndbGR
0IjjO8ja4inDAqLOPZyWJDY7+mlZOcVKQt8JZ+zm6nQq8AtwAHvOIwPEmIMcbpMm
h0zQX8XSGlFgxjIPB8fuDWyhrj1CdcISutX2MMvYn0qlrK5ESJFlbz9Pem7AVplp
zZ+tPVnIDBUBEDLS6e5JOkdWGrY6aU6L5PcLcHzDH6cxQBxZWQldf3f4HD3/65mx
of5Zo6csOIdxvTQ843QfTJZOib60Fx0uetI0Zvbx0KTHi8NRjNEeicmttu3F2W3r
g2Uvffffgfu4oViAhE462NPDuWeLSI6x70sDXKOe1asU3kw8v/HjFFQ42SNHIoJv
foFrAbfyzQ/GA2ztMol1odPaeEDXQly+Zg9gnPCH0gJDWzqAbPPyXDd518XQMcSP
DINYFVcLzTt8v/H5UeMFrhBlkw/s4hdMX+PyWiyHNx6OisWVXGL6MdCeLA9eClWN
cq4ybnjo0qud8w96bEgIRExLhxehIsE2GMTbVM0rirHZHUCfzUVx0NRfucq4ti9s
MHbQvPVmQPFRxnrv6MhWQDxRBbDy3UnngSWCBVFSWYxNu+0kunBahdXyHhs1rs2w
MFtQ3B/XfvKi4ZHI9CI5V0B1DEy4azr/H76sypOF58TX44RrJKqlhY7Kr9Z5QaZw
0CI3kILlSrVMlXEDI9KCx5fRYJpRhSQh6wWwuYdRm6cQkjsrrBAP9GGDarVyEiMO
+c3bbIxRF2ZAlRYerdo4WkVWABQiBzGOda6pnaB72lSykzC1qO2L1qimoYmyDwbu
s5QoK9OOsGsQ/+EgQ+SX93Ki2tmuPbYuTByLLEVH4STM7L7xYPxur9zXh7bP1lMX
rh9vIuupzEYtvCt6OQ96yKu213EUKRY62WZOayRg9oN1k0Xgss9+iHJ3zypecZ3I
9ICv1AU0pWEQ++x7jR+dMlTy+imyLOJeYmYV6/j9r+i1uMkXt8J8bTzG+jbgNvNy
jvVPXehv6Aw0PQu4w2sFROZQXEBrYj32bAiCyv7pvT/cvkRFvcs46vlMDWq746D3
7RoKOrGgXO7JvGn1s1TzYjRgqB7IILDsS9XXAxnjqk+2ohhlGzrLE42LEGg8iSR4
yJ88oyeyGCQ2GyzDO1fS3l21isBRlL5mj6d1gOixg7vomi0o+A4M5eRzGJcGidz3
C7O9VhFnzJ2KT1jSnbq5bsh3HoktCrNsqcUrO7YyeSEM0McwjY3qXR93sdxt1rM4
CLf/orD/UzcpEe52QSgl/KIgJufWlZDA9g/b3u81UYoEGXx59cvAC4MB4OviU1u9
9+9q9AQVyMqrnQh37TXfCQwXZ4xKlwIwa0UYX6kV+awnQxsGVfDikMQ8bRLpISyG
zHohzjsT9v2ngwN6WaN0d8WLnS+EfgTGkAY8Loak01ii5twKWykr+toYi1vmOwJZ
JTiwhJdyyvl7/uQq5zRgVvnLDR3zIUhgz9XogcyAQJ1qRDjKoWGN97pgMSeFftpC
FFr3iLTUm/+Q451JCsZLaxK2sQtibZD5DElz4vuoqJqQOxUpMof0QVfaoPZ2dCtE
aonYK7jvDUeWnQCLEveZwwjurVwEQHk0G8khXhgY8cr96VHoRkVlUoMuVep87/wX
M7H+pyqPXaMXZt9jA7hwRJGMoAHRmnfvsbtQA2CcaUnOJXaBtkIrPRQ7fn+MwieU
mM0iP0+zxqQAkFxlbqJ4N6M28rBtQQNTe4WTsAIkad0tc/ZT1t0/09T/mDP7K7DZ
YwFmIjmX61FKyPYw1aAkj3Qo6821LF+ka/s8Ah3u3MHiMo9yim5HCwE1+1aHoh9E
NasjxWGtJ38I/kByXwG/NPBPQ1aJchv1YQRdfL0QXnq+xx9RPuWB1qWb/bMd8IGW
WjWMpndGC6MkbA2DG2EqEu0vba2EZAH3nMGJuCnNIeWHW3gZZv83uopEJJM4VA1l
6RefcRDj5db/jd+yHbh8ZycC2VmpTsN/EWA7STCMSNdlR305g/O5HzzHm4EdeqVX
hAtFmM2qIgD1F6m/IfooRYLbE62NfMe9Qt5spmVFpXVdVF7xbj2T3+/nAKOG3nYb
t9jfkah7MUXGLNM33TjWQRGzqDBq1iZxwLiEiOKY5xnoepuxPDAmyrWXrWbdEQyX
pbsOnIq8RwfU7r+ptVutJF7ZQF7mXzDgTQ918LZ1wFEoc6YCbyitKjPwRybdgkOl
0bl6Ma/+FJdZhIAkVOSw+dvqlKB7nKtKVFjYkOTByjO9TsZRqb3Lp/LxWppWwuab
Ynp6Wyd/Ql8m4Ve2I2oFuoWqMl2sWLJkimTdBhLN5SfQav4nuZzW7mElp2Ke3THT
4O1MFAOLoPkAHLZyDOUFqLw0/2569ohpcugWgCjXGNCs+TJ9G3yu+ALI7wdXjMgj
KEmBqecJ675pXvoX7vrW5rZcVkh+UAhWbPH0YxT6rhJlbGEk7AwLjAnIBeAs+rd7
K03z5/E/bdOuyprwxuzkhhhIWXrVbIR/5V1U+LRDc0ux7Eg6tBecTYkg1NibexAU
gloyhgTUNTwvLC9ZwpObEiAkJcnc/frhD4C1K2cRbmTWnHBCDSDD8gb89EcWGS53
fEqgg/y28Jbiz/h6lxpmJ2bnnbGHWI+nyEqfV+uyk5euuFrGzjTLCGlDvXeJiZLx
3NZEuv2JUHdP+sRt964aqS/9prLP6X7zzBvULm23iqRl0yGe7sBONdEXMVWV3fBi
1+Amw0p2k0gwo7juJP2+6tAX8YOrXLHg5BrHus5JirvApMXm5hv/I3IxO/XPq1og
PspBXdKdziQce06KKp2lIn9Qw5NHAh3lKZNi6wAXcIDv3SFNIi6F1ge9Fdy055lf
a3XJi5gFJ8rfWi0qmQ0+M8uWbTlqEmTQz2MyN2acN+cza4b4UHNlTbejNfhDF13i
ZVwH4MPeXp2wylkxZMrqKy8YgOMf9FarVuYfSIsEzSGf9z031izgoKuEIFBbTmns
7G6RwznIG0PBimMe6H9SpLda3w3MLFu3mmzhK5zIn2u5xePMDAIpMLf99q6YIdk9
fxw4Hb7XlQHnOonst5K2xR4KwGldobl6avOme9MwoZsR5kp1Rr8qDJggMsc4v1iH
FO285BSNMJfcarQa+TPiYX/ow5mGCUbz41C6NUrcjidWWVYSDn5eDxf9pFmRf8/X
WoMVTqptCnF++taOTXrRqu2nls49RuQuAoaBnk5RZgnUXIF7bK9B18iepmif5Iji
mqcah2D/1cGBARqiCkPJipwXISgXj9D2cMCyi/eFaZHPV/Z8inUVqN7fz92DUYX2
oaR2v7JZy5PsM82ion0TVbChqpYZkaf/dPAxSKxshyfg/fYB2IL5iMuLOnFJoUbC
f/AUgR6Z33Zj8eXuFg2yot2GmxNHQ5BMdxus7o2HP07PoFY7kXXoHBu+SJBoLUbC
9/2Luu0A0aT1EwODRTnrfDyGjgkENadapoUBpLNMBDkBdlJLyznwvMgks18v3XIr
+upcf8fwLPeJ83j7S24A8iYVeraW0HiFpKM5paYLXndQhSekLei5IP3nqDOtqb4R
Xzu4zjOQPk52gXqA99R9tJWI1GjDcqgwALNfMw+cv5elvfELhbr7/OXqeedOdsbK
uwLSUg5DG5WBorG30yoWAfSNooribD2jpOIUw6W59cY5sKHU3hCyOdbj9NEArh3P
k+M0jMBiicsmkyGtk/WG5xt5ekx+19CHHXzCLg3Fh2govfNRXKQOQwH9K3AXpy8N
pxTLc8Y+aeU9H6PIIqeiE4QjsDMfGSOc1kuloNjK2ST9A/dHJFqSeqf4fXRLvtkx
WAv/p8gpTO987yctPgQBzT0fvDn52/UP4HozVxsN9XcNI/hkNSmqabQjxH5H6Pvp
ovFPEH8+sl5BHP+uXRA2GKVplCWkQSdHBE6LkP+8gytMjC1fYqWOrX5SL9pyFrti
DXoyGhEveSOoIriC9m1ThgKXhECwkg30VoSqZ9hOwLi0FWt88pQ3WqWBMGZ4rYu4
1lgnhv/MDq5EeAB93Xzaw6U9bmldm4e4zKxDDtFDNlgT54xVCDMjLU/JKFN+k4ik
YDgcIb3XvMWGX21dXzQfuJ0B6r8J4QGwN8jcZD8ysMMsQd406ya/3LKB7Ev0nSSx
en9O//CGsMFyKvD8o2KawP+W142GiaIw5ZGXhobRCdalToP6hRU7Hkv46YrZ3PRe
9km6WJ0JWVTgnhpqVQioiHpB2h5mqsUwTptxSbtp4afA7CtJMfnqJ5QpDpqIemdF
TXtRA5WEE2KQjUjI1Y86izlGN4TRSFNpm5JTwkRI1Nv6GNDWfUnfXyucxLWhwBYf
4FqnFtfeuv5iM4iJnyJE5CFv/0lLFt/4cHyUAz0SXOPEfq5qcxHdoUQbcsoYgD/z
n5NWARh31tmvGkJlat76hmDeIGmsO9GIYsb7FcS26OaYcnylK/trw5aoEiIZjWDz
PzKjxSQWlxzEhjBEn5KiiffoeAccmgvpGMuT6tDk5CtgisoBuLqWnVuCtOU96jGi
S8RLTfa8Q86R30M4EqBYWrJ/Z2xbqkSlgsFSLyOJlfiT2c/61RhEsJwGlGaiFbKc
vabVHuO3RGYIJrbDfDDhGF6SQny2oUdY+PL9/NunzkKlsyhs+sZ0RuxfmqZ/qDo1
7K3/HsY+ON6Z49sAFK4ciAqYKd3B8zdJvhpDEA/ae+1W5+XLbjD/+at+Mw/vmJYc
AKDaHWIkNYaIszVYrFKdw2kkTFqe5wWjEwFOziMI7vPt+A924KqTxG/LLtt+qQD5
mx5WUmC9c8pWjNPSmk5NYrPmX3EWH5bWIlG8wtCfbqGFd6zxwU5wzGjI962pawx2
Eh743r7F6MjcruwDIMdAR0fL2YUkvnzOdnI7qn/Le4OXJ2KPpkTksmOFk4fi0hs7
x9+sFC7QOJjPOilzf4f1DBQikUoYMgL+M5KYdzavbykUoDXrjLPRG+PorwOr2BVx
DdhxiznkfwF/4kwJTl4Yhep9tuGN7BtMcWsB8MicwpiEum1UugAwCpT81wVggSHu
42mzxEFjUo02A3YrxiUIgB3GIwNzvnfzZy1jIJJmkTvsx7rPlqG9nXVp0rtI1S+R
ZAWpLxFc0AGH2B0qOCZeFpCYlTovd0NAaVV7+kIawmOMtr8fqhT8oQQ2oPIzXSPS
BZmRmXQDjBlof41Own1abhyVPqfPcpH958lNsHiu325hwqjFSILU+z/tLrhvxcgY
/qLK9Kqg04hodVE4zRS0QmDP9a1ifMmR/RfaQSxi0n68sozEX0nXEbKJP+YjCzug
V3QLEhzQLm3oy2MJCT6+f1+qo7k+N6gSrgx3eyIyAgt5NXdoSb7+Hmyk+XAPbc6Y
ORgk2TZrp4N9/VGVRmakc7VTCX9JsPgTEPvK4XXerb4ODc1gKGWjNNmHzbSLTteQ
P203ahyDbkqvPVLGVtt9ty28Fh8VekdC4jG+/31wuoE6n44suHmlXN54V0W654IQ
BsW8Hg8sfHEV1kHxK+u+Y1KJMDvE/wJjkYfyf2iwx1LoOeoIo6199CgTrh0rAa3R
Ioy7SSNGKBq30vTgQ25flk1S3eyIWiT9KVHILnm5pPZzURA2w9AwtItpsgjr3BJb
Z8FxAotwsWYJon5G4+RWl+RTLTTVAEnOW9n/mToPMMhaBHpgYcYjwlKUoe8K9r9E
857Zw+6rxaEKWCVOtDsnbJW+iWkixtgdUshGnquzmYtIDJl3JWgKfnJlsC257l10
mDi3GuU5AQw0QiLAm6SYslovLK9hdrmIR6mLA17x+khECx0BHBKkwmPtFVGnrPiV
MdExq6dtij7w4t2MWZVWSimlX4VZfB8w9TEIt55uQwZc0tduXXbcEYOewZwu7IOg
SCaEZpRSqXSq2Yjl7Nq4KxsiJwO9QiwPhRzM/pMKQgl+YmFmWrLPqaG/pXuYzEBI
T5OcypZlL+nDVaatYZkoSC92HEg97dTMtYnMpXF1HSbfODDuloGsFMNI7n4+i7Ib
W9XjnCwDjjUPmc9mB1I89nWkz9d/vzCuEAlaYcpff1n4B7dGMH80hnLCjJdQOI0f
KW018VdVXIaVlFymyxMevuibJSrrMELQktJU9++mNnDiTvh6XdqKZfxaZsHUIzla
pR9XGw1YKpQ7M/LwJYxehFOsPBfOaRi71SphYQc1dDPQgo29gTIEmM4O6d5N1Wkn
UqPEzwq8OAvvwWnfQY4+AEMfDq29QoEy1hG8vgqvEv/9+8lEHmT7nv2Q99UHFzRp
7ABrCn/Qg4mp2HQIZKofS0nsD2qjgkXsCsz4dZgYGJ6hJkHQ+YLuhe/Zye9uGVuO
`pragma protect end_protected
