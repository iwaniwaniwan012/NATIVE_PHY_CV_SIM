`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Bb0Bht5aZnNYZ8jtbj9W6Zft3GSsNVOZLX5Mq8f8U+FbrnvyFWfznqF1uqvbXLJo
//K7P9mDUZnYIti7TtMak7FA2rC+UxM6nWMv7YdUldqMAGfIUDqLP2i7P78vhSkA
dqTwEzxU9HD3FRRSbx4bYXOsV+sRagG03moXGXEJvyk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 123904)
DD8qdaVDMqIKB0i7PJP09vjsGsKY8FfWRss/+IPtODOQfQoz/1jSGgZlQGKvTvKh
LeqguRiEAuQWU55ZsfKElQYhFjVqCTynoEa5nLefsl0CXFNdzcMaNeKFKvkrBYrG
VGlY1Zfgb0eahfqt0bxWs2nNPjZQMQDPEvVU+s+PGnllJ41bqI2JpFcpNxapIms3
ZyjMiGbPD0qSWaZrH3FdxIOrO45n94cSs1aLd7eh/T8N1tlFzEk+lB6X7jaDWnqq
tCmPgBkbA3Zd4TQkULdHUCNlxsE+E3Q7hLopRmOsOUE9JIzwmCxIA/E/sp5dohV5
P2G0sByTenTLgqftnMZokYIBTnWIJhrpS5rIWw/Q6N0OhN2Nstmo67ZfWKDy0a9E
IH7lTmf37of+GlEPV1RYPO0jIJTQvDvM2TROoy/w2UuRvbmowz2oHlEbwYv0W8Sp
pnSWNn1ga87Y5HAzU3crhOwi3YrcjDRWci33ZFvU2ohz+I9vD4oLYLesxjXIWi7n
Su9GCbvbnlHfaNpFewISK/WIlQmPfI4fKB2s7kDwyGWdkQMTX0LRQ/+3n7phxxEe
5WEc7Fd3MXjGDEzKNFSbtzEkcIpfM159WXxukVgU1I+sroO9CPO5w9H3ghbTxOBX
M40yqjrY/wklCHFLjVHb2KnC/yV1aqbqi35XSKcpNDBsjFt7MBJUhecv1rdLi6DV
DSt4E8lUpq5vRYJOAB3GIJ6koZ6uTUL7vmpbVeZ9gGdF6g3AJKwE+48SAxGJvQTJ
3+suoATO7aMSUYCehisK4QRsz+ZzZvGwlPNrhVzZA5nbrA4aTiSFnScj4iF0qWuh
p7OvRX/ogrO07y1W1ngf5K3z5224v2UfyW9JX/Yu7MdrfMfvbE42DRSG5RvDmH0K
GtFsS0HyxwbHJFMFlv43HpQx8XiTPleje4Ijwm5rJGAUhlk52nifJTBU1168TLJN
AgalhNL7uw4R5cKXf0jUYMvJ8OzmFxus8jDg2vjP0kOVsrhOp0BdPVDFGVAjAIoQ
/2oLeN2MsgFuZ8PayIaO0HKNAc6m6eK0Gf+AlWE3dE6oB0HNy9m9gYKDWWYp+m+D
yt+Gqylpug99x+wbVaVTaOwtXytsZDc1x3GNpUTPT3ISUTNBKvlUeVfDarohJ3vY
J2UOad/5HrLpnLCQZ8ni4zB76YE8eidZtPGglWu4e/OlIfmn0GrTAHmIzL1t6wt8
SfSLPGfWeA2b7YCO2s7XPoTkRiha99Mge6KyyLxM7ix+JEmJ58c+viDAkp8QpqZA
jLvXZp56cMS9VZwT7qxC7f0dkHQ2YxgzBE8t/A2IxsC6S+H4RvHgdRP0LPrIae+I
crU+9zlfdt9TV8XtGh4BbEG/a0GAysmjGukg6FS1VGbzFGzsbfWBaL6NmQig+FEo
MqDYmD5pUqwrbHrqxv2nNR5V4L0RsEuJ+eCHn+TBm6LmwJrOSY4MIdvzNyLBIFUp
hGSXGHVRxCxjJo6+OtyYAIUepuGzWDJXvDH6ogfOF027NjTlIMIDyqgIjizKhitg
f2+SuzUoSYABo3KzOSz/1mSzD+Ow3dATcO8eW01mb3cIiRQLfg7MaqiVSiEstinz
+IbQkfKCi/9sQsZfwPOWBpPrLboE1wAk3/2/5Pzinav0RrfNcR4ZKEQza7OJWBdd
5uhQ3pEiyxxDj2kFDEtdXftR1zyOCq1BTggPKLqLI7RWq7pqwjhyjY51kpmgKgEd
mz4syTKOC493cUM3l1plGBOOBNIobjSJVbRzswHIdgESG8PNw9IDvKSg06Hq1xuJ
u8jIubHci1jj4JPY6UHmMmGtT/P18Rtr+NW7+VRs62Wfa02NxsTylMQ/61gL7ozj
ZdF1KUiYMus4/bIIkMtMCcys851cGSOIJi7LdjfeHAxj5tVVRvkNdLJE6YIWELdc
Tuk8FHtCDULd1K+JbRexXc2pNk4lwPfSuBaUTYcf6cDlpLB8LOblQ3ZLJx/qa96b
pJ9Hi7HHkovUhMLRTsaymmTC/IlwKmfi7brSvw9FSfFnK/ZEIySiRg/Oa4aUK4vB
4mmo4xGApQ2nV8KdEtMleB4Rn7kUin9lQj7zW50NTWCKCZGIRNSnij5S84EPOKt1
I+op45bAU/hYVPPTXrYFFHBpX+ad04TvT2KOL3d+APpJdTX1Wi/MFaaPMQLa9zqF
g/pTbzAMQ5I1Wzdc2X9VzOne9GxL2Vqg5uaRiPncpCsoDHHNHRb7f1b9Y+fWS0N+
w75l2/lk1PAopIjAJvymATDgKVTtYZjWdoDdbySOx7AZyk+0dxcB++ZWdy/FQL6J
i+nVkFN+jGdr0yYEzsfmKDQmX2Lxz5rHXA9IiHvgDZayp5J8GJl4n+agJH6vbhQH
rVOnk1ibrNAD0dN91UUF7KIK8luG51DYvfDIb2SFnmctjoYh1Al9WXlKJ9fDW2OZ
/jCoe9Oc+HlMMWwz3NRqv2Ya83qxt32nLs7F2dxNky6XFrY799Sj0pxIaTDRtsjt
P2K/TN/QQWZSv8rDEmBG4Zrzxr3f3PC9Tpy+pOurYHObWsLn81/qFEFyErAg10Uv
Cbg6W2xFM0vFQhMiuE/hFKKROW5fQzFDPbZXa7dC00wte3JzYIIFTgu/Zoz9WR/h
c+tTrk/6ldyr2GcWpspWQkX64bCD1OvU47gSVOunbhSSi5obtexXBjaPlijPhqQI
BRN/PDt0pMWsQSLCeS10LaUdeMkZs5fwnMCRnpPO37tU3XhuVvKvujrtO9D0bXoM
gUFGiWiyMzyYwUkAZQZHl7TNxOk/w8zhZnf7wS5Msx5vZZiAYiqCBOlgbiOlurMj
HAoTQtPgfqKmcLoeoKm6blj/7rv1xwZsvhsel3Xymdzx0sXOhxjQ1zmQXeJ0MQ8k
ABA5CzO3v5ee13gbhn54pKBX/fqDgE87inECN3z3mpPG20PV2soa9Tlnlt9mrwuO
Z4n6+jdmGITBTyDf92ANKXSuZH1fJeAutDiol85Od6kI6iwOQpRydNpqZYea72pq
zn/qrYcy5vGufMIUHuCIdxG6r7920Rc4SU0hZ/vtU8TrGV2Vqmastd+f9W3fDWlQ
uKDHEwrvr56Qf7VYaxXTOxy6nJIQQ2iHuPNUgtgV3RcHrgFLDKsEXeculkRT62jn
FVhHnNWFDCDX5ddS7u+EZQWynZaUdbN23+rXIfwpFkeGxMDUB6y3OKT/fZENzuGP
CfTEByZKxwWGLsm6zHmo7IMjJWDdBatmUZHqjzNx6wYvOiNg+ZHV9QnAdyZkl1DC
1uoED9qW5HYrXT2cXxnMiTVHP1l5euQWaJASxYznf+6uZVE3Sx16/tBMRSfW/nSp
ovT5eVZvOYwhqvtmRPkP3kWY7BuLVQsQuoOglcI+SZz2x0nnYZ2PEZcxh6NkxIlv
muwvEjgKniN6ISdWr6oJVbnXO5NQIHLSnFyuzi9aYg2H6IXlyhDde0lXBZejT0c0
nHks+LEGZxlrfb3kao8m9yTWZ4paD75wikvVJEpgeF660m9kGymTmsyDZr1zvMLg
DYHpIiE3WqqqPZ+s8KWayK8YrJxkj4rBxH4SOLbhSWWaPuy6bYSzuJerd57+53KM
EeS89CncRflQs6eI6IEq8db5Mjw5xED0Tu3zJ1o/IFvw2e2tCZEEoexYv40WnH4w
2qeAtpsOSQHHe8ODTepFPtfGyBZ+Mn1ArhaqO6+vaMDrlBBIjBsSc2eFPSknSEy7
mzRbfRGC3iM8uCkoVUQax05gTFoZh41+X6hU7+kDWHAQ9Mkwlb/ST7axitXAbFKu
S9QIizNfdPN6g9a213/gqAhf6d90GZ2yn7H5rb3ScFQpM98OkixeFEQ6QAVzZHJX
Esra8nkrl6s3X0n7ccUpVay70d2qZKh2PkxKRS7LIveyBIwhc/1P5dJhttMBqa+T
Zk8UH5uhu+2Gd6mcS2yXW2b7haSwMbYGDsgpVtlTksazfvKRiL2oVXaxZ5U+iwFK
MfjpI1mwyGAls4mdOBvzoocJVIImsfo2C/lKHUWtOhj0qHii45ZSsIzI9p3Nvlq+
MfT5ncbEYaaihEXQwBEmiqOow5Y+HL74q5tO0Wmkq7SEtPrzrJKjUIxyZS/Ju8RH
UUYWpGjF3sGOt7IOsllZI1IYLqRt2zpL6krUDqnGfZyuL69GgmJNJJ+8XWIsLfu1
X3ApyUaAiD2YTt4dVwgedIFVGvb2GTGCavioHCfRwK0yklRuyIsTLtavvyH26XIF
NNImVrzuChl/XYUte0KW7R2T17Ke5fnd5wVLw/hN0fitgddipTg7r8qT5z0XLVje
29PJ0aIucQMKnracJ/otoEVvcsuL/H0AUAIE5q//H0NWEszAIbGJn2wmp1KOtvZY
RKZyDK/0RQt/2E9q6ZrW7T00UZsKPBNDAtWfx6tBGZqbA/sM3II0znC3CT4IhVsB
gas2xi4VI5Ua9Dd68/bF7hEE15DNMpp9yDA3i1rmqjDuFM4FK1ISTMLDa+wJM9YF
1pUI8TXtF2imv9EyXMgaKluY+kaqN0tjgJtMAt9yeN6Ha13DukXqgDpF9450061X
ZmQDSUmYLpu9F1zhMp1NrZWFP87qk2fpe+5L9OjtmP5tGQjlCjEAGL8WvA7SA2mN
l8gsHcV4r7+chq2dJG7dIqPSkzfEL3ACN7En99a4CBHGQC186JewwWZKQ42ZkhxQ
BTybW1HV9rxRtIptWTC/8/Erh1n+suvfLFzXSlGlRznN6jTjxQy8zjY3PSnWoNdA
Kr2GFdoUfXGlLuywLrt0QvIUyhEHkHVKrhtirSntRjQ7XQIvmH6LuYBeXDD+zrL2
dPVlyaLk5nTHW0DJqOIhbhp3BNsiThxG0kGSXrkpoEavPd85sgnIL8ZF2HALJX2O
bz79LMbGguI7wVEMfqH5WOeMNUryLr1v1f3CWlejwufESsOCsa5baVLqjDw26KHW
jPqP4McJjQiTZ8ajHc4G66WG8Xq1toOzCW2rnwu6PJofKu+UtJL4ZKJRJS7guJ76
beLkIURVFRx5B7LIRjyZxK5z5GT1FwFYq5L59tezPo363alzycX/f/Plr1qCNOxr
HuS7Fm69Ip2beyinndq1S+BBLSwVgBINdFV+paiipEraoPFCsUS2h9vC7CkPlhJ1
M9aEdne9pw47d+yYNJxuedZefnuSJ2KzCdAkjFFSlCcsMJiLAoqK5CFjRM9IQIhr
JXgGuf53BCEN0cD2Vf8YPBbxtb19e4YbirmmwJoN5A2MWp7adSkiWY73g9KWUGZJ
Ir/ZlwqPyNLsSndSKVRuQa/685Qeky1FAJ8C1JR5gNcuJJp5LbpP52qrl0d0VQ3a
PCEk/m4QVcyrnoyktWMZeBdIoSNIjab089f1/9Sdk1Ur0scO4MK4TyNQV8TjJGGy
FcxfPhpSHbLWsV8ASdxYHWIvLX4E1XpOLwX8towWPG72gbpWMRZHLTvOMyK+72M6
K3025jCF9V7XoO78E2M/tX1HbhGbtZ+uLF7p32jrZhbxCGS6M4bKgdTw5PkF8bHt
cexZKF1uuN6uNpt4E/GcM8xcDICK3M4WydvIQ3wuGm8tB0jxgKQ/EUg60oDw0w3k
AxpL1wVdz971IPijoWt/LbbqptkI1f+3Yz/SskhR8t77Z4qHRPJH9gLCkdcrcGo+
FdKmvyM1aXIUU7OrJzpOc1rkUgr5qTmGbYtYDjmURIk2dniQXSPAJtLS++ATLWRn
ggNmvW9ydWqoYLrOEuu1k6zVHldnzZXYR2giKL3d6w5OeO+VMR/Za4yNIONSBGE4
+SHLz56DNm8Xn+9ADkDpnKz0gJ8QGYKDeLmtwqRFUBR+S0oE1ljYeR2GTiqF24wg
VFhhgwArLBcQ8X5Tr3U4cQpNGfTasSZ+FMj4pqSVzlYrXSNkYTDWwFya8AmHEB6e
IWPxD8Y9B1QJeIpA4YB9xu6S+TTVBNsZbz6hkCZtwue5fH6/CRMCk9eIZlbyscUT
EPqs38erCeExyhNFhfV1eAE678dMq8N1Xyj7pkLslsBN20J8D+zvUmdPbyQlzwAG
rMK0IA4emDMhbpSme7GAJgx5OdBB4Jo6fLbjyVy0sICPAhVVhfz22X7jxc0WOFRI
+RBub0p+LFTuQHYFYL6eYYRaoCLnccryBYFe1OIiQP6aDwhKYumGlIE9LCLUFYuQ
vddjHopHur3k8U36ouzoOgWMArinlDCiojSU05+ZHvRo/CshUqgjRTXec9fp+95z
qz5sjOTkr7Mluk2efhIOfncOP0TaKPJwCjD44Cn2B2AfmzYmMmEoPB5UhU16XubI
x+D+qTLN1UYSimlZDrbMr8IUxOjkaT3CydIE9Zw12wi8d2njBNaofyFp49WVraqp
5ooYunSIEI7r1l1l3+M/ink67FEOqXMqPSQvZKNm8kRPDvJvy0R/kgPkHkL0/Dwz
MclXcRR7LgOOBUjUnZx79BaZFYFm46sIzhpCUsGzh9zkYCYBrow/4nB/8fWGQ9cc
RciK2lIGCSQ19OoOagA75cfyQ0TLUxxLLo3ZFAmk/GrEl9m/aLO4LlTU11IZyDsC
G6+CVvi+55ILkgUHwH+l5uTLmE0RXAkiI9zR5PAmlwgn2xn6suK/fbOdlkhlE2gg
O1b1Is22LGXnbanf65WtqjNmietv6MKBAAWJsw3n+FnC3MwwY3pPLauvV1Y/sSf1
74dVYrxpaZUG4gu8IyyRw+8zZF+suy1g+T7sxFhXCqaanhbgFu641so4Q8qXUJIv
sSFnlqBcbegvM8N+2OhK/mCeDpwaT6wHp2Vup5YvAweduuhgPbf3N0hf/WlEV4rv
4sA1n/MDseX3P8kbBefFQ7IemL7yKOPybP+o2xWLe1a5aL2gYh7GLgflGkGZij2j
EVCVR26JhZa9nsYD9WlEenYHOLHNWJFaBb0KvtaXbEgXuCOk9GRgN9WYqxHMFGY1
xQCtKEK8ow+xcY/wYMCXC+bte7b2RKzZyKwcK3/ASKlO4HC03g6+/b/fUva1e5qZ
s0E0DPwNykIYXz7+3S/jDzSG7G5kJNtDEj6ZjxIOiEN0ruSD3M3XqS5JWO2GTCRJ
eDqr8lICtvRV4qeoUgQt3y6h5Chb8f9RxWvkqkUy+k0QdigFndUtG4targ9IxNzF
Ms67xT2C4aaZhcnAlxgLx6u6fTm9HiutxQruS/G7MOz8Pt/DpS5QVsyVAxnb4557
C1tZNPlmsyhjWd/CJPYJhVPzgonMjHQtR4e6j6akLyt3iabTeq+N+BgN5NQhNeHu
cVmRk2LtdgAbi8+QxxMgjbEF74h9d7kNhN7a5RirWC7w5+XWYPNomnKwwzFGWPlH
p1cd4tlaAMpn9srQyT8KqeVZpytYaRHvP5s0L75dAE+jDq/vfHeZoIb7Dc0Vygf9
Ay8SkSFG4eOn2caAgMCMKEHggFY6wS++/VNzMoA3f6bs0rmjQbBMtZK0X7PCCxhl
bgwL+61bLrfUba+7tkpVeXZpX8uAcfiz7GnOT3oKn0XBrmybkBVWwARemfNIbXqk
lDgPk7gWwZa6TEvj329HsbGCkVMCmbqAJsa0tST07WhZe3KRIhvulSefTABxuGws
+VyQyghc6CHLbplyI64P1toEeMZHPlY5LiRiA16Ngid0mQFVq+ylW19DYPMhdav/
UGzRK+RxnNoeauyZ8w929Moknm7F6d0qw1QLXtNTy75uKY0ssfinxVaf4mZdmlE8
fROjJI/rC+gJz2D/4+9dcpb1EzLxB3Xtha/lrTciDlpFjc41fCc5MEd4LeblNklB
uHpDyEE4J7NCOJpAcCm4ijZZTkO7F/tDKljDo258vi1A1tmBht9V+2S4yjt6BGMS
8LvmTcR78GC4zjuNZrIgagpPaIrRjV1FzGa4mANq/Q+a7sCx4tGqi9U2VNwGIlFC
NO+SI8KqdaMbwJEXpuIm+wJTz6UeBJ7tv0y1UDG2S6CPtkaF7hQtC2Gxv87QNAOY
Wn8pNkp7dnAqWSfTgRwuhWoKZA8DWaR6uPdyKQmg/B/hMu2T4oPjkVujIwwGPldt
VcqviCgKgNbxre94jONOJUSh2/N8c+n8993c8Nyp6p7CQbOmrXNUCRgUIly0GhA9
DCJ1s9T8sPfW+goi8WvhP0msIVagM2Fgrw2hhk/SvV1CDaa8QSk2IDpcUOqfev6D
LBx8ZyNtj+9vqjYz+d/2zmEhzeJImbqtdHAnr6/c8vGfEoya3R53g1V7n5ymJ/xo
57knOHgkZihCt+3rJn72YHghU36jVo3HAYQpJtn4nDMuZmCTCb0TAtY1KMfMb/Co
bZMCib4L+pjKi1S9jerlZJLYw5ZAqnTJZcoCpuQ5IKwUgbTwHdUEn4vHWS+g4aC7
SmaosXiTcHKgQLxrE/MtICqTOVv9ooEqD4JIeGmjXzrivLq3nA0fp1tajikFl4dM
c9fy6HWncbIBs8Z9hOxr5fE6WYUj/3jicFHqX+6VoeXlZRmjaWvrGlhp4rOI+3dt
x82OG/5pVy03YrxnTHMChe9EcjSRd0iZbsJhb6f05OpblfBy3U/B4/4Bt323JCSH
MlLThrx4U9CWpNhSA3Lq54Qiq6vymj6YuqKk/v8bqCYjGnEpn47DA+I1z+Vcq3H9
CgaekD8zTvWL7KvmDsf6ng7esLwQQGec55eBsWoGf5XpocYUza3txpe5lV4yhm0n
cdZ3waiMBuS4/F7eSIPiXTYexOU47acMn4l1Eawjtl06o+NeqzQS5YC/MYI9cNdl
1ZMiJOMRTcfKJeSsCQnvy2QLfgqynm6fAZ/MG9hISRwSv3qyOU2HKygWrBcjI5iC
+4St3QFK97WI7i8gixD3Y+/QfidcI1GfxfJ/XEucvIQ/JuChL0govVLwi3nKZdsB
K+S7cnzzxQOMnK9Zgfst9iVaRxvGI6l6uoFmxu2atxJEPOg0iLnyRFGUw+Rojwl5
lzZgLnK8mYeTUcPIjH6QVOq0dScKLONsW2h6tdKXHABGZTDbxL40mH99ABFZzRbP
wcXtKQmWCorYG0uz3e7fDWOci73LSh4Frn8w+raGTDX0LoTCQwvyCWW16NuDfL2s
LPr4FAJd8ZHZIGmIHKRW48j+B0wiEXhTJESq8mCdYkqmnlXeHcjuqh2DwsK0Ii3L
XeDhWgv/FkkUVyhiSewYF3oasiHMwts5/1w5j2iGWPbUDOWQQ2YOfNQwn9NJhG65
rYuYmHQ7KW66w4r29rZdcwUKFNDHOJ80UeBi675KtS0UYOQUM2U+7/gfLCZ/MA/i
k3uy1jIqGoXBnucVyGASdTpycoNTNMu7noL8/FMY/qUPNf5QFhfS7u5xyE2iq162
zGYAsos40zmbnBFtg+yWn6MaSG5mAvOPMru/FzeZH/7438djkRMf3//JdvtQuvIY
syBSeddzbdr0VJR8ODM9pQRTJZ4WT3GjABaziIES1XAZy3iF9qPazqcgKdQXIys0
ihBd2K6DPbVOkDPESS1u3OgQwKnkomkoiG8LuRxfv5GusAF7z41Jc6dw193wDRUM
CbuM3ImRE7LOFIXxHXX0lOV6brewfUAoHbhIHB44zrhL7Fd5VbgRgzcR/YaVuH07
wt0QL8cdX3fKr4J3WpKVKRmV+w3DxKbf37aeZcJVmo9DtxodfSF67L/6fIrDTWHM
sWTxMilms+xnmUv7+vuN7rAExu7UwZQApgEAIRK9ErToFY8MfIklgyt0k6ftnYXH
PZo+BMs9VH8ARZ9wnDe5o0sbIEGI84wRDrqLoU9a5bWqXaTRWpFeENSKJGAdgp4t
nmK/xKeRMYujhCTdl4b269epZsSgscgBMNV06tWBRKX0FOdNVgm7NReBuCUbcSSN
PAfaRZQro4aMGC7MCjoHntMq6C7L3um81tGRxXWSbmLjsTAUvQ1FQtk65km1/Qcw
UVDshmW8mnCKkCg5T23nGg96apQdcALhXB+hXqhliTJuvWgsTPQmwvpSmBwscFZC
3/a6otfLy7+4AdJ9CukePUViPuRdJvWitUpTMGpAD1RJ+TVXq7xB8cO+hXzBRHcf
kMd9RH8r9Kw0Np3RDh+nwGKSuZ7qBu9GCpJurHee38mvQP7Sgggfz3FcdGPQ/Ag7
sUwPwSt/vBsdG6nUOFy7lQbT7obssYCt17GHZBTpXTmMBL6byQLsprdpIeW1jWKT
AAvvjmvsnYROCOeFKpTz20ZWaOMIlyInOFlODZRnyPXPq/BsO4mnD8RTOEzdVB/C
lBO8uQLCZcDsia4K+dGlVV17xOT12ARUlptLIeqDhAf0EAEBdzaUIfNDmR8FVx4d
RImE7lJEfOLxzqS0TP9b2bWgBcU2F5C90CtKqd1rxsxazZomvtOkcemHu7eegm8X
MNs8y/+vJUcp9IV0HFJLbR0tppwB7VHPOeOqU4T6S6T0QrkFmodqvWk1JnFT5ipa
981JnkJWAlgm3+Xgy1CTSykcFXdYm4T/zvpztryThovYX/QEZfvmuhvt2AtUkUi8
PvpEN0zv60Gvqna26hagv+t80ZkbtcbETXwivCFt98lvxOMbCBEt4EfCkMZMrxA5
1UAKoMzG2pUj4fZjn7vDsY8KiaBcLyM7KjE0iKzAcwoEWL0qnl5UBE/cEKhlTCMr
eqbVKW7nzqybkeUsfxB+muXoJ96cQoa3aE7tW9wEodfN8+fNpNbR1tx8KlzslxJr
Pyg/kul5BfJ9OFNsvxlW7qIrznjgTJnAU4zYGDa5ZTn+nCGWs0wIRIg4cBKEOMQr
5JybYC9S4E33B7N+xYq8xlc906EJXIejTlvBuw9viVFaUvLnbTRS7x2I2lZUfLYO
aFNlmQjgiNHesIBqM1gC8nJyHQDWW/MFwydxdMQ17VKqQqM07xuLJC/nMz2BVFh4
Sh9gp5GsSUpIOYMt0bgVLVnsJ9EstjKdrI4HpVG7E6u4vfjawZI5jCKhGefGsKnY
XqTwPUAim5v2mtj1twIalnU2szp1DEQw/oAjVDCTnTWrfwIRBbtoMWp90r0HJCfN
1tt/6p0MsxyeFUe7O5wihSFXlPs3lcJk9H2AhhWoYIojl4rJ5VUUwB2zZWZh0HVY
Kts0AkWwv35mBPqVwEcKHZtOCTd/4/3eOfRvTFHf0SAz/uMvJG8Y2A4z2JR0cDgP
pCJlfsGmEbrNRdnLWWxCTQuiNyDk0dLDjRw8jOCJI/LCPRUWxDsWgc7Ewuona8vs
kmoQ6liBgunUO39HblmwEeMF4GYzseqo2gdbEo1kLM+JhU1XYKoEj0t1OdhWBM5U
A2Zmy8mdmFSxvpoQ2Pbj4Z043cj7z6oOpGm2tzUwW78Jo4Rpwj2liA79/IKT2cdi
2PpqAdgzioxdZ9WSMOVZSTz/b8TEFPlPiwkNbKVZ10on+j2jH7exxlx7k9HToSoB
9k2/puS4BehH+D6US4QcRVKBaSTELPrWdIso+6fEluLV4KLJAjoFIHyap4gwU4+8
nTShvJ5+Tx/h1VHYtyoTMFm5bsgTM3frHRHMfd7JjcvWkHB/VgOnI15zEp9GjjqJ
xjCB01uLli1H/5BzPMQSzpQ4g8DUGekFgYmr8HZCmqWMODSd1oLjWMwl12tnNk0Y
jTd/7LjSk0hT/7wfo83bz9AK/ge3D49ORwi4zLg6V60EchXGprq650kw7J8p1iM7
OqOxMGlkQXZapZl9QOzwEizgO9jAxFYyLIirWekt3I2Elk85qWD2xkmsR366Njvw
7hbnJ81QbIybSLTXcX1rC3zzwj59B4t8BNqM8WeK8h1lvV0k0HnA00IoYyFwkZsL
OKKqwrHb9BM+aRNaZ3ZZKsPmtlJRFdY6YAqs5g41qXtbS8ZgTje+VwUoGttFSppa
SxNgR9/Qkf8Dwkm6xr5pRfDi/pk6Wrl7J4T70JlUZPCHk9ocFsMz/U5bA1lL3mEk
tLcteDdHTrSFtFiZIT61ZdSku/ESNzBTQfWOtBoMPxDk3j/NKa/ANk0hKvto40Xs
WfqyTXwBvvTPpgCTfOkL3N3xlubAHAgFJTwNCmOmdMF6Ygb5ODx48Q9WRTLNYr9X
70Fc7O0AZh1FvG60XgPNntA2hRIJXQaOlqvMgwT2RShp2XjU9P8KrPRr0i6f2V7t
BdcaJXiySCGezQZMTk/RWtU7rHFQfHw1bu3OfgLrg6i/hXDbGU5ccZkBSMEccyoH
zO43btMfm8zipixzj4ISFuMphpd0Jxy4Lee5wYfg6bgFXoQ1t32+N5MPnqbdpphw
vEMehBwuJw/BT6qPrL2sIvNIMm6MNsBzF6Y39BcddlEWSnCqqcBwUHR4dnsVArEI
LQgeBnpla7W237BkvIw87N8I9Cv6AOnGAk6FqLyNhEFSJTdAULB+BVJMQqa6bx+H
FJpaqHSyemrLBsP14wzF/uhkPPJjGi3W6dS5VkWyh7zmEgGIHbLd/snnEQes/aHj
cYSU3kIJ0J5yB3EyKIP2WOhZr4dTFtW9dSW7yspX5tvB08OCBqJ7A6G5PXNwjvBw
JgWKAzv3LL4KedZEQPjgrivdTroQEqHjuGG/DaZOy/hHoyKMUUtVgRlM+3VK+aeY
IO1kt2sjgaRpRzEDVX4eoITB7OE1KL6wiz+y6xPJnQIaI8xMkmrtVS6uKkCj1gpD
D931Lz3EsIdNtdaHycV89XNlROlVA+Huu92yef/Est3dcm3Kd9CCzwyO/cYKSGo+
hdq89dAax79QvJAkMeGuW54/NSKDHAKVxAVSAShG75t7NWv31xRXxlpAfwmAyJk9
d3MgI70iuXp20fBObsNoFXkT/OHP4XsTwgYaufm4n2tJN5sFEkSj6qPXYWnEQCuP
BhUJiXLEwoRQcUVCowWbNcLFBI1AARUTcd0G7mPs+sZ6rkdp6vhhwZshKZF0exvG
G+4brRQpj8sgp64qvuKGW2KPmxy4cbW0X/KcOTjnlI6E7+3SpbpEjB30nejkm72f
mLJOqHkwDQcI+Lt2ahE1D3yq7NEGzYHPpS+EeRudhIHf7gI7mJs5mDQFkHA5Fa6d
WUuqfDQoaagQ5aAnhmtfuQJUGV383U2PsvnClD3UGF1ELFE6KebnNTC94xKz35bN
x3JjtHZ3hgxBBl+5aGSzImCxukVbJNNptRAuwmLcRcv6X6BGFfjY2bmjSVFAEXpc
W7EJWN/TKt7SI/MWXDZljvCCiAZkP6LMoRKlpa9kU3coQ70IZq0lqtNodinhLZAt
eXyRRvLoM9lxibtltPwCS6Sr0tVms+USSYFl+Zj1SIfTPVwEC8nYv3HE2S/gw5WY
wxiv9k7D7Z5UoYV4IfJatpAbHtxKf2HxJttAkMlSyxkPFFtalDwD5CB/ioU76AOX
ZV3Pgm/FHloSt2n7nU2uir1Noncxa7leTy2YNqbPp3uP+a3kmQkhPdyCZAUPJyrX
F9AoX+1PvbEsGFHEZPCI2F6lWvPYiy4ccUzKnDs6FGOjnzv0nE9R4A2AsbqsVulp
WZvO0OCIJQqaZ/fkkUBl8fNEHM0IAGcwnHcFbojQNs9YO9lGnZHbT/9WcGMCX13A
m2xJfiZpTTZYPw0VUWuAq9ItmLNZUMMik58NWoDQkyhDvVzbX5d0rzml4spJ4s/H
QNdm7ZkyB+ruBU33h8zshC4I2jNAjvyndxm/ZSVZt1Hjc12NP0L0/dr/NvZ8O0iz
PrchLentqFAwOxoPGNudpDHOolHcyrhusVgVnsNG7ng0gIaaIhV46pc3UWDXowvj
6In6JatNgyuOCXUjevbUJZgTQqmddd8sG5JQS2aSxCbnk3hP7J+7MQR3wbbPgqpK
hdEkBihOQRVEe+eGd0/BOsb3szB1ZVhShu+OjhFti+6MRjgQgfklm+0Hga+qtqVK
ZXdsA/7ky/PeJ7gtuUd2lus4iBEDmKc1aEvt1x6rY/lU3Ydawf4pknpdleewxEQX
YsxEzSpAHlO2AQgzdH86OiEasPutCMZ91WEq5G2F6UfGv440l8gjj8rVmzD+W6U2
vHEKIzfp405yFnRB7waD4+tT1DvJCKP4PG0gDJ/Zlbsv5Qr9p18pqLosYK6Yf9c5
Q6MsdeFOhRGrX5M7qqHc2OBJK16oZgfBHftrUAHzKAIOEtHrca5/9QjTUbKAiQwR
r/rui4WAU+rUsiQSea+/V8IAO1YcikCdFynYrvCb/JcUi8LEmlHNxyOUsejYns/l
R25/F5UmU7cGmPDrFS2EXHHaHTAhXh/geCtWrygDMk2w2bprfAbvKq+2gLVIUrVY
MK9ofMA55qDUs5XKo18bZipafgu3fc/d/Zb3uQWth8r+2VkZpwd1W/lo0XAp8XdH
h/WBFecX+sVx76H3klTAtF7j2zo+8zJgR2djxHYYD7IVH6CYGe5aRb+j7d5zzZT3
MnOyn6NVn4+qMY0HFw4xq2Xa565JrbqTDlj41emY4qF0DTn60CpeWYOAEZxnO+K0
FA4XM5xtjuT8aGAbUbgR4zn7PBjiDpbEnxHnFE5vW5+/YjOcHtLIs/v9btE/xWkW
U5xM9dviMShdttNgpcQPd7o1MhFEruMvWUfZCmX/IOx07zPEC5g9/tTvl+wNhce9
hA48f+qW4tUZPG9h3QV3G0QsFrWCwfEFDmrKbYmxncCgy9dRUg4Rz/7SN4Epnj6I
2Y1SPPRRdN98JRhBimAg4idmB84xJsj2jHKUxrWNuxWb7uU6VcpQkggwqT4Lx5LP
KnlsL65lswvJ6x5TIJ8Vy9t34LmG4SC1GECOAz2ftiDPSUp97et1OeKZxJbXt8e4
+6wZDxcgm64zgicmkupUg0x9V3UKoBBwnAxAzetWkbrvIVss6pgIiulKMLtI4TWx
Z+u0OmaDt6k2igtufL2KMBurWGQ9bxdYNtTzZoGIBAY7Apuy4goOETfXq6Mc/ks8
iTFaLtsGmoZC8nmyl99ZbBXKuel/WtdlIIlEBTuoro0qsXd60YAkAN4KG9yQM7wl
YMvWj5S/wJGeakuyXF9RL1OnesvRE5C+wj5TJUQaQKPwt92SyPg0HVSg5nFk9fSB
ZxlVZOTnimg/lCKORPtg4tKCbS1+akiogqX3KjjHcj1IhdeRmuZwJK/XJlXbvlj0
UdeYxHr371cGhSglJZgB27J0I1d9+IzlXgdqCz5RHokCoLnp7HZq6QxfhGfuYVLo
k9NepFZcWZPw5qnNsFhQ9VT0jMgwqM5RuyNggz1Ku7eJKoN1DMlXpWTQmAACl3Rg
kgqE9dYDngzUVML8Yx+kTGpIiGot6YeEDF4JR6y77BoCZK2hXtjuvukGvymuoOSB
wEFRJBHdTyOk1YOkjrDIFFx0mQDiJxmCWoZiYYM7wBF5E1TJp4isrIHoAZDkbwZY
ny2LTBIZaecTj3vOBqBS6VeLCHJCQ79GlM2xLmYVw6oBiYCOTHMMoPqkT1eQiEe4
st8cRTzdzSdc7Ceq/LTdSWDRypWDxqOm+169ksJCKMHv71nxbqV1gEroLPDRjL47
YmUOgX8oUkV5aZTcJ3YmE6BdrwwhIRaz+qTT/frHWO4I/0/11JRlXXu1RGxhHMI7
7757lB6w5qVnhmA/rvQStlloC0ZB36F3KC2vLrquzZ4/XgkZw11LUL/ScZMHQUBZ
m0U3WmTCLfuxotPVvhdmlKyKfosopa+O9vtuvA8qW5K0eLdVT3+OIFSOiSbhUsP6
ME1V6sBsOACLHIYnYaaQW+U1YY6zFss4v+mR/iecfRMuTzD29nBEa5HI9H704Zay
nKVY1jCdbO1agqEoTMVbcsaTInkja5QRjGZ4mYaSoDvioS66LQ3nh3N1T6ohYTP/
dJEkBgHC7Riy2uWHL5PqPh7pqFvQfm2sKZZP9iNWZfWnkzFmyOVbF6lVn4d928qu
RSTxwidzNtntsQiQ7Q9y77QJB2nUPNWMYSNP+zj8vryd3Hn9u/IVcCW2yd9KgiOM
jZDex9MJ4349KhKT+w9sb+27T4Y1FSa19ZXlSLPPwolBsvxFr+RVIq2oTlHFRg1Y
byyHhxOIPjtQsjQlSa8KmsIvXo6mcweCKkkUl7mik6h+UWKdolAmeUOWgrmmSgmx
u4PEt4ehfb0TVNsmPdkV2MUZCqZfeOp7/euO3+PhQK2eZYV2xiXopjP6Sdog84zE
w6ot8hfW+9myb3Bdl9zflm1kClii38XiUurX75wCAigiYzFFmWf1Hl1VXNqYINeP
0CQE1ew63vMUqtDs2cYsD9YTmc+w3Wu8YCifIp/byPCKy9P15I8ZjRoIpfnTP2X9
DHCcUn23ACLrERtju2MSSBDuFWDqQcIRcioZLgLYHDU9qh+JoaMJ24yqjt5JPmIZ
196GNzfXR4wGkkpzO0JVIG9wL9P4rL1Dm8Gnt+murzo1eqwmEq4xzPEsCedDw4o0
fSLP7UgF+lRfdq9ULaswU1smM1HsngUBln7WiXSqSoyB6i1H6jVjRpjy/eKehRG9
yKmBKL4cB5u6tNRd4fp5yXIt5deGB7O+5LrZzny5ULmJqeKZ+BeZiORMfvwJsrpX
Rnd8SGeE6kBt28gPZIbccnblUiEUZK1sACpH2g6yrZxi98FHljV60K/kMhxP0oKN
mDflrc2DkGmkZVUyzdQochN1ZFyKtvdHqudO/v9vAwwgqBrR4lTVIHcwYEhPW71J
t646BMLSUlxpdlwxnw8BKL43xDNO1aCdT4wEZvYx4iegIWwMH/Sn1jTHVdW+swm7
uBllr5QapOzjzrFpwsKeURsJYzOCHtRoKjTj4x+B+a4oh6lUH+MEVtunV7dqOfSG
qpKUuannVsin58J6iIdy81ebvnXcoznLakroEeW7ftYrnogXSqO9pYrxbowKsRYc
ZXK/qnhX50qIaeZpdTkvXJQox1ED4BITR6+oHJgWAAOZFWq4dQ3fMvuZSugiht+d
dfBpPzCvcEgg6GwG+GOu0R7BDsZIsAnXHPVSBtX3h/vKiG5QQyXQ9KsjAknC0wfP
1CRt8nViLcz8psfG9ta7ADmcy+182WwwCqzKoGVuEPGbtiNLhBZnflJhKCSqOmEE
ZfrUz0kd6zt2Az7Npi81ujORHJwcyDeHZdaDHL2pppb9N7FCmDR1d+KR3/UdS/T7
u1z8woK1LCtyp+CCC8RFdRcu7TR8zdJ4/nUvVlL7GM3Xwqx3usNwVkaoFMwHwu2m
C3ummkNv68IkkRl+KWBthqCZ6BX7lyAp0y3a3VIVxdMZasRXaovsKjrs6YZv8zhg
YY2caQrP7uqpyHtGckzWJAcPuXg8lGo2ucf5CBI4NIQl0mxvTrxQUSsVCsVhqajd
z1HifTO0vYxh15qxtSL7Ieq2S5zZ7JBvvSRAxi7LYwWTqpq0cL06MDPeuVElSOad
xsO7AldYMLJdJ/8oak/8SOQ3aQ45LaMXdXafcz3p7NxChXpwFR3rxNCCWSrmYHhB
xFxKkgrrY/39kikCS3vC9HhBF6aeaRitVVbmhVzRkY6BUyDlIb9eAAiVlcYN7WGc
N+EinJ7sYMVyoqmePKmzD4OVZz7qZ6Dekpn8i0vXRcSdluPiRdXXbjo4SIQw4Pf7
sBRTuFFKOmYpadYy+APsu3+4/u3JagnLgo2Kj9CItYUjbwEIIiKtbg2i6mklViWU
bzgvHMgxA7PlHM+H33J0OUNJxfpM4BNntitFqVLDro95ThdNS0fv7uv0jB6fbcE8
xJ4CLGOdOCg3SbjMIpXfQ2v9vo7ImP3lyNVBLSRbSycZREfc+aGPysXpHhzXKZ7I
dtASEVpdizUQy+VRd4KGyIUr3iKQ2lm0+HuRUCskwe7vesmjEytsZ8QAPbA3TKGo
17Z+sarTT0zYW6hA4gKiv+tdVC0uqRMnGquhPlJa/KiM9h/jL5JIrWdlkh4ha7TF
8cWd9vuze3LupnWNkRhY9c77TpkDgSaRMytMYVuALPXrM0yWpWY5e0t8IH9nxTRD
eokYqudBqUD/HthmzKpa62mkLVTOAWzdCYYr0eC1brYPEuLnlPWRurQOMvf3SNdh
6+44IRAmx3Yfy4FASWkgRSoGG/1RrW/gnHAGkmM69+Gi2Z6gxpI7LcyoqsYEtDaL
q5gi7SVl12TV6qYs5svgRw4s2uBe+SUBB9YT6J7EJeTcLw1cZChvJnjg1irCfKws
aNYzgbt/LQxoYMol8Hak9TmitcqiDGUp4GENBD4LN0T8PO2nJm9CtibpfGH73j9X
v3WM1FTVbiRonmtG08ZKDzanv2CWCNCcD4VTb7cQCr2P7JVL+rA/ryNgk3zGuO9m
QH4g87fa9l/Pa/Byr2dMih5DpGihUFs616Mebnd3xUtVix0grvKgLla1Yl0yOL6w
ZmlB2SXBFUC/d33crmO0d0q6V4wu87LouJCmN0VnVNC4wOIzLIaTh/O9MZuPP+EH
7K+dLPOnKCRf3/lP5N7drpzYKOAHxUkCGp2evX/zo57kAINc8SjejG75rz63tUxK
g9tVwNkRyWe8RqJiTTyA2teH5bYH9WD75JIf7Ro+iHwGMXMdWpmyNG86cY4PAKpd
rlWi+r1btohcaDODIMDEJ22kq4EPv+sAWmLJUSGtqB4Prtvnlos/zk/l0qbSdBQA
s45TLScCv6spIVAS6fF76bCr1zqjFH5/ohf0ncvN5SQSGUeXMuKwcG8eLSRDNvcM
49HiKWgLU0SFiM/odU0DNv9xgsSEj9/+iHATTJ+xtJwzyHbPJt2ip4QfHVuGyCeH
Gi9kqJuVOhjmeffBpNQwbgbEBkOFbuy3mNLpm8Ug2KIIgJhAnzXMQXaRIa3OgeMr
icE3ktb5CGNkUk5hSbDlf3v43Xga9MbSMDEx3HFYwe/ykz0tgw7S+a+EtG39Lgp3
awkCxIEM8G19uIqUQJGq/FK4Ab7dJSXc5doj0esjvQhZdQKjETumQsnCkbu4qG+5
X3wG7gdfXmcuhWXNMDKGo3iTQbksndq1sih46C8UH/9RJMUeXsK+JzgzE2Vml7//
PorcTdoyaQYXEW3TGeqQsSdgX7oZc6UOEtu0fwb3MNal1dhFLBHxGPlaoxVOLJWL
mpGq7WeO84uginaR22FSqTlgy02iufpL+LVIjE94B1rFL0Duh9OibqyWNe1j+8gR
BsdZUtrPGqubnpPD5dpG54R2cym/htGa4XgqV0RJF/ljF8e2UgA7N+mt2KaQZHRq
o0kDI1zeg25jKce7g1lFdpkaBTzFwGU3QEBy5yEzeaEkuWhc2LC42rZ2zpszleB9
GzK4mop1bPlzHx8zO24k9YKj9lpVRh4nRYc990VejFBbVz0KVxZpGV/8EYTjCBYZ
w3ArS+iV8FUChy5KHwnZ+kZv1OYpZAdON0Rjtpt8em1mnQOmhnWBsvMweiufJhKC
p3NHrgLybaZXJGi+Yh436EQw7Pvf0pwZSBVcJVlI932V2542Qm8OR0kB3HECaF/z
Zv7hGOBK1fY875iQqZFlTNy31C6ZJarzFwj/VQf1Yy080KKCdIpp7888I8D2KfpO
RtMivIMm+zjMhdck9hj/WQtTVh+1bbPUnvip7bwrq/Buyx2WNP54wEQ4Q2Ar3QY4
NQKCCYxZ4sG31Eojr6KeOHpDPIO2+BDjzhh7T8MUTg6tPI1DE0ZJHSU7xnLGpWWA
LC4EhCs66qqujOGaj/W8Pf8HFZT4XrUO6XvwTlczAM9QzpCOKZZ5PDI9viHhlvvI
8q+Yn0FDiHOqFg+ZlKpSqya0NuTv+O7a/gIr470K55Bf4zp3iXb/6FDYY7Eozr+i
F4Yfc1U0Y4gbSgxQCHM2KolS+EpKt1ljvLmAZzoMzaSUXRfVV0MEMG1kSztIhoNi
imb/y/M4J4IydLpNraE3hlLVX4vQJU0t59yC/Ds1TCo5UU+NV5C5lcWGE8T5MqpM
ziFPJS5XZGWbupLAMVY6gkWz4ezpn/Rba1t3YvXOZeNC8e6M/fl8MByWY2fMkgFa
GCNnq+yUtfSTwD5DsFZEjREDM4ICnB057nI93l8UFJTdx97BbYHn83KH2pxPN9q/
CslftLVreva32+AdDrqQprjDNpMn3SG+Xcnx9/jWfjn/q4QUyMLFYj+3teMvpi7C
JA5xrIUIZFBG/lPjDsZmtRdU/nUcjvnNRbuJJtgxeRljuHcw3gw9lIfB0DPt+oQH
uJSLae37/rvEkFMRCavg/GED0lCS2Ccj6WAzo0Txv66ZooYRQ/tY85gr4MF9tsjT
euMWKw7wDSDKvwsb77k2fwLk4GhSOZQVTESwdMb/4SF5enYstRDvoiNGg7R2ISrX
4DafkXCp8rI5UM8Mvsbi8ehaqIwyGzq/3aXCLLKEPYO35KEsuZtJEd/UO3JxaMHH
T0FUE49H2cQiFfPFNgAroOp6gNrzQiW+NKrKjDqcMgQhNwk045rsCGk/3cwukL6F
A4afSVhMSTtuwqWNDN+nBteMO78Y8wehxZApdridYGKyN/7COshDlgw3XC+KQN9f
7MjC4X8TkPcjVd7h58HyZ6yodCnGhxboSk3/xN5C0sJQ+5nLVe8xI23SLZW9p3wM
YoMj5t520ubKhkbzc3rs3d8wV1jaa9QigZOD8RX3MXvDCAasnHV/BjVQj+4XLLtV
Msy5CHYRDImXBu6BfeHRYJoflruHLtUGgyhr0SABzRu0T3kyJ3ChrqzSHTzpfIGY
XEvM9JK9jWgy2KXQGb0iYpvKApf2S1kCmqXDZhzXBqt/eWIJkT873dgUr9g6mTGv
1mefMwGEPPBZST/7WZ5LiGFe8RJaRG9jHPE+EIpLIIQglwdwCUYAw4tujlb9Utsn
SdLdnGD8C7JAVv/IEMbFG6tlHeTV92yBQm55s9xboOu3RCe1+RRtn7JV2K5k7pRd
EIK1LfxLuCRXo8sKq8PkxDlmlD7lhy4cA+DjZskOO3IlC3P3JfRMNGYw/FWc829/
QFswjynS0ILQfKzLxGPTYImEQkN18EMjYL57c7LgD+L2SgsPxRrQ/RhGFs2k3wZx
32p6x4SMw0HVluT7anrAIBwea8wyBSyw+5C+jaJJGkb6XUStWoImNC9r3/o6nMaN
BvKNM3tOo97CMiWFo5n6p5ivHSaHlgS0mxTBJ/pzhhKyfi0NdkW5s3c8ZPzlIrKi
5PjxaCK7Tkk6FDRDL0NY5IH/jNCcJNInXVA6aeUJpI0PhfB0v9ybVkqZD22cY7x6
Do5jn8E51pwRqWRIe33O+sI4KCPR1EogujyYh/ZP4pnJ4vE4fEL+/5eJAQP3zDfv
dmyM+wdk0PkKk4oKJ7Gyq2suA1MnpMxoYWo5o3geBP6fInK1mIv9cjO05IeDcVJ1
WU1bBnqfUHPxDHW16k3kMHByS4q82oUcqc+/R+prD8VhJR+o+3VSlgrYaORBGpmD
V2saUhrgvvYNcd2ZuWp/YCpdqaYcKQbUQg4foEl4JskhZUgOv9pJcj9OcYE0soLs
rJARcA4PS4vyi3sN+4aVqnf06Sa9zFfbjXgqbuJYndZyB1aSul4cQl9wMmFQL2Jf
hLvZpgvMfp5Ssx7pL4lQrfKBPKjggxo8Vgo41/wtAAmJt6k/CXjXXL1+G09D7rV7
sQFhVLPq95/COEv0PvHkTJ7FtJZAZUEprsxkuQJZIxe4t0L+3ZF8T8afFWJXP+nE
bG3pwPS1DI1H2hjI8a1fuuVV/6v3TQT4Wr3exWldaFQlt3JKQRqFsIsyj3XzFg39
5nOPAzSxZA4yLeBPexZhQTmiscddv4oXtF+kE9agbiLQynR+GeaA+kghYE17PaPa
imM3gys6U2PNMzaV4zOb2xWzJhODcAf/H/ZAJoz/EnsCKFgE20iYGD1vcDOBEg8f
CIRJZtxLkSt5g2weAl3jeziLpKpaaN6d20X5STprP7ITlnP8mcQ/wYyOF1LHyisf
jWjUV1MmuHGE99gMLnNZWjpPpy+g3dZCoNkypdWZMrKDOu7sCAn2P7WSdKf1RZMU
QJrHo5eBzat+U+B92IjvYJKyEzt5xIvdCNaszkMFmxdUs/IuiN6S82d9E8cJjMMa
cts60rjOYsSDh1dxEtSJ1Asj/59xuN+o7iMsPwyp5tNLZgG6o8dzKjpj5y6eIYPX
bmU9tw+VLRO4WoyTOHLbjeHBwV22eetydQzUvbJSDxoeIDpZI32X3sBKH/ywFLEu
Yqtyw7GFBG9haqg9hBg/rUZq2n3IR2kwIE3yre1oKbt0mLfBVrz+vG9vV+JcOexG
VhZEy3KbQgmFLsM+RaXZ9+92HAPLwEZJj0aDz/Ex3Q+sHp/ChPn20QA6oJ7DtJ5N
Vuw1oQsfz+L+ayMwby6wmRAkkfNJz8cUZAVG8KBbveMWqfODy6++Gfa5B9b1kxON
V2RtbTOm/ww5kQmh5gnOV3CLNqTykF1TDEW6HheV3GYG0iRHifJ1D/aW4VGRaw7s
WyGdfGERj15tYhRV7tAHUKSjY63gNIFra9BSSz5KNrOVtI6g+iLxJRkppATLXBKT
/G+60t1lNq2ZihOGVCfwjuaBidWTTQeKD4lFuGerrp0J73WTIM71uhP2a5NLpbNT
6RXvoLW0wJz9roS30VbdvuFqyy/N5S8uZ8MONlr6SquRzcEt2wS9XALWx6SEZCLH
rOrK25fx6m15vYxL9Rz9vWQB7CYOd4TyTxY8apDOrz1X+Lwy81u9yUAtCCrqOMjC
FGfvS9ORJ4IBUAAz3DOvDzb8PZZ/IIlfDJPxZdsCUB4mwTjIMHpL4YFELKXoIwiC
yOfO1a+ypu6FiDaFvgXfQPbR0d04vp+YfoeTCve7mEHlV4hTRTPStQm0XmSOaFqE
7wltamrXEkoqSErJ0voNEhwFw3Y8wPyOc430iAZQR1JtYOlu4/c+yDcrLtF87WEc
6UEbqB0rxVLwLnqeIrLpLEJwIr71WqijbU23PFCMj0fnwdKWPTOubMT/HrM3ZGTP
eagzDNec8Yy6YlCL7JCfpocqMjroX51/88Ih2/w8Kpb+6dbVRJaakywy91tQwsub
VyLm0CWPIjfYIxsna5cmxV8AEvZ8siuuw70QtxmiJ5FbujHPLrnTNYsHFlriy+8Z
g6fn6gb9t1xnO6y9kJM8YnGUk0hjZ1afRVLkZWbahFcQmLJefGO6ogBokTVxbwV7
uKiTugRYTuuwHoQ6YUuZRM9eUJGDd3rwrMhuj4nUJBsGKN6VOgRfQsyoKWLz1uB/
S3p2jSuQ9zWFeXsoomqOy3kGMVq4JyuwbH+FRVQbSSDHm1u+gIBsGmjJ5b+cCzop
Hrvcj7hAvb/DRBY8sVfYW1hYYkqtvWcgF+UW8/IQQo310vf/koIjHn9CANeSdwAE
St9A2t7sJOVA8eQWeF6vYlD+DesiXlyh4EUzM7coSMAeoFZRPGFg1p90xFBQUank
uDlUS5L0FW0nOc6cWhx3hlx1mhE15FQiuxhPIicfxgN4tzT+49NJg5OOXBqj/zH9
EnsOBOgBETLdCcaYvl9uAtwq7hy2pm/pi8DplxUNw4MBCEm9kNiEQlYArFL5veAr
L+f/G/eBG2zDs+M1sSPCGE6A2X2sn2KxNtwK/eAprqT+BETDGQX6H376+9Ug4GF9
XLGnY2XquA7wdkHS1E1/0OHKRiK6Jg0//5sK03BYL+lknFGwvJmZk6jTUVEYbyYz
hukMDzKX7IOdUGV5Ky7Mi/fMe+V5Lyj/zs+1jK5rffaBVkwFbnckQHGPOqzFAb1v
nkOtMMiYYoNznua69K65I+NpGiA62PvxompAffWdQdCKuMzhF6wtC6kr9oJWfl7t
8XnTbQXfgrXVE7D4jPSn+Gi0X0rtLHQPmDNoX5trIPpFnlw0HwjQzYPrLhjgaFpt
vKPHQu6pNTFzkCnw8YUn7lRSOP6g/taK9c8HppcUqcuDJtsQ228c2PVnI9Trx6DC
OvoQOR2MZYcQdDA3Tq4DJvNwzewTZy94RIE67VJcNVbdIlUy7Wt5YABPE48EdWpj
y6vEP7UAbM5zRJS60Rsz0+wKNMf59xvBWoFjC+U5tELh7du4COUes+L/u6ZTP/1a
6Mog5jsQ73yfbrI5e1vjVkexqssFBwH4CY1bjSvaOdKlxMgeleTvsCTtswwSArzI
OMO6jNLayfKcgp4/CpgJLJXTQBxizHFBafvL+tAc/v83/boP7Nk/4xUe8F/0ZYlT
W9+YOkHbVV6/4H6KSiIBL4m95uAzNCm8yV6bFf/VBt2XswimzkDKyetoXdezYitL
tmW/7p3NYujySuEAnilODnjsZzR5hyJnwGjqnyBEvXmQh4H4JFwH+KBvoZbg3vWx
tmWu6uHFo7pLqgWPZoJR/bsE9L3AwmMlVPjuHTr0740EhxVhnzqUzG+7qU7vQJnJ
1JD7BQlDChm/PdESJlXsKx5ApyEnGovwsWfzYvGh7vRER2oCr0PvnuY2LyGGs00M
TsYFYhMDqDtKC9Mcp7UwwMnXEGittj/hCoORFZFQDlSWboUnpMH1oxoau0X28es9
4VT0gcTy00Hc7DrsfFikDfRgjd1eXa2VxnquVkddoFuqEfGCcqDsUgALc4BUGq6r
Lmcwb9G8nNiDCFrzZf1tElJ6SEbR4JuXRaAsuM7gEwMMMRhX/67OCHM7T/5OnDJJ
twdPMDZcSfMcECJfuMLuF+bnyWF6IQbEJ3lUtDDvE5Cv+1FfLl+L3v/mAO3MV2bM
ayV9WTssiDq9OI651mNKfp5GRNj98fgRiGX4Yus9aI/QXsSsH6Gtm8WW0s9H/eM9
A7UKS+caZwgxWI2WyVSiBUnx4REvqvrNuHlxHukqtZNxQwBXT8g+nMS+QmhLS/o9
vKRRxZ1ITSjc0xtmrz49CHfKRFuPmwgI46jsUKhgRkz2jiR8oyQLBaAlvMO9ZxRp
74Q7YOXZKUYSurwDKnPx4TcwMRhWPMXj3QmFhtGVEXfUHyXQxjN7544nm/8BvZKV
RVGwwzHba3heBrC8tgTYweqO2HB/Vso1rLFG55x3zD6ThxhL/0+XakRKSpFFgOwQ
wVdKf5TbeE5m4epU/PDCEn4qX88xqtYTvfDg/n+NU7fqO3l65wREyvZRt6JZKcwg
Y6dCnSNwLg/RYr4FXTCII6eNP1MBjud+vnzHzz03UmGcZKTEvEw96IsBMHbES1/t
aTZfcZeKt1WmR1hhztMrA8HAd8eIK9XYb/LxZ9hVAXa+eJPWxAshvy5MbmxJQa72
48XsxFBI+Li8HG9WWzctqBAv+LOvGXJ2BvZpGbG0AyLir2EJS4TkAwYflrf6ny0I
pfmm7QTqxYq4AacxmAvibD5PkVTYDO7Mycf7PoiWopF057k77zdl8mZiy7Vfb+Tv
yh4QZ+ACiheZNKKbMwb67MiXkXSOj7Hg1TFZfyTi9OcLOf0oH3M1hjoQQqtuetI/
bVVX9nEZRyJ/EH1QBFBB3X8liyDcy+VTDHI/EdB32Jr00Zg7hclZH7ezG8OpyjS2
TrESKVTqTEUb6JVWZwUZe34jwQwVph3sglFf2YZ7/svy30FFNPOi6LU9rFUsSO7C
pGk/aXcxlvhC0lxlDrSHR97U5lj2Us+K5cM4pxX88RlmNxI74i3b4h1GQu6CaTgG
yLnctW6wKy0KZ97XxyazP4/2LDpt75ROO8hUpGlPPghFGTaMMRDd0oQy9osY8uo0
KIAtulTc2s1jDnk0u6W6UCp5B6sXD3kYUowJ0WfpMtFYrMozHYz68jxt/E6JiSV1
skpLMAaZgt6wublU7eMSd35aH6wHMtXEv03v65yN3VA+2HW9FsgJQnZ1CPp1q1aK
UbxXZztD/BBKVluzLhwd0ZZ3n2yk63J9BpNYQuUalClUV6eIjUXNmCcY9xf+h55r
/MZPuj+pDHMWWuE1y5sdydOeMear9IyWJevprFQcupj1kKkkqom35nRlDuco2fP9
qWCGn2oE2D1W8oNlxy1fH08eF8wAWFLDyZSZ1uChjqBShJBIgcFNxzzzI202AGgF
LzIwfcl5J1kvS9JY7cTQ089JgQWstO2qpnyWu4xvqsjoby1qIun6TpjR3q7M7Acu
3pSoNVn7JpNBcdtpwC5iAUSYAyrHchO9gQ36iE06/9G3PT5VFig4BosnkquyBXyI
BKLhr/w8OH3F5Hb/HHSb3Z0PNPbPCgoZyPOzky31XUGChyfmugiJYIL5rvvsrz1q
awaebpEF0wr7ecDOixK3vfPAZ6lGy6izay8wzuEa9OX9TK0zzSMcsXrQgRewExEB
tcUaZP3y3A1d+b0Ob+XteQSHrL0KGRI0/DQ+SR7lFkvI/rhvALYxUg9SCuOl0xIS
zq5Gj/2iHfsqGqvX0X9O+EtkX5UnmoyWyM6bU5E67e5l1vlUFiU3s0ILkS/a4B6o
lRCzxbD+9DsvtWb/6cVrRCfWhVTdrckY+HBotYiOeFrVwVkTgD/5a0f2C/jjSrrI
XORbXh+AP5DS2tho/zsvWcUV5/8ND4lyNxED1jt2RR0+BbbkaiSQD04+YtdpubbB
c8ALIMATwCxTBIcbkxzH9ayO4nsbN6yK5uLPcdqzJSazb+1yYoWfym/Jl8GanyXb
g+0BZF6DN4usAwyUe4gmEUtbuwXPtCXvtc1ooxfP4WzIbP4/kOSlYXbI85QneOdw
/ocrgtneCldWMN67yiqo5xdT5dQ5Oej/tMCcH/84+V1msS6Kt85zxJkpKJqVohXA
Kaia9uUpMwEpiRe9jnk25/9RRmePmxPsN4auHdMoaJupclrznclje+riDbjyxsmf
uO38/ROaAYbouJq3ek8Gfwi2lLJyeURrjLnbp6vy/KdZKOWzSAZTRqb4Y9qDzhP7
zUwJRGRQLer9fyjCVHcOt3Kg4r7P0MlwOhyMrAuQmMwf8hIaN+7b+eXi+9RTzXr6
P+M9eS6NyqIDJEyalEM5DuIw7i4FEtABbk8+GZ3Lgw50Uti3y32kYa6KGXkaPshU
XYwv2dMp+AQi8vixc1ELczEHcflN1FpnngLxSyYxhTYvlGFfeucSGDl2T7t8eesg
oFKFl2YeMAO+7KkXk0ZM9C7AglLffZOkUaIzDyaJXVcatVZ39JCLWrmSE3o5j2oE
KN4PiXlOKeMj4G71LMD8kDc6xrAKOeRu8erFpSslert72dr+aooDrMwh1M0p5XsZ
PutmuiRTQdOYeeCXPnWT9lnedbvA/qj8B8T3vi0VCGpTxg8K1qLKYXPWLTXJ/hc/
SJ4ASxVO8r/iBeccx4lRkp97Mn6rIkHrqfbL8nsbiDtMMyTgg+kOMO45A+lM6Y4p
mjQMUNdI9hkyvI/vqRGBqbLtMneiyF9lco5Oh/WtEiAGqnSCNXrTcHY7X9m5/KVC
fh6ZQa2xA2M6QXNOOBIJExlvlcmU/tZiz7uadScAEUk6r6NKDGZ8Ht67KNgDG/tz
vM90bhdB3uMH0+wIIdSZmurNz6hS7K6a+5bXMAsbQBF/ekh+z6p6tTHgL1y3WExf
/Cz4SF7SixzZY1OdwEKe7jWgkKXumrWrrcnXUB4qA9QdMTaerDaacBmNAdr3WBJg
sQVed1ewOyFloZhU6TL0tPBgZnE0ond2qje6HbrcFsYxE0oYtBQjzdV5dGfeVpGV
K7+DiLyg8hZReYLpkN7pKna5uoU6VNAPKk4E6//OAp+/9nuJaXsXd2O+QcifhR5z
/AFr79U4p94Aj1d+QUj6yBNKZR2wFhMoKEzREcqJxyXo6wFi0Ar0wwFMimYh1hBb
oOXzoYlDVd+xKsRCEOmneKqjPT8r4i2lYsjn+Joha6/dih2DF+4M1ecKNNhePHhO
vlTpIm3kUAXDwcbjUOZxkvmTTFMRX6+xoh8jtCaq2sID6UfgGw8VPbL08lleSK6s
ymiP3Yq/hfJhIiXvdTp5Fy5QIJIBU30sIddMDK3aRIEoopm9Neb5a5apM5ooUWy1
ZZnAj6BZKa2YeUcumpln/DjalHnvzAhUHA/JYAtQ309/S0704pTlJ2CZms80/w6+
rbL0t6JYBjzEDZi2GMWH4bW6KELYpeuueKXR+vxv3G8Sq5o5ZUI3vlUNQATTyZrG
xdy3tjw/oiqK+RfnBPKU/5WiRpalwM/rZr6oDMjfx0s3MLpdBe9FAcHlcVvSI/5S
Ta/fSxUr8zM3UyKU2rX0zPTUG8EkdseAw/AAaiL1U4m67VmSo2UkOCsxRSFpIozK
OQg26CgjmoIIBfna4Y8PdSvbncrTahKtbYFO9UQmQy4UPV6e+ZrxOr6B2k2xiZBo
VrnOmlj2Z4jIBPY8c1PUgJ4UQUaOpAzFaghN+RfKDjNfWXjXznzz5Bn/zj7p9eaU
17RY/MaK+D/ZuZBERJ5aD1Y3FnrcugcxTp91lsRVRQQ7c3Mu/et2MClIx9TDXAGh
6325iOVHT43ATIrgCOP58lvp/iDPx8aQrhz4gjTrXm193ps4JNY/Xo3LAVpU0FL+
310vOUAVvGI0seWl8VE59l+RBHcJuJ62a6u6xg4caAdwivxhFvMdD9hHURkmD/Dl
bjkIVWN+P9+vm5NQWgJCRShyJEqydT/09BLafKS6+Ki+9w/PauhVJjf2F6pB16QH
Oi7t3+WJ4um0SKtTSveikjG8UoXKv+tlNJgXVah5ZGd1woZBTTH2OlDgWQYja3rr
0dU6twK/vmSZ273kjtWQ0znSNirsEkwH85LoAGJA38dwqmIjUw+x3IQJMffyQQH/
l/rhDZZfhYe9sf4QvHmUekLE8bLq+FBOPf+xxpDFOiGkGeW/OpXrPOydkv53QQv2
7n5oHxV4L6v201EV0podMDXJ0ws35kR+/zi5S6sQ2YnQDQWCMpg/1h8BXyAdgZN2
tVUcey/NaYNl8e+X0ynyWxz8fV17NjBdIPEleOWpQfXQGO+dJYF4e8w5QNzGjlEQ
G1ZHY28J+f/8qmqYM0YIwUmjlDhZtbE1kjSux25lAzLOYAdQvI2mPq5QU3rwhMmQ
nDOTjT1eSvjSdPTnTL0FX0Yam3vVAiM2dOpHGFlsT4H9B4MJjpSkiapl4d6kwTlO
L5rYrtmFg7oNK71yzKHn0fw5rzyuqslETSqp+RRDLY8JARc/DX1gWuv2ojqsN8wN
mEK73BkGxzbywqnvYiTq9Hxr4O3XYQ3pMVGlQ76N7xq8Deeja/OzHCqsmn4GOzB1
wbGfH7AK7AVTd842NlklKzlV9REShz2yahUPbpyv11xkP9esUXLpH/KtLBzOv+Jc
iF8z7Dq8A3bh+cUzir2ttM1NU8UmO7w15RnPQBe82wmy5OqewMBem0PM27dGnziZ
E4Wwg1josRIBydio+l2R8O0lACxVuk1x3ILwYH8D67jOdM2/wOqMa9ezWMXW6U5V
kggsARn/I1LE19lRHO1XLgIz8yFnGSBfKpKmhNcF4uMi2qwyVl68/gPGNnTeg3oc
Rqg0aETwtRmH80nwA8FFXEnqee/Pzac5k+bDs1eHc398LbM+tAKi6D3WM3gjL78U
ReZx4mFxYjUXU27SvXKQi55F74PODTE7hg3xqxkZlbbysW9dHN06EUuVi/+c/bEJ
LSSw4ZgjigXNLT0W6CuttNaaj/++KVWtG56Kngve14/Q/jTjr+rR3tTBWWWtUItL
0eUlXOeUgmTGjflD61A0/geharu2BOgG0Ss09hBUSuTjq1K2js1yxQzR9habgMoB
M8FCLzou1vkd+z7LgWtxovvnfbTfL61EL31hSGkleVDcH2nx3UQOE/PulmYBHzr6
le8if2/toMMzdPorha27hBMb5Fb3wxBhErJQDfjD/zJoOaUxkXe2ZtOgcffq332T
sFvRfX9hrh1LzfphV3DTs0aCXmBZJWBiJMO6lXeZiR5i+uNh0mGaafWueSaeCRZE
tAf73DS+/rCrGNhSpCzxzAyXq/oQBXh9/zMTqt32sgQxijAHGdgO9phVTi+EdkW4
eyZXAJ+qtUq1l0ZEvkRfeXmAArC6WY25jXsFQWEsjGHOwOHtfaVog2UyiKq3hLAQ
/gZ0H9XvGYvSAeK+nLb3gE/EYtdhIKO1OvbTjgpCAU/V0pgf60reZLP+S74dV07J
EXxj2cFkaZJGUVaw4/EfzrME0Q5ezN1nreZJ9CByOFCz80RVytZdbKqt1+gAIOYr
hsBkVV6htf0kENX8yHPRRBNT3P34yID7ra7blmI0UghGPB+zJr9eEOKU7lapZbNx
m4pgPtaQYeUy8pzyu217O8whXMteadoZkUCGKULJdBirC2mjW328L7JxEyM1OzRv
Xgt1YxeO5QU//QQhQ8+BZ/Jbhm3KbPYq18dp8h+G/1bP+ryiJRi1Ndf4spwdELsk
v0u8+wFeVZJgUgi+2sb0/bvnHzztmqJ+gJuCdQVkAqJr90makp5duMLvJjEtr4kF
toGCaPJ26glO2uJXDen8kVXVgMca75cHMn2Xwe3TuzFppakMBv5xY8yqKkOvC/JO
usWTO7cErXZY0XD6MzL/mO4dX1h/XUM1gnCHAsePcXuzWLsbIJEYmK7aRkjGZvLl
eYLtlqRZvybdjkmAKIL9uKOq/W4JeWju88kizCnTQEJ1sfLSLXl1Ybk6Ig+Ym7VI
HgRbrDauZwHDaMru59SfFjk+jtrDw8TBMOjQ3Lz/fJredDSN2qPb1QsJGM6LL2HH
5VRZmDzhYIAgnbR8J/hqmh9sCfu1rvm8Ilc35oOEzT0ozPyZGcmSe2wnzSQEDrB1
ddzTgEYfGP2OHBUlSJqiMDjvSkvu32D+PeTBtDgKQtvQ5beiVB7qpwlmj8L5OqDZ
C233K8S9tQTshP7rrIhRKwNE1S6OkRfhim+OExvXODPyN4xShSJBLy/3AbDd3SRS
+Hyp47u9L1uOZuagCY6wYWWp+2d+oQmAPrPSGWd6H2v3vqRr3SHHNciAM+inbtnm
YxEL51LPrhEUsN8cXtlOlRrpU5GHIGoOyGBacgY/Bc6Obt6eTpToZ0Q4ciUIBQCf
TGgAy5NlqtFWAcuuVjNdinJ9jdBnphnUy6f9AQsA3r5Z6y27NPZZCAY76NS+bQYe
HPJ+ugRjFCnvzHgweeOGrnsBobZHNK1tbULb4dxUNEJlz5FWFNz44t5Wc48D+UA7
wb1MrvHEjh3+wvBf5Uw2EZVYUvy2higpmIP9pjrx8xZJvPIXOyIMq33HuuntUEmA
YL61FMm5gc1oUcyF75hOIa89B1QX4M8WMylVUsVnw51XwbDlwwffzzktDFsJe0OA
ceozrMj1e8749hta0UyjH1c5zPeQHjcfwZtsb7c36xCLk4m9XLBdUuQ6hGqWfZKY
aH3RwvwoKXVTzdWZ0Mb9W+NI8Xihzn567ZYhqmnRMkXgdrYYK7Oi5NYAkwW6IzTW
dIDOTvrniffU30VdcHoGw/DR4uI0lj3IWAxp103eWRmE4oEBFXdJ34wSIgrA1bv0
hceJmYo18eUIwS6bLD5w1E+SPOVl+P5ti/XpPTZ7WPcPaDtY1x+/uCKZiaM9I6ly
V8AYUgQ2sADuXN55FkMjn3rPvPwYm+z2I/GEe4hs7Q+h5OGP1d9hYGh0qTAxkKKd
QQXneaCzjqxfqs7bSmUMLhXwaBPjtj6FYm4j7NFLn0OCKCrJ03meAVc7cI6Shkvi
CAnp36QihTAYFzH+hkvUiZCbf6+Yj7yjU2ZwcGCSHkE8GpRlpCF8pl8t1Z1HkWTD
cd0Ssoks7pdeK7vm+PYOfmFXXQ0sd0btt2h6sYgHPZ3NLAEd/mNaBhhbffmCMdRD
TrrK6PM66v5XAmv3Es1ThLbonTp66/0fdcLaUFUeDx5Tm+OnHW2TkNUOMfm7BCcr
rnoKn2OxGJO2EAaS6fhW6f3BoeUz8AuEb2wPtC/nNZ75DvscFv5sj2ZFqW42lM6g
L+KA1/Iv8uYXB/zxnG68x5+xaKh9dw73xHtxb18CkR6cZ9ePmXVfOgE6pBOPy2Ew
u/rqFKZIHaDupZ3nOtug3LxOfP9jSzuedMzc6drqefU2x8wvIZY85bK/UYekY60Z
KpFMA3EHcjIrb4HP9q0C3bhsvB7ecBqsbyhtMLIeXSm5JemYKcaiiKA+mThsRRFO
tP/4EYLNUyu2T8xaN5b6Bz6eCwtvl4zwYtBkw5kgPxPkVuO13FBzz+GvnNmCmka2
2Wr897/Fug6C580k9h6M3f9W2hfKZJ7CjBlbUQSqY6+3/1jZxvJ8AmnAH9cfz1SA
+Vv5m2Bhhr+80pjN0GikCq10a6J8NhKN4hTJEeuSynN4VD3H3o44bCNySAn4CmXe
gBfK3+VGQxiugh5kmfd2ThOQqqSpp+/VEhGQEYxOyNlCQfh+AdG3LkjHJkYG89Qh
FvEsGAwYrwzBWxChlZU5xiYDaW5AHia0gTcRktYDKfaF0shi9POtB953jQi8mdRk
paeFiQ2z2sQZ/m3+9cFqUJ0OA8aPJ4DOW3RWE549SlTivGzRtHdq5F0bfDT+KBfa
UYRp+gne6teCZaRq21HjaheFRf3JChzUssvOXy4iqu4HmxixVF9DHpqDeo0Wnb7C
vTgMh1U+6epviAIOy3TcyZ1NoX3hheIITQ3VzL+8Puu3JblK8Etz+yzu8ZZwFmoo
G/47yArH3Myx8pkzJuH1XqiphQaQO8h25yfGIMnh1z3tMYEBYjxAfxjWiWD233F/
Y/EveYkF33CA90Qh4gtmeHncJ+FAFFTS/JyypzAtyPqT88bKdaRiKGzgX2V8DE1D
J36rcwRs/MmEW459HTKeP7jUstn0qfFEbcROX6Y28nM2ngFos+ufA8ZpaScTk7sb
BD0mL2SFIrgHxLuca+rPzsS6KxGKNKiiRZ/UIli/lsVXwlJByh95wPUqeIWklPGL
S6GIEQ3/xceNQKvA1srPRqPdqUjde9aIZD0Z+Ujtc4pjGqY5LkHXAVGJuubV70pR
DjdfCCUaUBsDQvBTIwy+uRZkGTzb4muB0tLDwnoa4sXTm/r0N/U9OoWJ6LG2jxXP
NYlpOyCJItxW5PkfblHZPKAGykU6AOpLVZLmV3BzCnMIxTk2EwPFqWUa9VqRGwbc
UtKlhWz0wy6YoQOEE41XJbJPXbC/DNAWqMTKLhHastuTjS3RpLc5ErIF2IN1psDa
PzNZ9C1hEkQ5ZmwY/icMNlPJwN4wJAQha7rwTrcQ1kzDx/VwbW1FEwYJjxL4d8mW
GIGxh4qePykVdUnwvZJlG19nuC+4asORu3rRGhO/mA4jDroU5mb5vHqot2HsF/A3
YQOIvWoy2tpM+fkNrqa7hQRddRD4L7JzlbwaVNFSW5rtyePFnTYKIi+k09bCA2Kv
u5uj84lCNtkFwBmNgWE4qQTeOZy1C/1EgITXJ8k3NahoolPQ3rIm0dQKV3/WCxXB
uMu+E6dQna85KkmAe3lmRRTWEnBziwbgv8exFkm6Sg+5pTX8jFSyVy1Zk+mEZWnL
vjqPR54ufUoNiBr+Lc7fQBEZxh0v1z51V+fmADSkTGjHxwsnVPZ071uDQGXLdGP/
jRxnoCYWw00Xy9My7gx1a2y5wY6OMPQAL8ndJ8ITRi/74VQmRFVjJhdBkIBhT+s7
896r4epU9l79xR6zP61BRkzIMAeOqt9RlMhZRsgtNg5NqMkC3lM6f0a/+P7h7+lD
YKN8H7IjOK1p6m8iBLV0oCd4EyKHkaY9fIO0LWoUQUNSH+940kugCQuJFnQr9WJx
TIzLp1Z9FFR8EaIEMFVsh/bDGcbwjzJanQ8kIcjXj2cdc7jZjbWr4TmxovUOQqKI
wXLSaE7AMlkMVTLler7TDLOGlpQ7aX95JqG2MVQhq0UjrV6qPq2b+e9cYc3RmAER
6JX3hluZe2eSm+uIE39+cK+tmHawiapnTmwrUTHiwOqfK+xItYfOJTTNOdWmf9/m
agZusffDNEUxt/4TbI/cJwtSgKlgnlk02d0T1QTvI/QE0eIYiFuIAErSeVM0aonF
4yqC+QtGicKBszc9P8GFvQz+BFct+xWsW2SyEVf6iFIIZGwpeQYw1CfnO/t69xWC
XD3LuQMfDK6EE7eQDMs03vrQGe0ew0ICn0puVxxTXxY7TqGtkzkXl5/Ahl9H9l4n
K/lQTxCy28UCMhYn6fCzhmBuPGEbzUqBkmSIelvzpZ2KSt+VDylt5ut+91reHzOY
YbQWHFGUNHx3jHuXcTq1/30Q4qwM/Pnne4E2bWOXdgx9Uaodheu3cbCAlCAr5XpK
4ouEcFIqCQUx+NtjKTjlo62vAj4xs6CQndh4lRrfh0n6jteMMrTvp/G8ULecUV9q
o8XfsDFR91zwl5C/UOj8ahCvZ1NizK8KKURFxBzT0F4vRBNEoRBmKjfHqhOr8xkP
xwZaTp+rzKp2DCAcSIHvTeon0Z6wcw9pi94B1ZrwYHpXfocbPWNhddOyZUK/ZKXA
tksrhnedcJKkni719HGVvIfS8RN9WZBJiZCAkBTToAS5ywtciZbtzO9DGHK/lWyG
r74jUNPsE+9XkWEJgyBrVE+9uvXkdAABhMuNajOG7GaAcKrY11eE/i67n15A0BwA
qtKpqF/EWOcSfVo84jI3xABighjl+jgVzmO6xb3gYYHUvBQylVgeP80EeeK58vUk
EH2Q1COPi06Wo9NJz3hSOyyU7zzT6TVIRERbHdumeAwOly56YLZGuBGuJ+GZoiRQ
znHjdtidYh/oytTBiCZnWIG87hrKm6/pDhHiMItzgXvo/UBFAGRyN+Yoz6yLrttc
+b8TVcFhaNRe24nesgff9hrkKfmZy6fL0EJJ4dzSFJyoyl1X2aMIldeauDNiLr8M
GwaXvtRzCsQDqWks85LtfIKvg9aoG0iuArnGvhsS1zN9RoXpjxdquafBaUPXjyVB
LO6EHbSBE/H3F12cNb+mh/vBHYbzZf+ao69o1vTA5TNFd73T6O+dlpo/bQh5OU05
untWSMgkkzssBnDOM+Mq1eyChTv/2QJyYXYrW8yi2YIwBiHZQu0GpbgZKkMl83ZC
JlqFnxLJl4x0sJTRaAjUT6/GPBzjXQ2/0IF5ksrcxxqaQenHLq7qSz+CMFdYWj5o
Y7SBjmzDBtu25LwW3mv0NPMIRh4TLQsHEnTw1ld+XAMX+z1UHev7PMwg4z4HEfaq
mQPXd4HIVINQPhbFbHE66ee4LXOjLzj4C9k5/i7ZmlHIJI1MJ1CpPZ65gnOEGYBB
20KdZTNxKd8wmdsoYOcPRStfn5m+3afquPmpPJYeigXT7FjggbJPJFjKCMjA84Sx
stgxs4ygkpTnVfhVplGj6Uu7AedeAtz1swqp8ONnHSiHxti06ARs2qNbipOBuUXK
+2apKa3VQopOGFpe8/XkECM1Zv/WUQuLtbohYWnP09h3LLBfwQIvetu5Sq8PFJQ5
sD6L0UQ86w2OUBfAJ0UJ7eq/lU0DTNIRhnauBy7zFi7ztJp3MP+Z0QJXddXOO+ip
dpeHt+1UK3DfjvMEJrFPoXxms75hB6huAkZSLY9TUaMR15eGgivv72/OnArH27gJ
EKkR6iLBz5ZJihRsrQ0TQy19mzqLC/vgVRyKV8PU+j3afvUengk+jRSpLc4sXtuU
2Q+4nazeSw0bpbcGf3SVb5VapqGw9ZEY6KpvC7nNPF6oEvkqvQfN3czdjQGeWXfv
H9lcou6C8xVjy9WHtF5DVYVCdFEs+69650LwCdtg4ecljHssT53pDMRJY6WIzSmR
VssUggjCI1cmXHYsCkACdGVWMMhvLCiVs2QnQJD54Zvy1fxAQx8d9UOvQON+sPJs
pZ8/UHqMDUn9vJulsn0WSFhCkYePVrLbe0DnNuiRSkk0f1U9o14o0YDMB8ii3lV4
r72kQ533HOp2S+sMfhYLJvmeOF7/OD7U3Nh7o84muKuUuMoiT3/szWKeuL+l57MT
I2AzEvFUEGaaXIXG2HK6+BH184JJ8wl8JIHQ2Ocmt4jWZ11KoZdkd9YnqzRbhHcO
okfkh61vCiuZQ94EzWmjn+0NBtjvpRJNbWNjU/FGVOuidSLKk7jWg58gdZVSRlVg
iQheC87/wasYSq9AltigPWLpSkwMNGSJeE9NFBptc8JYTNfjgEjTPO4SbzCpA+pL
fzJR3YY49y3V/NC9cwnjHXHHhak8fJy/333FPUf2S7NlnsKMFyx8PHHFlbY6F7rH
MtVnZg6zKZQGlpZsKS4fc35gKgDy6tVuCmL3yRq/BGjPs2twUD4YDgn+ati+BpQV
p6hGgJ+OjKdV2kSGZEv/3g8VW4ASNYbv4+BVTeTIw818CARpBRtQhq+B4KZNuwx/
RH4nlg6nlvgCovaSQe7/fMri3VtUetZrdfd88TL7bPs1qIMP+/6/GN9bQpY7HLFb
HH75hrhpRAwh+3cK1Wg04qVfB+qCj09/tGHOeAovxKllvkkJuqeEQ084HlFzIjTm
LYKujn8LosRZICKFHBEaYneWe38TqxEx1R8hjQ0wbaujgg1dRNCtSOrxjUqZeMIY
rba0Xn9RyYR9+oPmYUniyfKrZtjkxbgUiom6lXpGInj2Q6QpO10lfq513NzVQ+57
LpdZ1Obyjfu7RNiJ7bnz8Lk8psC5+aBj4W5V2uiSGl274ECgb1qb2zIT04XyzXVw
9WjKRGkKbFkYkV4/0czAVP5HrMX38giSdOnFcXEU5svDFQ7ol0cFkcUIgBs5L/Le
2QgbZ+m5/1reiVpT+wN11IDoDZTG5zejfV1huPMPvWTrlVWBmIhiiFA/0Z5p7/t0
sY5LmanmAvo7Vy/KXDw4XoNCmLpLtOz0Kga7PSKfYOl98NrkvoU3AQwLKbt5HE0l
5e+XbhQ+t28De0IbgTebpxJPiVCiUSHtMhX4bEX9rLEn0Y87g3uPfFwtIpa8xkXj
MHlNUiaNxLJq2GWV1F7VbyI2xtyusZ0wnWihyQcLQUCPafUbaIR1R1+XIRHsEeL6
MvPMx5TGoN6lYuYU7fp5SvGCeLwjaeCf/IPLa6URLPkGKneLufBVsco+9R2HUnsC
71Q/8lHu8MU+5DC2neLpQkNG3fi9/WSJ4y6NciQ5ZldKsVwOmgcqXGRdM7pobI00
4FFOX7xp/wIeMtvroAiuqsZkdK9LyB3jRGoJmlIL0SCKLumhj7jG+HA0DZDkGt2P
9yXjfESzdwT3S9z3BteTdrW/6aPp5QSocOSb8gyu+sx6hT4nNxHi67l9Lff2P8uy
tjk8+1F/QVmzAb5bCfzaoLUj1c+sJPbiKmYT2SWZAGbOAVvYTDKIYEYOPUKhfyQJ
oSpZtUxCFRnxl1ZvDwOi11EVrPNEI1MO2/zd2ltDj3YPpqv2pV4MKb9yA7msRmGT
jyA2ZmKsZHkRBDE257WXL5NYIBAWtOwuriplhJeJkXO8YUztQCCJ5jojkcPiOSSJ
iW+JF9PJHd2jTB3oRG4r8FpYsJ3NEmskMctZTz7DOc97HRDZxdMuWm15/BFmSNPt
EQgMo/VNCs73FMjt5Nfz5O0MQ6lM3iwz43Lpr3E4AoBcyX34+nylGSYdalRfw2uU
FN2ruIPG4dwVVy8nIaXKNvTR6O0h5/8PWH/zBlItpd8EwJYna+ckKLJLAzcIZxNN
12102ncOlPago+JjAULToSM6xk9oLF7/IwQuYcfaN9eXgP1N07coTqwGBPqL1EL6
DTnBWGd+BA1u1hj/tkmfnwDt1UWs5goHzNwEYrbMpMK0KYCO1aGluBfhWgs7ahwF
PwzxKcj5UtYQBQ/tcvUhC3zkSWd9hBXMhPvXacwLX4kyqLTFbgjNhEJWRgfnI9jn
/cmRJSpUlnL2rHBTf9oz0wTrAxhhgqXmEqU/yaoxRk6Kt7/g2KPMbVPGS9vER3Ea
8yMmhFe1C8nBpmQOGugkyoizPC3tX1854jjdlN60KImQzu69K1QcDIyLGzFAUs3u
1f7a2IUyubcKAVBgaD2s13rNLcY1tKP6b1iYYgBlxOJHyehn7zdQS7zLxKUzJIe2
BXf3RT3RQqW8si4yeWoRFfo19rQEs1y9V5bUVo2q2lLYRl8ogroTqj6x9Ibzrns1
xdZSJHuJ1fVC+J0m4cd6mntJ1sATiLNRUvhBZ562bFoMJhpUhz0JFBpopL1Itcp0
k20qZ6A+8C2sTSDiHqIQ0wuuJ6xFYrMwWO1lEY7LY4WtNEvYc2MyjDXZirFFLfiN
WkX9hCvbG9HcLoU4hkX8mSu9QNTpH4JrN9iNTe1mLBxs5our+VjlU4BGtvZbB1bS
RvVZQdxAy3Q26TUsl06N5Y0CbetYj3UYfUsBeM3rNiUgMwlcxc0UCqOx2LoSM1Sp
XtSUU3ernEjekKIJQoU/Rlkj/Ao0cyjcVkke8gtsy0h9Ee5Xbb/pIrvurCTcbXmj
7bc7Cg482YRUwhT5BO1ZvPoeBkEwqqfWVVhlNZCJb3grZ2EGgSDzMx9a7Z7PqTbr
M8n6iKdbL+WGcELJMoyGzwjAeNwFLoAcdUVkesqhMcLWhlLLEn9Z9pBCp+SVCJtS
3xDTONU4tuFRRhphdPgLu07ViNrg74qEROQjxuu/63qNCMX0VdLdH2kbccJzYXL+
oWwIiI+PVpzr/1sfiS3gSGuQ9+HOriCi5zaaer/v8QQlw5up8tyusPJyF47mm5pX
TtlTDE6NiNJ+nUOlAmCn454QmSfWUczkakPsbI8wXPnwgqOQYxLmNulozKxm30nt
PmT05wMRXd/X7bq5QD97Wy5JoLdNKdeucEyHjM3zfNj+G6dJif/4/JyzM+GSnOGG
RlDnCyTet2jwajk/l9T161S63feyF1hOfaoLHpeyzTq3cp1fTdoKlvadVvk2JIQt
pc46zVRLn3zCySZdkW81SjiUlr8Syf8xvwFYRg2kngVut+d5XZ/L3Hi0Ve7e1BjT
6iZHML/FH+XREmIVwVe3KiYqidsuRCd1i+dOXp9800G/Ow1ipxVmx+HNBW6jZw4T
RprJiVL4EsncTCdT3SzrxIb3bYcY8PljdEs7QcK0X3irXgO/6w9CbhcPY+8fXjFA
2Ijcdvfat5e610h2v6g83VGWW6qg385Wfy21nMVQlXoEqVFhQVyUBmFlqrReWbMA
aJ2FTwbEYH2alLJgPvg1ZfKXlF+Ied6ULcxu7acgP3Q4T1jp/FPQCcmL3Z6EA+af
Qtf9Iy/VRRstPNHczbxLf9uNmSCZwo6DO5vR6wLJqSCPh2dO+XkYFq5+y624Nive
BFvSmLUGOaEgL4pb56aGDoyOeOV8BcNPlrYukITaBIbZ62xKtgm3X9xwA9WIz1p/
X4/oWgX8eXR04pvw608W6MNeeITot5485EPmZxXNFHtOQusGy7qHItdX+OgGHVy9
K4ZSKJDrOHAxhZYin+GUzcv/qxQO14yVSKn2tTvpQQuOo/4ebV7oPfdsrCAbUcEZ
NncUEaPnfJ/L71LmZBxlkFQKjiuzQXksTvr/RrIJYJYaSoz7PjjQUUV1vVxHObae
jFiuW6NNKgmj3te6Hhwb9EriI8U1yl/d+uORIRFiMRzoFFDSwzrobcGMcDAhyW99
wQfenmIOrAMWJreJeoplcIwTu4JjuSfgMzAgkzSyTvoCbNnDeCA/xuiEIKQVqr6D
3ux9fD75KRCPF5q+EtpP/WeUCVnBB5mGv7JEBwDR5NBXVINXaUXm8x8+w39Mshec
qmAck3IXMvcXSyFj8gxSkBOxZ+drZxlEraoBvdVyfR/1CVds2t2+tDCXvwwphv/S
+ufwX5PlscxYvgbHXdmfyjj+oXzRj6npXTMnawJTdjUoqMDbOPty8gwKLEMXGu8z
yK0eMlXg5n08qEkxmjCESRc3oB4zphuslOUFIU3zNkHBHLDEpNBd8HSeBPE4B8iW
C58KNlagZ4vZEUVKlKVbE2wRFFoXNQdTPHUKg7oniyEhtgBQwSlMDG07ak8cmw/4
sF3BWm3HMPisoJWoWr6BnLxWSZEBYimqR6gwSqwXUdsWywnBagC2qVvOT4LgvxvQ
GX1YtGfqZmbmSP/Hr1U86fyrfyTar1r60jLBRDmpIpWPQAHWeviSCzivenlwZGuM
aEzgTUiUl+vCoGK8jfn/9Ssn1JWfSbVU5msBIJ9H34rmhjfpXor9RXQnZiUVF9A0
fGEpP72yCUzM54QFidFrEo9I30P6vNjFxvpHAO+A97+RpVtV//5Lb2NW4Z1IXvyp
+cf+I++o7W7hzVIWY09mfHweiUGF+3jGsRb0DpxkUKnY8pMtjdsp0q8lXLGUqthi
L8uNpXPV14STWJdtjMhQCIEg/lT/T6i4HtCpUTB2QyW4gFAzaxaHAJxxfIyiOc8P
eqYUyNPaS++VSu+SPDlfJo3Sl6YTtOqhur9lcfI49HX3cjnJIqW0mrrFG7rtJpD5
ai0gymgHrBHL9DmyaGevQQXHhgoBuXki9luMLVNmwRzhdTSMtlRAApCYzNbgGHGQ
zXG95FvFiHJLIA+KfpuUl0Ayl8ZaZmo+EkoBH1lCIALuLEapaP3Jidku33pgkKDL
HSODtRc7oBt7nFjk5ZaaYXLB60uQppG6Tdz3/XWB2RA5aaEU16S95pSzTDcYhpOX
XWC7IAKE4E/kEY5k02VJtBVq5rGS8PjNeMqZamUmnTiYvX6fRa/uOhBDlFmM+HAN
VbV+tQ6a5TmAoytQekqvslWbHV3zUQUhuvKbSIg58Wu+AleW7xPRcnA0HRtrWes6
CxSZMjql9YoHrsrUs90lHEdDi2HLJhsv5RzHt6YBeF6uu3N6j4pRBVK1zwIiBIS7
RseO5e7jka68wwN5pC7yp6t8m/mDG5TBJGOfK6gVUWF5XPz7mJLy2o0Yc+Fl0J6W
R4cmL/3Emcfs5alt7Tq2557Q7Yw03VRmbYbAX6OCRV25htfsOQRfbJi+uF+fvUij
7pj5vG8/UqJKFdUFPbCa7bcUV5nCUK3QYs1Ne7c6CG9DqZjwRyS/NkLTPCuiZ4yn
srTtvnHbAEku1/3XUbc4jzezew+pnRlcsn0nAEg/RsRc0++4atbIy2WDk/9Imdtz
k7ipeBY7rpdLB1SV61nR9bDqFmbY3MLnuC2JZ8Lxp0mqdUojkN8Gq5bJiONbSXPr
5Csnl8uZGaOZw4T5tKJAEXT8gcsOP7Fg/ND9+EPMf+8Nwprx3Qn66OgsPBMbV4wX
1P4s52jrnT1hVzb1PIYZaPpW1eai3DprUUIIurmzQ4MFvKYiN2deJnE11TgciYD8
lQaGYLE+J0WJzBpwwPm6tiy+zuO6ILtC2s1hQmzxokIvwdtECcS+PIDBOcfrA7ZB
UFV42CCt6BeQpbJPKehwX7LtATRh9DH7CQ7Yidyjd7hRgynLxUHSvnGzu/gQBZt9
B/eLsiPhrEwIyhKiyxHs4N7cIbWCASkjgN7BOSpe5uJmgke4xAvFnUuJu4HgHpyB
bSQr7Zk9C9qqaABQskj38Orb1DUAcNKN6/DFI2vXYTjIy1nxvCxkP1STIHTFNARf
15Yb6bQRkbK2GVXcgqHdBFn89z1xmy7bf0+bAQX0a6p9iim8oWQk2ZjVwxzA382Z
X9/0TbhKT3j+6S/xt0NpYNTarbrOKyOReROM0o3gX7XXAFqvhzGOSVQ3nFXXEASR
PnHEQ3gKwI+JFDF+Gp8GWCvZKQ1zNl07DX4ik95NTOQolRoNQN7Uscs5ly15phIR
Vs+j8hqR0n8SFePRmJrkdV/aCVZ9SXUzqvbaymQZxZVWXAFKFahUQz4NcBZcI2OI
KTjQhX4EdnjBz8fG9UrBwAuWkSKTjoeQj0Tkb9WT0w+iiK196N2WixSYkeLD1lUR
Xkw2O0hotXIk0hJ8i9021SF2lpvbowQ5o93oq+wWn8m+TBh6+H9SA9ONyINhYmV5
skJtBrcCEOuBUABTyQ0l9C9PXuePYTS7QvPKd9o9oz+rRn0srmjO915A2y/1hqIf
s1iC3yzL1dTvEjqKB8xEBenRnMKB7m8eJJD8MGUf+EoYF9HqXhhdSzkEdRourIPG
9s/m8IJnfHCZ25Yft1b9SOqF2oHLkEN0IekQR/lcfQPhLixDWJQ3cV2MEPTTFzGh
8iTL9KvgJe7nlzL8sqe2VPyVPB2564KTznrlysy+LboleTbUeLx7soOwXdPpeiwL
Z/vQvsOnlPQP/Gr/28a4pumKS1BhKVviIWqCazjdKWBOMDmvWqrx4DPtbn2jR92a
3tJAaHxGz6CffofteNhkwa+1j1kwejOMbxp76C0tzfmR5R5gBk+tUSuvm9YnxWFV
1QHGK3gcph3i2LAyzoqNskUt0l7vP1ZIrStdc+pGXMvIT+EExsT3ceq1XeUgbqoN
BqZQ69Y71cmhb0OEXAEKZbVkMHFZtLrNYXncJlrAFD8OdF6laxIGOzbIs3duijG8
v3D5lJQJyqlJygG/v+MLF0/fNdFc2mY/BHCFAnLNfY9miYxkl3rJcfkcyU43VIsf
1JN2o7LlTmcDi4ZM9qrL1yjim1PTgd3QLEHIHEohg5ytO6CT879oe/CGcptApm2B
GK9izCToGFf0z5yeD+yUkuJ0SZq3Dgc5yRz7NzMUlbS661ABUSiCgkFyE96Xs1F5
aGIwASmg8sKEhFR5nz8VqDApIK+II3yHlF2+kPx/stONlh7ASjLrCM5E+OfCt9WE
BNizOalcoJDaPSrZzv/sxAhn+AjYYYrJev5XD6nneBUTbnmjx0iENORqs7rNptew
IfEAtzZzzjBA2Yh89Ltfm0fEQ9LIJJu1qNeUKD6Lxgkbp26/IJik4zh5cw6JHsHE
9ju6j25AzMv+KKxilee9zirRLoxWvaXAwWcO398aJYZGGBo5Gt2wopKYj5q2wM2f
naqzszFmrhaxxBAVhwd7LhlOJrkU/ocVR6xa5JqsuRHpvkjGZiJznVdy7AdW5E9Y
6RtrPgjuSQRhK6iFf05J2O8crQd0w5acQPDz6nz1Elv77mAHps6GUFM3rA3gNdgD
TEoSma6rZnSLDA8dSh370tq+WFqAk2YQ4rpjOI3V+r846TBTp0p8kZ4TdRbAz1ln
iUgCu/9mDqc2JWx2vRddZ6z4qO3FPNLTc0Jch7uYGvtSgcOjogrHqWd19jt9tPpH
TcwGwbbD1+ZywGpeV1w5/gGVbMDa8XWWdgdug2n9ck4symPfGN1n5RdfrJuS1FJS
jb0xyM0umRZH3CnhtiXeAzXvLOacQLRepIEzpxCAj6EV+CcaeJ8ENcixWMpUdYo+
rA5R83f9DuG5KvVtcp+9zJVB6cgZ3L633yH20I2vZgY7z/OZgi25l6t/53PBumyB
llEvsVW7NZYoWNKElcH0V+DmTaTiMNhFZJf85jMBA8Ojb+00kbVa6Su9LxNK0OTz
FLl2IudjaE78Dn0FutpPQT/gwGtSAnbwm1C8JDXjK3xw3p4tcaL8SXpoA9Ahnhk4
aGk0pSDFcqlVhcmIiHMDbaDxveXINK/7y1SEsXz65jGFYTggm+iJZj1RueaEx+IN
5x7C9nVUB7/kymx4HXL7kS+eqB5nIwtni2Mwo2cn+b17vqgJsxoHBfcms+OjCBRU
FV547Rpn1gHwrz2mXGRkZcz+VRMid0zZOy6S9m9/F9iCdrbrE/nXVJQhbBBHTfCS
JwuMAMhMs7GjKA5/CupQjtQqXs9t09qNZMgXqbUsZCOP51wE8myQ/wKGZUFzENvA
SNWDf/jU3qDcwOCLs/DQ+qI9VjoYS8D8NBf5SPh9cCgmxdneNSIAFOsg3h7FQopR
zn/Q1+SPGTFNe6XyKFMpezGJeONzvAqzRr0/fkhgEhHO9e6Tr6eFrniWHs+hnOHx
oLSpvdWKsLqz5To8zQDXHS70I0tnc7MPA7yw0zaeGKP8kvVkangvDo1XehqSMp/C
nSc/aeq7vyj26o1n03mJik2cG8XuRF/X2uViImjMdIXOHAJpunVQehjVPS8Zm3oA
Y4mKMu3r5JouzJ9ZYEHjO8aneZCTXBtKO4G34tT7/VzJ/Xqs77+PdQPDhiD2IQir
2J/vJfEOXD6096HPCCxIz657dneaeMt6VQySf2Yfva6+PF6lxsR4d4VVETX9FrY7
D8kTNDOl7MHwc2I6EbDQuH0GphSBbzX72Wgt5iQx8vxRz7XHz0SyoHhVjLALuOT6
T3qQdlcdLEu9PoSMPCzGjkrrmKAz2JQCv01ESkFaXxs/0MYSYa7mQcUa4IdXRB3e
kOzPFSBTZ1AR3Gf2oDmyl4TMMi+lGbLSd38qCKbEGOzgYdKdb+U7sv5kwedWP2q/
cgFxbxN5LYzAQiCnPJw0hYviV2OYYko5oi09E8AI9B0jITpW9YezClzfyJuXLPaN
7uq2IU6CyBAI5u88DdIlIW+VwGjGjovWrAywpln7JsFpSoEX26GX9XZb15niZMIJ
VEY+vli5sDFBgDs8A+VGo3Wr8Sdh6Af9xFd04dC++bCyGL1XiYhcWwmBCw/QxxBe
uICM2ztPUkaHl+VgJaxde/5Vw3y1pbvRVYOD9EEkj4mCRDKS9usZGEY8c5b1OXtJ
SHDY245uqlrF1KrGbfaXT9aJiHdzitD/4PmIeKFMUbpRrmHK6mfHvoomJ0PCobKM
SZhtMwNSGWIRRPlQppCMu6Wvkke0rDfw2MpPsMRS4ZY5C9LVgo1vdr1rcxCgFeLE
sIyuTWD3INvXL0JQbAkeBcXJgiZedQNpY5FzfhBQbxgxx5jdVaTIzMTT2svXW3Kr
ZBMnV+YQ33zavQsdeKC8brwu2COPbwpVww7WWjR7G7P/DkSS8SLPpDkElaVDhfDe
FxRNKKai30IP7H8A1ot/p9boji25u/Bfe3Q4fdL/0LuTt+tckQMDaDoQQKh8M6KF
quvDFdLb+0/ZpoMf6ZTplbr9SIQxEalVVHGUrEngLboJJyMyANziCM6oPYT1D1LM
BsCuKOewmwNhsb81FseZwNqnOSI3ru/I+qj29/Fmt9OBHIGqoHGLO4zzc5Z7RTiv
9k1E0snSTMHZN6yd1povn784EQzVXEkITqB0pgZVNZCcBUjVOi7lN0Lb0A3v57tL
rs8McH6Zzdhub+jZjyoG4+FDNFthvPNg2bvs1LaTGYCV8PzSGYvI9EKXnbD79ayH
+bSPKeH5hQM+rFBB6fX5Zj8+KAt2Sa7vahkfjsw92SWJpcrKcOavO7CvFEo+sdDy
0PUurPhCkT9emEKeI0ItnKE9ARMA3vrpgtdpOVb8uxUwk8QAiFvG/GFNRHDRMfmW
llv2RnTM2fOBKm8ZCrl6LMgqZDuvyDhRxIrm3nhEJ/t9dNqhiVWC2pNz3ISp0ZK3
LoAp+Uk6SBvSjG9SvS0v1m/JiG+FEHwIoPbGBmGxTjUr7LM40SCDLCQhCOTlJgYU
T7KfZmpGOV/iv/NBNUpVEbbXfrekIcezqNdSv9L7cpMGuEcfhPzjvK/GPJoPbtD8
SZWN8kbzPbr0ye5jcHDPSZDx+7zDwzvl2kFT/E/u0y+U/jWKeZFE/semgdoQoU9p
dvY99MjJnGMwQZmIxjKgoPlQV1MkG5I/Pvng9BdUV7iw167Fgj7vWhOzwADSqW3F
SbBOrxCuF8DXiK9sv5+EX29qM4T4fg0mtI6f55gZl9mZ9v+aJ1pWPd+pfoyRdKZW
7SMmW6yTFxmRjXd5lhmAc1bKpRB1WzLVqIe8gJJtXM1sCX31imLBfQOwGI4WjkTE
oKMlj+5blP72OqsXhBKEWTFGMlsOICQgpRPDVaxUM8T1y6tvB/ND4xxoaYXzbWbX
1FX5MY7DpRSNW4jw+6RcxdHxMniiuqFHppvKcFS6XW6Frp7zav38PRP9sLrglKXJ
uJyVw5Vaixbnd5A5HgDWtgyHnzVI0nMlbl2tAtEhFAIWvTgr7cy3X+JoXckprKRQ
rR5+t+qS7P/bGlVjn4QJiy0JMTrX7Wa1DGxRDs/H8L9s5R5SvY8K0fNsezGBJemU
wzJoEejxAEautL8Kk0whoYkhtSA8gbGgCpDx74kOM4JRUGa2sTunLZ3CHBr0NlMF
Rrmcah7yWhRnIWfmc64BFbuob+As2lEJ95g8Vd+kqj8vFw7/lTIz81fhWzLHsi79
ZFAkiJeugqlNaN1glcyq1gJB9RSrppj/HRRuzwT90K/D0fJ/PSk2R6z8OCS7YIYl
mQ96GxUcVvsF/GFFxwaHYZg24eI2MOqPJ8tCJJHCy0wGot+EzYvzZKrmvy7yiJ91
Diss9WdX3Vbn4D1+PvzwQ1dN1D4Dww56b7d2EQfN4ZSTG9amYV35+vZyszBLnXey
Gqc6X64gdfikrnPic2OAgbeOMh89O+TI/Z4xoLDc9A0knGpzSYFisuTSn5z0cSvR
4ZRHhmNF8PXgzvA9THm0V3qne5jXyx+KW+i0FU0DBMahrFjbLK2kIqKza3XEqI4j
zGES4I3ZsrDd8PgGcssdwk7wM47imbVEgwX1ZHQsKSYuiEFo9Y2d7P8pUZcGgFDj
G7RRvoN8gaaO823L8wYc16V5A74QKdYZRBrGiybSgxmKei+ZBs7ySNJZhgGwRbbM
uc+09DeAGYPGcepsrbaxvrSoWiwoMGeM1U0wkg+2laRaZ6eS5mEg1rBo5asFr4fN
Dq3bCW+9y2U4F9BeSvdHvTmkAEX0olxRSt3nspFEyDIm0IkfGaARf0FPBAmzhkG+
oJ7zNGK28vzEcBD9StPZhZW0GvRcs1+FwiVDyqAMw5XTcp0s/yPtNOdGLkw56ECA
1VgjbC9YVEi9bZaS83t6XKQKTz0RhsK8tE+icd2OwdYIl/5W9nFq2kSr3DwW5CUh
CS0QGObB1tK/bA/t+65hcyOlD5L9To4DWxkzISmosKkAUIIzRZ+1pzTg54E26mRl
34I1xBui5zBC7+5ctmGnbGpYBwyRvtwQA63RvtHQ7UGuh+7d2xZzv0KfOD3HVxRe
ZJvvcHYWV4JxrM/bSlJeAt4nacqoPwtW8uzqvg89nkHOonNaLl/DtujS0LjzwB8L
OvRukS/gG3rh+gh3a1ho+JNqUNe9cMwtZcjjNQuJvqMQuk4NMr6vI4Ei0oIJNF4O
oprgxwkq1hdAlkc0aH781KgVBMJ94OGOr65wXJ0bmsHKC635qi9RcrCCoFSjNxTx
RycCMppPl9ujF8M1DW5sdnykkQi4RbA1gSPmxsBBN0twS4F6p87Hxnz1cuVcC+U7
1BNlDUI7n8ZpPb0U3we3i0hcbnh6StO1z9LPw71DdesrT8rIAuhkqH+L8i9dQy1b
H67VmaeGeIy/5ZoMmOtsGKguxgClPATpJsqFsFgVmuS0Hvm4Qs0DTjCILcC24DHx
QTk3p7ExYQwCEFfCOCshZ/yhm4CbVtcKLHQwauB0C/hY+PzUdHcXpqcBJkiVD8+l
TUzGTM7XlZVfbP74V2eNa0k8G6TpSk6D+luA6X4j1pmu+lyomTv145oYN3sSMAmH
rw4EhT+X1EmX82Vt/NgcYQhnPaSn+EahVZRcYF5wrirMOxN3D3AWPtZY02C6xqPq
R3AvLahxYMyjVG92ZtvRPL8MJkMKB+zbkwxXTMo/hXG7W72q5dNm7NHY3QVaZgBx
addqF03RQLmbFmQgUb66Zal9e2YabSv0MJ+1+ZUp2mNEyqn8vyfrT7w6gnSL0Jtf
gIl5Z2JWhfy1R1JhI6IY0jjbnytK8oHCV+ieTLcp9OkxGZPvgJtrJzA+YTiHWSSa
LFFYUZGBY+UAQ4AR/gSfZOxjvNGCiQJvm86UZRWlTq64alwOQE5iQdanP7mdYNNt
56bU/bBm6QjzwagBwcJQuymFeKHE6zNoB2ay/1vOCnlLtzhBYHs+mt6L+VoG5zao
EumMJXbkeuOXcPBLqfCpt1emM2a22cvUvFPDkber041Sh5wfIn2si0ikMcqAHV/8
oYPKFpSQ5Jpbx7o+LMMdNskWbISjuUpx5KxFddWEmJK0gJCRBj4cHHFtdTxqlUgO
E9LeN6Nxguf5f7qsVYaHto8l49VBt8PRpS5eCQ4GqdzN+UwsAA+b9hWkc1pCB3zf
SJb5s+I7BwnmKZlo0psFe9uLLi1L9Qehzyqudz/dZ7vU8JKrmvPM2YuR/iyAaU1Y
kEOldXCML4UKGkfFhl9b3wJ7e/sO9m6IW/nwFnKM9mKmE2/1YD+moH5Ue8/B1SEQ
5BwKNm84YZg3ikTFZJV794pmyskcKXsQll4LF8Yi8guU0w75mwFZQMCDkCGCm6ek
HxwMPM8Uck63cyCUj/AavtRvJuTx39TuoZENrPYxbuVL+AMlCmqjl5Aou+B9/NXI
6QWGw5eg42/UUo08IG5qxbEs1QacjUOh23xmW6dZg0vlHO59jo/D1jM4Jca1SfOe
0+eqiZA/gUZQpF8rpJCNpLge29GQxG7U3joiXf+zG6FNUCn4raioqVFBTJ2M1STR
XLBRmvl0xT0hSw+pemSTjPyz4TwSixp0te3dfuR6WZ9gV+QyZvdnyuTdkdxi6V6R
g2y1GN4p4Z1beHqzihwI/QNZK+4KMFldIxwq6AvJtxEdQMDhwkVBXiQwp+8X+2rN
sHMK7T8m1qfI02KjmjwNdR6Px7jhScebSCcUqQS31pDVgEfVAg778zIr1pYyGgpG
+8rW1IBk5UjPNzqJtocpPMVCKRrZrdp/gvCaxOTtr+vH1LdL606i62rg2e+01Dmp
0MJmCgpQ7lF5BeUR7yKPOLye2Ngn80xorRMnx9uqCshTNuWTtz4nd10XxtbHpR4M
pVQE85/R+f/PtkbO1qtPxCIwUckvYGCO5IMAzcIoLFOrAoE9ew15MlRGCpUlF0Vo
6ithGTog0RQTntGtQ6/Hagn4dkjHRqZBHOBvoLG7QsZnllCF0KFEsyQxtz8C16dG
cZWDqd5/SBl7ng8zhgqQDN+wXEWTCB07hkciJ73PFiP5hRmKJyb8DBrmIP2YoUzY
6nTcIyT893Yu6BPpTEjN42lFJF/ZqKLbS3XmwMi4uGHw/4cM3qJDjsqyq2rJy3iW
GMo3Y+jThcjjSPblP7XH8mq2TnFmLgfiYEmrUDLH4MSuqbIioo8aNx7x5lAvKoyk
nYLbXgus1WTWUZ/WHv/12eZLUvtR9n/PnhuL4fohLAs4Qc6dFjoKEpEjYo3hVfCC
MRwlE66Rp1ng2zCRA+8o5oVv89V0FQPVzLDy4PgsjcLBEHGXzlpI91A+aJulEKc3
bSwJ6h9H7Bbuj1ZBXa7fO18/x4WAyFfGeqJTwBcVZxbcPbX6TErETt+sQA2GYAlQ
I4IVtrHsXLVSALtnNAmLpbkKtZDlkDqfIuFpxGj621s2dkJoXxULlqoBcm/pxHOL
nZT7sPVFLrjId/uroyS9NhAPKJ1G9JTFTfGHuSkzsjE08CLhjF9dQJoTux+GgwWV
DDk5KxyUIcyHaMNl/dazh/hqnn6v8Q96loLd8fDn8xEXpL0H2my/vSTxj4lyJmZk
ugYJNlW2zQ1zWC4aOwgx+e9tctIiclwbj3QPgB/GkDrnfYrQXbkZrcm38uSm9hlO
SwGUW62oe4+ouk9KQpqrUxcoFIncrT+f440ACzHX/apBnYcdGxY9rbiN/QHReTKN
dMBFirCJYNADdzINB3VROorqbJ+lT7pV7vF6wpv/Q0Yj4dRMv4p99aPUX6WEc/wf
2EjTuoFaNYQjwsUaiwffbuVi0QSvmghJCCDG88jWP7WqxMBGbbTL6ojyOIybTtCP
wb6QxJIR06K44eqESqVTJIB8bWSDn4FLHQWbxd6EeX+qamdxXpUFSbDr4gHLTI95
J8LuQwgiSBKaCCUQ/N6WA8kdAPP41+BYcH1VqFKEgm5+6hEmf7T28xBpHVfYwDTi
ymbQ2EIygyNCJGUcC/a2xJRP+2RlKWFSMP8gEaAgqhMapFU1TMVNAArQFMsm2ROh
/GpT//9OxXb6ibL+aDaj1TFSPMUdPKQEPAzgl1112ZgBKKCu+tyWN9N5tWICrXhm
IiCP0299zTIkJhxlGGjf0aybymfbBoGXGMigdccysPEHZJGmPx77oTE5a3hx3ZoS
RecMXKVknI75GMd4001J+8bf0C3IED8WzJPth2uWQ3cx/wBI2QiLSek8T3lPfkFo
GYKQhUvOdUAiemZK17RRsZ6D1V/ArFPfGpmOKXpz6cNoxAOYWhVAKRh0zUXu+RhU
ow+8++R4la8c/CExDuz8hdcETYbghLlz1583A5UH+kKw8+01k+dN16mB4ZksrWW9
zOPbTuLrlJdjKvWn0XVXDL+A1K7f102XwpPYeQ3ravnBZBSCaemQOKelOXckV0+V
CsmBBTdTAUCCbEu8f9e9F9+gi8PWrktoyfspmvC3aewutha8howRc1ybMP42NOr8
T1Z2Hk4A0te3mhGBC6iWyS2v6niMKObNCKAfWmTtOVvUdz+Dh6EmUBmu4pFemOFf
Lhc5XUR2Q1/Ygl0i0NmZNVmS36O/xokVux8grWogI9ZbrtIEruVKoOhJ/qzkQ714
gB8pDKJGebEd/ZOtEM6L6WAcLusrhnpw2U/MrWRZU4rxdTl3fSiUm5WYArMymtHL
NO9DBi7iibDwmtcQKO5fwO+hGJKu0JUohg7ztrptrrv+xy1AbKyHgK3Y8UpxhzZS
9qHi1+BiYLVmNq0CG4jYbhLtMrp0n6IqMUE2oDrweDNGH9RWenktuIBmx2c2O149
74exG8kKC+gbur4gyS1d5WIowA6G+QDD01OsibeARCFbp66VN4MrUJmFCiSIalz1
SXCySW5e3UzGVcxWRGqmakMhg5b0AVvWkfMC928fKvVbsGaY3MR4UF6aOpPRuJNn
5RErJ/Hl8CKylE1K+v32++TqSkdWFjL71EI9NRA/EyBJezsKFxBDlmUpdzPnrb1V
wwG209wsBOPDQ4PdHjx/xPTkpYI1nojCMiRgTKaaWyfdz3LqYfW0ebeyyQWG46vr
0tY1VYeKF0Yt25k03H9C2Ejsk6QdDttichBkU8ZQRXWA40AJhrSkhKfMMlLxRhit
19Wc/9doaZ/b8fkktcHoXI1fLZKDZLCT2AmK86lFr7nOZFtvrPpCMVBFjU6oZbiu
sUSdIcfm3/dVzifPVGmdWv1ibWBW+13ob07QocImhDo6mxzV7ig8l8U+D/P5dJaZ
GzCF5A/LZpJ6HnL11q0CWVKHK10MIgCJu9rRFa0H7S+igH6Liu0kBSSdvcRDmFJW
ZpeNdjCvnNFSYVylk27qoeEXaVPMGuGDbGDmNPU1q4tEc0kkrPana5+CWH2M8AKF
+R2r+Qo0crrjv9lOnlKelCDrSsieZQ5Hf0UuOSeL4o0F21NgDeHeUQs38aFWwK8b
xhuf78KUBTQwTSgG1cui2Fc9dYFIjne5O/IOaAEYL4WVNWZ+e5NPUZw9xHdCCEGr
FEkt0gBeT+aWQ4CLgBT6oaOZyI1lUUkX+TXIXQXfs36vHJw9Ju/fYXIWpLWgXZl9
GR8An7WDY6gLQZ27ujAnGn9Fn9plg+8MzD/jXABP/Z9Uh0utZAiPpMjexKw8uc8N
QEPUVSB9/bIYfTHSDlL/0VIN7M5GSNH0vY4ECByJeWNCo/n2pKdVMxk6BCe+LieB
PE1S/AX9DFJjPpm+GE4yUOgPQhWnvrrkN5iNtNIEXxBkPCBnToRGtkflp211eHup
mbKbe4kNmFiK60kyoMRkEQTLgh+Uly0yKV5fRYZ1ACNGoRRe9Khp0eeXOJts7dFK
uYWyo7yX1ymc7jOpRhHh9v5I8sGINM/uzsHUGMAY/8xRe2aGABj0Fr0MB80g5G2p
zW0djZL3OvGyF8ZJ2vDylF+MfDTFt/9YkAo9E3SHqNFXCSerr/cRy+YAH2rc8uUX
bvLFNuSMqfV+fDenkSH6kJb7fRtyM0Zfw/4u5iYHOTewNmFyD1Lb//gueik+rVvi
MViPDr8oRfdycGkIYa1Q5SO1tl0X3Ml1Hk0CuQvm64icow195MQWR9nC1Qj3iF7J
EcRrJr2SaUnwZfB0M+yTtX12hC0BqN7y9CI78wv11QRSzTb0lH7MZo0NzncCNQLe
2iNWHqDhHFarZzM3JwfnjsUnL9s7PVQSz+yGNydy73u6608vyeK2ps4XinjQ3ga0
R8K9CRLkEdeULyCjEWWXNEAekzpT48t+EcpvmMAB/W5h1f9VSPJ3XzSGzYYvhM/9
xMafD6OQqB26oe0aCJoowO9VkA2ADYQXRLtk489JZ2vXZFapU8XMuo4OH4iIZkpk
kCmXgbm0Qgo9z4N95YRECCfLnXBnNXNx3x9C8pWEtmB163KRBVDlIrowAScdw3k1
bcyMr/9iVg1JOlj+9yn2qkHvBV2s2sJ37zWNrmrAgXqFtn7nFICWYt0xd2tt3/ih
jRR+cOS79LNZSOSPTCokcSBbs+CoHB73IHtPd3CP9RfB7LTEaCo8ZO3FkfHD32RB
vfDhWLLbClVZUY+a5+WbLiOK0T4MWzXiMEYP42ccRsHM6Z4tzgT9dxa+YHbKor3N
ntReRR6+AUiIttKy6BKSGUgvYrtV56u73BFzNgBxm+THOWIi/ArwKhrWGCy6vlYS
wrRcCFaMx9ZDOUNwbd9jIk7ob6DBRIyl76xGUqU9Irs/Jm6IS2jjzq3OUPBFDpZb
mqIX/7N2q8Z1s1bmd3tUwQqDkAD3fLP7VMdsP1qwRMDDwVNCwIoqTqowTdzqO1dS
Z0d2N2XVe7YFIRblJqg7+cJWM9lanbiwAFi3EWYqtgRu9E1mUxIRai0+4jqnj388
7CnxMgsw2GuuR77LBesvo4pYUQBegA6SkChru0CV/Xa3YL7d9Y0Ecb7lI8/T3eMW
JWGYxMLXQNIy6xkmqCf+pmi6t4UDL+e4upBTW2Hku6Onskaq7QBQdkfnv101QQpL
AgDkIPDUIvOM09ymdLS5zmibiaT7eXKu18sJGEMzuLXONPY7BT6AsSZXwVvJEZpe
gvdQQv7BITXyX3cefJBFhVQDq79CvyhUHLGUYp6lPfHxkHa702yxY7OWwGSob59D
fIJXFcBS7+LrCM4OWBQJKMJOuXK09v4DdigYHw8SgK6VknlHDY/JOlSJv6Kt4Pkw
p0EZZcFdSaQ+C8VlFfJ2wfJbnyk89NZJI6XdcSNMb1XiT7cbB1PvrT14+3BtP9OD
i5/RJZgj5KdQVQaN47eWMeLnG3wda0Uc1u+VMhh0bFbN71wjS3Ivzr4XuCeRisBr
ij4H2fy9V5j27BnkK4YsDI7w2FjXyXSsHolZx8wQDObtaSGIocHIeYiv+Svfj7mZ
LEgxZEDRrJSC88QcP5+u1+RdHAy5k8QA+b0M5KgKTw0T35JBOunb/xbXhlNYN/nQ
BCG9j7Y/QTM50BK9+g3bpol11dImogP9UqtcEWqMSCU+vH5T5Z4Jkkbom6w0yq4e
uB1EgqfMYVwTAgLzbGBewbfQiYca66d3LRbP8ts8y/RBNnqUK8VOiUUNW9KQKymA
DUMTrbwrfjvN9GFd6xEB8Pkq2v/bou+/GY1jLolCv4DcdEEzUmwkgY0U56mSeGMl
6JTwMioN6dzLy5tVVO1in+W8PtxwzoJQ39334V0SLd8w//YmgI3rQxlJEJN8b1WE
eVFrsUvGVSCRLo4lO/2dFX7Cu5w2jJOo8qQuHFKDMW6IyhRwwK0GTQEGOmdPfI4B
doS5q5H4X6x1H7KCZKANW/DPvFBBPCy3MgsLyYFau26VJtpdES0ywZ7n+sPyVGcE
xBs0pCnf9ogeTCg8QT7fZOoGlg53rMqZak1jQv4NK+79uGioPvpOwT0xxn0Iq5/a
AK2ylzEd4ZOSkfUWZqWlPFUvpqabi2UF6r+AtCYMEg2dCg0Y4yiuIf+nhFLDrWsa
07IVvXh6HtXb3qj9TMou3Z3BJfia8G8+qUoZSc7BIpaY0F9Yb/lZoiLkIr8OOGcL
gbCHKfdJQcHH+utu/HqKWdpsgNVK0YU8wJQRsSVQh1j1aZ23HggP8BlehimSF+I1
WT4n9rucB9tzMXnAKyhHOMpDuyNGkw2W8V0873dlCH4WFIHG+InPhgRsb/eLUPXO
rYQBK5IyJ12rLEz5uVSeQnpsU1RERFPqzbzU7gBVMHq23OnzZNPRMls/6oQyo/Xw
ZCp3vyNQHATk3rNyUVk8h4qvihbMZKGs59Sa3Ulu39ZXE418CC5JfKIAEybEU2ng
VM5m4OqF6u3JmA4shypgycgQnxfyHHwsYHCA1LZ94aBRzGQbQjJX2zGZuMemcDO+
jykpb7WZMaiKh3hbvlvJsxVRUj0JigMoWToqR7dxMCZf/N5m6PzP57oI93nUnkR6
A7oWyN8SldeyRpyjfmWAKSiqfy+54SmP7CigS0jVvELzNEcInB+O+hYtn/VQ80OA
Ubhla6x5IjhgiJSVe9qtzAfzpT+Sm3CerXmoarPfsmFgwlyyTbxMKVBytNBroLU2
L9Pb6gSN/Xk3rgGn74NiRT9a7Gs1oYDkS5rch43Vw27XZ7Ejjz2LWhrroPKeUdsf
FdRNu73hYXG4A0Oy9Em5U+/6OwWN0+tCRgzNV0T7AJBNWi/o9pP1EKYCvHHNV8RZ
okJvS1qZ5pGoeSHo0j4LMBAU7B0oAxiH1CMGUzsq8iDwP/grpSc4gvb2yippp44u
k8XXboVl5HHrMpJgJRm7IW5Uz1cCpe670vw4ugrqjFtpxx/oRyzQdR/l3iVIVXAN
S4eioVQTk2MUJzy4CQbJgVA37+iteZTvvfG2sgv7MnKsAnuhYRzX4tO6oQWA/5Yv
3cu1R7yJ2af4kvA6Pehk9TwdZCKALiDN5m9dGjrdOKswl6RGZHGQcX6Ha5I2MLQy
qYOIUUBJNsWS2L/5S8iGx8nacsY5D8iwJxiIl7x+BlJkBsuzqIdrEuLrWfEUYhtj
AoQVpgqwwGtQH/5gLak6qUARji4O6RjOeba3tGXGEQEpqRfZb+B9m9sC4K9I4m1G
7o5VcjrezXM76VoLKNaL9lhdofLvprgTFK4Gdv61UVL72pQF9fvFHbc4aKfc+50M
pWdg/LAiSVRdbK+57Jqs3HGm/FWtk2he9dj0OBJV+qgK19iN6A1eKpHRuiYIzPAt
QEqoAc2kdNdqIOSvh7I77TDYSyhdZ25cMHMQFFDXIxhQXpTwmGcb+aJtBghp5EVC
WtqAjrMlR2zWa7WGXiZpumaxcwyrfGbD8M+Fo2FHdkHJEbtzBcGobc9P+D2yjZ8p
RT8oC8+wqrXR1r2SGhhwaTCVIlHW5nBvnXFrcW9cF6uoxeEifT1B6nxW9ZTMQ4sN
srclI9bw101gsdKWrhJJHq6e9RU4vFMyXjzkcbCM7vgFwnU4gu5am61xN1sBR4S1
bBCQan9SBrcMJhSRWDlNr6nBeSRSaUn68eM4TWgXSOTqeb7bxHrbI1Q9+8KPW1SX
p6zeK2J8CKGGmpRQ863IbR9dMaLugCE9P2Da+3+i2qp7Xy1Qt//LcfDd6JA7pL0i
4Mk+WJ6OSyo8t4yfKKE1cXwG6XhuQCebtrTFgZj0ft30v1Ccm5FatqlBHj0gB6XS
x+bNFQNcoCTWbFGpvOdRa38XGc6gjtxm1sy+I99LhmrLwPWN+rCXjnBvIHyDzIwp
hT1+HsJjw2YUOwfBDYTtbU4cABYPgXYfX98S7lx4n4od7KfJK0VaoefPAJBsLTSG
E61CJqgh4n10G9uqsZRbGOQmqPZi3y7Xk3b7L+tPlzC/IMO8JJSnQWHzFiF7e3EF
Z8rxE7m0oYLjG1bIXFSHQz+qyzL5Qlrr4ewZIM2HphlS1TF6zCUdatWRLqsT5JWC
CKyL0PtN5baO3vFFzxpZC9AxaRXcRcj941Sc8Hopn4Jd8XseBY0ZO9MUb5/Pjccn
hJeAe2vtnIwBFdCvgrl5aIjwXK0eBlAD5okXHt+5CULE5RY3FsNOjEbDWgcH246n
Xu+UCDmh49BgG2PzdrMdwW4M+jvJZLxF7uTAtLjSZCbv4W0dLy/SppwaKgi0wV54
tcZG/loihHv8CfeMgIFODb0mnyhhsomvd0CONXmZ0isZwyf/IyAApjT8UTNMz/We
29I4c9F0cEZVvIEs9pva0ODrdSkAopbBTAB9Y1NYaW9ur1L85izRKrULyFxdq6Gt
iuh9e5g+2y+1AK5+UNYkqkU+vD04bagnmh4uvhxi6GiDohd7sawfzVUt48KVQdXV
KSIcmXqPRRvHnEja+BiDtforA0C1eMyS3YXlO/5PJ1Ex59t/t7UXE1FudCftf0hs
uw0b+hup1RHP5ak3Q1IxF6uJYSnWGT1TKrvbb7/83Y1ye5o6LBjPpCsSfyFY20K7
/hFA+VbkZg0WzSqs2PWA4fhfw/tLYJ4N2jmECbIO7kCUVGKYx6Sv4PFR8juME2mT
mzAqzs3qZVYogmSqavr+Kt4D69SBZDzZO58m6JD3jvl4E1KUu2o9xgI3t4peBGB3
BHUY8+sSvr+CLGRWqQCirpDj5ynqpf1yn2N5kz8RjGq4iVSU+dVDzUNxKm4tQKef
Ei/b58kYCFZoTmB6bycpdx0A/QT+3pxhRNRDF9aoVtGPt2n8a4mwvpNs4PFAw8Ew
zf408u2TJ+t+ZOFj8VCKpGzYNoza4/kJ6K4age9mFZyrJD8Eif0ZydvQdzkfTf8A
EoUCVK5/gPTo9jyOnqBC2X3FfCNhcxkVBtUA2t3ME4mr3w6ajJYc6tE93+wJS9O1
iCEa4HAA8rtnlgs2Csw5iRkEWgmd2L4qU5hUzuCoXEnCcB9hDHJblvPOCdcytBSg
9hB/Eh+7uz0USEiWdC9r88lfhlAiahFqz2mSEg9ZAmTTU03WF8si5Y6UP28A685o
hGEharm/nCNnOevg6tT+rwWnac9pWrz+WHQZPiTpsRZsVbKjn6jU3oik0Fubsv/t
P+IsHoREGuPv6yKixPd2NZz4eg7WTu4RBAlnhwAj778wnMYhoqkvTDLX7XPGxxdS
ZVeBk04GZHRpp1Y0M9UC+t5TCwPkKqQ4wDU/yQLTiijDIbxsdgGY9hYNuTB18h00
/yRboY+Gy/1Rz/HHKCVg/skj3t4/v0t6Yg9kbVwUht8uPTxwWC9QF3m8U+u7clUV
FTMLCISb3yn/1fZdNaRfWR4DlQFkyDXKr7FhkqoX/zRr5BoWRGivIrfjRx139qTp
R39BmQ62ZlyUngqaX2DYrie1FBuWvkT9IbVKvprMkSMpgd+U/ZA/w0LLuZ1iN5vP
Y/9cMTSF3pKeXUErSxgDFTQOCyZfAV4Gj9f1UZwbZ3ZPNuyUQ5UAvur56Gk6Hfn3
MmjWdI7QQUC6TWW/tshLbU81p86oxQrF6mcetKjK9yDATbxx3xbQRoSbhYwO7n9s
sN3vXlV0ox9jUecSBp5XmNNJgD4rB5V5eTEihV9Q9R2n78UMKN8N7yMn6pcecI7z
ixSM7thytCIiIb0sWt96UNuXU203HtufaqOqPvIOYQ7OG51BuL5VQ3fC9dyUvbJp
PjUXcPSdaPBwFsug7sLN+9NwVgONcqFkehJEqpmMW/rjoQPz8pODPQV9NfPh2phg
bwZp70uekV9HAyN9rTeiQ0RghYcKgGEZ+RivQuDWLNAP0BtrD93+JcViSzTWg4Qn
axFH8+xOoihOFaA4ZCNxBwrMJwgNi8TXrjrUz3tr2EtUX4Uypv8VUCeES4bnwV+q
PHgBISJ667PX7Iwn2yRx3owCkxVWom2gg/y9Q1dvCDwAe9+fnSgEqbC/E4qW2csv
KAvihzSqqWA4eVNAU63u1ITfNXMnoJ9LK1MHE3+RK3J0dGgp4YUzce0ElNzF+Yk6
1Sg0Y+KEcK2NP8m9oGx3WiM23pzTCU1RBCDb4L/iH2FoQDATaqNrycUm0V0g/xrg
3DlRSA3n1e3KRTTcqNmqv3cDouNUHBPOSdOLK9n4F7U7f3cLsc2iJsJZwms6Uzi7
Tfllq3esEAYk50MSUnR+RB0MJOTJV82kFzCQsB2bwCnZGQumrFURuAHaChpuJ4YX
vBY3x1SrzQnd2Fl7jgWBIcY5uEAZ9CtZly0o9OoWpEMtkF9GIrnegEwW0sl0A3fL
MSU/nXwnCnkbm6BhqFwp+tgwtmC57aU5A6U13+We7SHViv/7N6jKFo5tuumhtnPG
IFfC0I5HFcvf8Jv9VSfYFfS1ZZ4OSDjwWTLMCFYVIKRHN0Z4KO69HTmojUNwIE/V
7ES6uMom1LgInEZvxhn7YAvNHhX7IJdtcPPthoJBeXSFtzY6KtToTpAIJYZIkPAo
rjUCdTc7U68So76OcGrwFZIBa4ZYT5DMtqXa6Ky/96SINI+t0d4ClQy6W1qRlnCI
rux9WAjR3nADZ1MOr+r3ABDOuPmf89dcZLaJXQigowRHGukbgM14ws9xtrVGbolG
4TCOOEmCszmaGTtT8Js7nrtj72Jv60guqeXwoLt3zY+LWDIM7NX1W9qq2ALOnLC8
70u1RLODUv0ESrpJkoVcQnSdaHj9MTEOoKB79MDktPN/Jc4CiSSikkILa4PD5RCc
vTJAgY14eXb990T0f3Ql2nc4YCzFGgVfPzAeR0KNZhdCoJmzJqZIBQ/zIWM2EWWZ
+GJmbrbV1xOtujrxXp17b6LP3hHzFl9UYVhvuetTj8vMz/22Gz6Pw+jyS/drkHMj
ai6wvm/ChOKTlLVd54k6o2/kjVR/tZUjXoXe9tkPRDVwly3TRHKpVI/lV0Hkusnh
+fji4Mv2eWotRtfjRRc62hrdHZYJSWioltnoAjgfW0D/C7tz96fiT6Iwq1n/Z1wO
BQDLqpRy3p79E34MNeN3FoLGmot//ufkYwvrFNNjdTWjVVNipE+39JADpgndiO5t
H75wsoKg3O9400GzyXjciRJXktlMitXYCnTFsew7tYyUYxtHKryEWcJ8vvdyRgj8
1dv444cdmqn56l+SoN5L6uKLiA155bMUTqDRGie9C0KFLBIDUIHlACDOefMiTGTB
OkHYS78B35LXGNaQycVUVYUZ8JN74saS7tiw8iBsykBlSdHJysE98b0uY8CHCzXh
dfb4Wx+PwsRhq2shbJ5HKUouJYDewJmv5/bYSpRitVzYl78fHBYnkuiu6vVq/UOu
HkjE3Q8c3iGYhA8lsKd2VVCJ6DUb8I85ymrheLX2eA7jj0+9gQG8RqRJ+gbIFugS
FTt3iY/col7P5HUZ2DWt8CKR6zxEgAD43XycMxDjb/3KuBGNZogAQmbT8sw4z7wZ
DEy9Bx63htPNGvMuYOT+5lNMyohDipVpZbYXeEOfdpeGBU1LyBmg7TvMf+4Zf9P5
hqMfAKWqDCalSbjxcQIxeRuAElMQFQEC6zuP3lLdgFufKm1qMPSWzT6ew+hJnizU
omMh7l8uhM9+UWwC/ZP/Uxwop48mHef76xTJaRWtuDTOSyU/33YdsL71IWJ1EKLm
n0WyxAff6ORyFhX8gwbBZhayFEG6Oxxyqq1GBZPrg/k4V6Q3NQfrvI6AHypeMsmk
xoRtFaX0/vdURVNrcrOJqRxaW422a3tYskUyyrrIFWqkW7ZW7s/Vfj+1Corlu9Bi
hz4xWphV+OpnczZzc55XR132v+IrPVPMLttKT9qsvDeLe+p38ncvqEq+5MtHRB6E
mowHcrzweOSMWnXkoeAaxHam8W932CpxhCn1qoDOOVNXuqeONwtseOlPuEcMKTBZ
25TNenGF2ap7IE8b2SAqvgh3tgPevDAELaSks7qDf0S2ZJdV7F/Gnk8Mlm0RWqeF
bE0XyA28Ylebub6QVXCqOWzEXe4teAnxtCjmW4lW6xp3ab6ggMuxNu7xZ2BOOXAL
Lg785AhrU+91GQAXoHIIfWo2mbZf04BCGuH+mBqDfejLl/lIYmWxoFLcrklNgBbK
HYYKFWqQ8xG0jpyyUmAyNakbdRJw5EoQgadxoGJpyTkXjodo1DUkui9IAzkEosht
CRiCFmKZ5LEnC8VlFzOOgFHsCgs6AkmXAvj9tE22ZLHlPG2FWSC2hfo3/6kxsuNt
wGq/jfHSnH3hHAIT0jgifZ21hfoSzjCNeIME0EfIF9tbt2jNWhOmGq7E6roxW0gY
XCegpEc0rbz2ktZ0zdMfvMPGNi3uBfx00p2yg2OQFgG5OC+OlBa2WwD3tdMXFFUx
XXAMzAjCnUXlTDTlSFz3AafquOJ2zOur9V+7cujPlLEtV/811UVkIbdM+piU0pma
cmmNqDgkb7yp+Yo32PF1UVAqoVVtVrk2OE1CK06G8g1jSguY59PW/yLXlgJYxAVq
s2VWy7nVZN3yJBGmddkwdz+eJjsLeVZ/OD4w3irhFIVAW7HE2P29b0I5jtyYcCs7
LkemMp2oS3TYqq3i4oulzH28NciAEJJzKGP8sS0DVgf490sd3duxspvdWg4VpyQY
IbyUv2ia9yuKN4QjASA+4g28WekSyFKwNuysfeQVFBNjP35sP6WxTzBL4I7YVbhX
l1JbMXEM1Nd1pG26gZWhLx+XpL+T9VhyRU+kNq05fXgql8uIYs5flRu7NeQm7Xbv
WoscYcwAi5wG/M9NiH0B5AU5k+8LbZEFjgcX8gwlL90f0lilFQl5fF89HleX1ZLO
Rnq+YcVfvHQb9WzMMe5oqFPEKuHf6lJnRiMUKVg3vArm77Ulf7t64j/EQZYziw5i
7O+UJ25QdMsspJm84Q4Ou1WaALZnm51ooQ6yDGKNQzz/lnVz+9/7ZGYVKX/IO0wB
DAAX4BGUEvyMbcXHFwllFqY4nfUpJtS3TxwD4pTgJPw1bY4w2evO749CMybqUyo3
aBUdMR/cfWfq61FOnD6BY8U2BtL0arcxkMmI9RjlkEmAc5FXPPv9Goe1pvNyLoWG
bB1j5JoHppP1hdD2vQoQlnYgyqWL1KxVa4DlxywJVVfPpw4tPYZDUg04H74i5iEw
aODOpVqafMAvgK2COaBJWvzNLbI1rSWTpZn3QRSpIJLIqbj9/lNGMyROSAA1WVtv
KdqXedrSNs5fImVtQGs2/Y0lpNarv/Yihgd7phmUHuceC/JssUOMOm2fE7IASPig
x0GeKV4hYOFTohxkgHCLUEppMhyByL19tHv5C16wVS/cD+wN9kgEYv42tGUrMflb
ufA6irAw54iCotcafGmqfIZJVN9cjJH1HaNQ2N1D2rY5kwf0rPHevBSW+zgSWoMd
BQoJFHRiTomA62yX7l8rjHO9BHG7ng8Mp8LaVo20su81in66nwHWoMnNODrLZNBz
y0CjyphuXG1LLas9ZQJdf8zU5D6pVluKCnoipaMRYBYHVeqY7rQYTaMTDnYGOVFy
Ez4uy2rbdyuj5EwQnhTa1LbhipD0uE5nZup6hQYjzWyGqOI1Pd1EtWYST0nCLRFx
RqBwBXeFnmTZAQ1KlLQlSufRXV38DnVV+8zFT2UActDfNQOsQt9V906Tu8oQLakM
DVx7uQGWB0IwQHL9q3OtyuvUtEzSnmnhRdi8OP9cHqOqrF0Jdokg48QaIvDOk1X9
F71XUQYGGjk85IMaRSaArThq406EKzRWH/QB4q84Qw5bXrswnQ+8updjyXfK6+Bb
9GwrQCA3KhUsDTRO73x0O35ksozzzE2socjitCOgBz9D2fpt2IosPNp0WLm36z9w
q9ydI6V6hIFDxhdyKsdZtXiaQknwxIe7LI8cZVqHMqOQ51xY2JP/3C5hBmSbT2AF
3k9pcvj/lQLSbHn/AjCq3aAhdMRkzSDXbxBTRxiAZi5GHb37hokYHy/bwaDVir3R
YHZYPxcTcErowzXI6LB002ZZ+dTccqKg9977OV+YxMMCslsFPGeobrpgvJceUemx
D9dmV2NxUrqsgY9BQm1hg+kzxpQHVMwaGE0Kw6RpguYBaGGjSsHe7INlaHDLIg1q
BcSI/Cqrn9g3u6Hga0Y33tQi6p3YiudCEST450+/0OwTKjZ6KK4Lndokh544U23M
Skd/mh9k7fzKkh2wc6qFXCWgWNHzAG2JGXXVwya0Gzb+tGOMFHayOzF855AD0oH/
0O9ynLFvSN5YIcuYMySCPq155kPmHbfxOKbOCiLe7yFvCJssG4VMBMsXRbrnPqot
t24lHoWA0kgP5MsTOi/oO+x1PGuFseml4THCKaT2BSx1UxsDTNqY+3NwAxWkzBXq
UbC1r4cB+xLVEcvE00zJtclgZAPFKSRy7OK857j0LWBivdk8ov50I6q9xJO1ey6j
nmkCE+yEZrZ2IhyJxjXrgeJR9IhbgEEK9T4VWmXLEL1RQjAmQAXrOlK8kygGywl2
SMCbh8rak96ecSx8YcysnTkCI/SR0AWWUlEzlLn2lFPTKHbPmeeisx5DtOs33VEX
aU280oXSvUlRrO550Fdz8UkHwrQQzEgHBzYMtlBcVQsq0vpRH8BOy2xgFN5sf4Oh
Db1Aa1azihcYGR2RjCQUj7j4PLIaBi13HLZOcFaWzTOEGKaIXYxhCJs9slmj9g7y
e2VdvBld8VLhfehr/SYGGirluYSMTI4dgLaMzSHq5c3Sh/UN8scvirUPUwvP9X3j
UfJ6wh18sk+mMGYqainVEFwmqFjT+S38SNSx3uYPXIrxlr9zm9Al96YETd56HSsj
znm8xG83MXu+B5SMPTIPxsZ9VGzgycJQOwab1GIybMS+9v2Ho7N/0yVIWLQfD15J
iNDVLMZ2xvJki5dKh+TCtR7QjBdcfDEWlsqXQVxF+CaZ4faHZiETUSno3FOIHL+d
RQz7W5+PhcfT8XkkBazINSNnwHY7HYpxQGI5xM++KSEJxkVdFJFZPgE8JeBmPfff
8TrQ7dKAArmp/Ulwk5nkV7JJlso628waMiQG5SUnoAwa/xvOvdBatFuw79Cth44S
ySlsudI7vPf50AG8Hg5KL9jGjJvU61bOxssGwRevx+2jZAJ6saJl96U3RFr0ekB3
0QFLeHN/OOec36ROAfxps4A9bD6ykMpJv1pMnf+GYhimTR8mFFG3sKI7c/+oDXCB
gPKgkUqjZSjd4s3baTLYoOHP9ieIvWT3B4vmWGi6cLiet3fGBu7tTqcRIOmh2EWe
wolLLIhb/+l/jIfULvsB0g1C0IIWZDSN+sXSTCSRB2yzcbQyFUNUgcHcg432QdpQ
I+JCEhD+pTPjNAkHa6+QvFAtv0x0trLpxSKcuL3lz43vikEqoIRa/2TRU6gNMOhj
HOZ6fKrKSvptHLb/RLaDfmjcQYbBAa4BdKR7b6ZXy3Y9ffsn7d8T9Prft9jCLHbG
GJN1hbWE4/RzI2Gmy+lgdkP2eWiJafd5wPH5VtC1PdM6tjkOfym5iN5lcxd3zQ87
DhCRugdv+KMdiz5LwvgejTXfGsGYayLA7nzUsKlfuE4LqYDH5pwNlGSrsk0izyqf
Kp3/M1hJ3wCb7xGT+DF0zYAcgFBkJpuxb4YoQIuJs4SDe/9Dxq4ux9yl8gmj3FA6
OTjPxBKVBL1b3XddWZ6lszVm/Qe3Dk0Cgt2b/zEMIA4vEkqVmPFfV647zn1dN8RZ
ejqQ2uU5N3IjWxRwQn++EODADxy5vCARHraVW81NI7v+zkVt76Kf9QovW80D4KO1
o71TH350+nQDh0g2pFSYkz0i8uZJx2bH3DLNqGYE+L3T16uOBZy2KvSSB7+A5Fbc
L9c9hre/ZQbiniyy9qr6PCiTHiu/Be9oQ7FDCSfG7+Q+m7VfUrxc/AS5waiWzVMG
VfykJuNQy/L2zrVGjGuViidEMSGT8RncU5pPooX8GUlRvBo8fwBY7YSsfXSsfiD3
zWr3EKzZvkNuqua+C7xpG0TdylRpvP9Z/88klnXoqqp6D8IYmHV9bBMy9dNDXuh/
VNo/1CCJlXRlQSJMDNEdPdkgYzATvQ3rLGwOA1iTxPsQWAVE1I7wMx+gkpIy9Mo4
5wLE7xG8XR1bEamhOdsmxnTVDVsTN1hx52mH2/DerxserYxEouTcvmlkSomYWcoE
zfk+4XwXS0LrtRfOJpVuFDG71lSOWu0IPQx6DuCtwLUyUYzZ4XspQEREf9O7TpW5
rCk8FQfmNPVEEyBUlekPZEUR/uBNdNJPVDlol2w0OJic2jws12sVNO1CyPMOiTck
tXWK05K8Pridb8OBKOPzxqoRYWswCi9UTS5oPEqcIHlcxIrdVgANK1WdYaCELehb
pzqRIwokt7QJeOfM4SwM+/pmct3uE999iKcDOD0lzOMUuMTGUpqx6C8BdoOAPzF+
DbsGwNCWGw+RR/jO7hhD8un9d7ZKzJAoabT7O7RYdFC1HzGoi3g/Lj4Vr9wYespR
AnBBJtVSJyIiKHcTizxcVgq0aH5tZqR/1HAPnaafpoa1pFWvJF+UG46OdiltcYdF
4g66sb401O5ZqZ8mlK2jrpA6D3Ds3H0bVL+swtqZt7GTsYajE++/rRhpMGmDKDNO
Mc4vCv9O/nqtU6aOwXywe9Njfr72hv/HHyJ1/TZAMVfRFnevT7zWJzpajFBaZWCg
BnCn164hgpW/YqpIyEgUWjcjx08BHdelzp7VbLUZKn3cc6ETs06qC6p48ng9TRyz
WvK4E5+Qb0L4lWoC6qJptO064awgs5C5NNGPw5lrCYPl83wgLtXKkHQ9+P/G9rUN
oGv/rldNgik9h18KlsZbbg6cEYFXRbwvbT6UQI7a+PEbjlYEN8EN2Vu76Cvprk6K
mnzaZpnetLi+ivoULrNb/w534PW+rhS0IXfmtRKMn/9d24FG7zNRHEsSR4LT4hr9
YRF7X/WYBn7yhEvZHXAzhlWAjUWd3ry46DS1eJiRucjc0KqblplVdwVEmNgzax6w
IeLPSynRq28xwQqbxn0sO7uBtsjHoBbah1kg3Tq0hyFLBKviQai0mWUc4T0Rwedj
5ssHYHsSgiPomyYyJ/peNtdHXjeqCr+lzOStTxo5JmUGE7jwXskhQHv4CF1mfXWA
FCKNWqy0AWC/SXxcZOuaqIEs46wZvanL+4dHAhJUcKy6zJ9+qREB2FcwVBT8sYMn
+jECXEOStYwAAgaZ6hM/s6gQE5UBAGpaEuJz5/RdQ8W0fHBFRddcHwB+I94E6NxE
gkP7KXAwPrkcj9QvXEi9dYv6x/t9u7h3UB65Ae2Q8xki3QTnmOVQkwtVXlWp2Ier
bxvKTT8uoonCanrJp3I0VNhcYcIYUtyEd87UlYeJo53/HSaHUpI0uh1PFTr/hLRM
F6qm3iVsYzDqOP4he5vsZezAbAWFk4U+3H14lDBh+WDfm6HRFQ3ep3d4Qjx/dkDf
a4+udjKmYM3X70ED1WD2cg/VzxmqDNh31G2JRzUqgxOIiVP5V3tQRDpyHe+xIQ38
Zf2y8Gv6eABQagCT5MPhekxgJ7jfG+cDIBuPuZXoRmC964zSNiQixDvlz+3vN7Zw
7Xb5GExp/ZmDOirLYAX6fwznwaV54hTrmFCSQw+eQVljS7UFDk5jcT0yVwEeSA7r
Qw65N/jUGx7mLbGIqehJCtbFt6qdKGug6gnSqGqHCoqY0l0Goh5N8u6K6mZu5RmU
0h+ztavQa21iN1S38Ef96FBmFB2HzrXTqYdymOTM9CUuteTEqZLCkOvCotD4m2v7
TE4SU10+qqLiVTVtZ3oKLmsGpvkyz/PwcJuoofA4IMLtK2C96YkqDzx9gw9S27vr
YVz6+Cs14qkvvytqukeGI/7wWiKgBEnTO4Bexj+OHe3Snqwa6BID2uYvgUWNifk8
Zh21tLBMvnzU6ELncvpfCkZgaXjwoShptKK+Q+IpBfFv064wGSwaHY0IIzK9PQ4j
DnH8wekxooi7SX1FW5ESR40c+XW+RmTreALa5M2vTHrMUxbHjXSQ/kEIGjcADH8O
itIsoTnOq2iTsg3G/8vM4L4KNj4fEsplZc9U9H6TlZhCi5hK1xiBOcar5Lf89AHd
2sK3o3ciWI045LLp6XNyVw/B66SRnVtD4JB2SKPLhFxWt8jkxuyt+qc5gRHSN9uO
/D3BePzEyN5hefEkfVvj4Zhv8WAT4fq3btANcqwkCSMtx/7JYnIvG2+VXSUjFTJD
TRjUVhpv5jOqC+a1k7nBvDn+vhWEpVoNjh13WoNDSF3Eq5qQf5T6+lKaY9i63eOq
bNT6zSKdlBc4LYZEPRzkxjCKuIxMWoeU/85GLv1Ovu6K1yJfqVvfqbkneiW8rbEt
U7V5Y8HuEiS8EVA6dH2KRedxRh4qyutZSsgxcdOb5DJPuT9tFKOC6MDJsZe0XdtD
+dB0cYCv0U11tvr5zcyUVnZuNN4KoBOZBKMWge6h8pJSxW2DyKIHfLQU/yWr1y+Q
ItmtvAUbGZ0BCnLgXi3BFFNHvIcGaSXHhzV1BHHVafdDfbhfvjt5XhOqf7LYr9L3
+IfQORAB6qzrgE5NWVld+9pXJVivZsUwOhLz548v69KVr8SpYuF/MeSaneP0JXO+
U1+R24msx5YRVrcN/s3FupqhJOMgBdPTCKuGaslv7AhVNCLVFljf7sQE6iuFd2HQ
lqFFTc+R3MPxXgm2ksVhCjplc9TecPY0OGUhypm5qOFYRxUFdOAMBIA9IzXuXKWs
/Ca4FecaeCgQKZn22eBAMf+ijFTJxZG9aSrLKroRZ+g8wkRAHIJxyOc2Ur8vlNbr
9kXJQ9ffcgJVgUlufqREa92fvBJ4fJcwNhMTMvTNV8nHQA0ZynE2981NIFwXufkU
hCJqEo7KWlXQKe8JbUxAhg9u34/ii5FR41dmqLtay9wX3lTyYd2QqzA9ue6JIYVC
yaQ96KqH96iDRDI6QMKDmxsnCVmo/4AmCCGagOKJ3MgMBwaGUa6r7zIzgNHB4qKs
v8Y+7Qe+GsV3+inNQmEUTRC/ZicclIGv904ANf8Dz/OGtN7hgCVAweuoNj7obWJW
jmRKt7M+9ZlKoRIMwueJ5g0+8Vu2L605AiBpA7HrKbaH+ZcnWFcXYXqp7+w6wGI1
TfdfX22JnQh/qa5dMbDmxad8Hg2cBTxstxdnO2OCJKe0/dxw+SQ2PzuRYWMIAqDW
C2s4BrUupaILZ+6NjwYXEBXAUO0FMrnkGgyqiaGiC+YhZ/wLbOxsS9kJBNwkfqMA
DScAH3Fs4LooKxg9vrrcDsXSqPjAAIZc9lMWjVu0ze++hPsuB27J6iU5ABRc1qmE
tIrHfZrVnin+ushxK2GRI3v8bKXO6bho1AmJBPeBXez8qAQJ7zts3eYyGNy6IUcC
S5oAyeSMLipB3L9cJFIALYuS3XaDNw1IsqqZZOayY302PSOXHPMtzmITtTApJIU1
luFhEcOlb5shghCu1YS6zyIHvZkP09WMdtWGjXdb3a74zpCkTGjTsX5rufPWlYRP
zQBEhz4c0L+fIovqFpYVApl/Ldc3OdtkkibZj75DtIKzs8EbwGTkRbXgH9Ms3P0i
RxxRk1RKlpTxehBahrEY98c8cQyf3XzHyyxwfy5PEjaRalRHghjbX/BafsDYc+n/
zPVT8J5bGBaQo4gDDohzNwrDGjjtgW4qRghHdMn8STjvuO+PddNU4GrDulHVfRaz
HonKjZn1ch/HR8Lb0240/dgncw+ihjYgtiPU2kuwHsm0rBACOPyaAEehEl44p3Vw
KOuV03m4lKnjP2OUKxBU7BLwtAwBT5GhxU4+Ze2dp5GB6i1K620GTkRP3zjUrcNC
pE7/R/HYXX8RwbJbPnVogm1oG5WZ5P9APdndBxRtByosOrAgETxJkfZ7lkGNjpBo
RIhM+KBqiKEcZ4eRIl6C0rMlbNVa6jCG5tKpecFrpeaIcIFKZnybyv/8ZDNRsrpt
fUL6/9k6kHwcLTaOV3bnMwzAmVqk9NrO+HxjFTcAyVtQ6PtBv/OOsNhQRN9u1Qjb
RfxbmbDxDcmG6R7bOqBPUu2Rpt9EKvvRYcJ/Kg6kZje/mCWeMtxONvOj9UbV/r/O
ssBbP42GDNlpzweAvM0oXuL9UulCTnJTRSlyO2AfwQkQGRYKFx1N6ZTFyrpH6iP3
dD0ugsDpJ7PZXukSiZfJ7iTzicWeBqWFnJEc7fatSNDAoTA3G+FSYqvTJkotR6d3
P0TpiyswPxG77pPu5CW2X14Ru8SbMKhPk/ZrhEN7xYRMFxi+KH/S61+UY7VcB5r2
exw0AQA9E6vu27hHRElCKUHCwB9XxpJ5ke2wKOISrg5x9WVSGu9Lmwaf1TR39OrV
5iGWae3IxqgEZqq3IdRF6IxBqOLAGVYkkfusv7VTgAYV1gFjrLS9dQycESv05zj8
WKYNuii0Ygd1YCYUCLy9LQ+KJkKEYs50aWUxb2DVOyisVWHBkTHELx6C/TwyXuSy
qaSAY4SxYgfBQ5qim2eVbPSGcRAt/J2dy0peAqjDqlXMHra/SZg5NztWoPr36t4b
xSKJV1+sJGMg9OEH19UIX+Yke1XcGNvoNqLUKzQxFcM23vA1Blc95EUsDZI+T7cF
VXhHNNeKByhdoqGA7K0e98RumOps3Eoeccw5FxYvQaOau5NVogHvpOdVt/k+sL8U
v377gOEMVj3oW8glnK1ZTbN+eGmRHi7txjPS3SbgEJsrVLKevH6NIZhWdPzNIoI5
pGtILmva6PesKE05w6GQpseMRBEU3LhEjacYBS8M7hIQlzRejn1Yy/J8oCwQeeCt
gk3YYqED0hl9ja6wZjExetkL1YgKPQE+n9rwtevHRoM6br4TUmzAKy7JlKMEOJJb
xkKkQBwm2Ld/LznK8jNHl7k8NDkFqId8QCR8CuMIvyRLoN2SSb8o5GUy74n0FL1K
d1jhSuRWBkmaaLOtif+2D7JDgoe7Awzsd42Q7z0Fb3pdS12AaDLlBA9PCZNgumbf
T+mtHu0UG7MhA/KPAUrCMmRHxuwLy4XpV1ZoQf+tKhMNmE2ipQZ2h6lyiGqTDDgQ
BnAHFV1PdXtJujcRUDW4C8M1a+1kjk08ssDXQkvo479U0772Jppk506idGbVNfSQ
1gjJX4jyJqCZ7haRUvonRpvRI0J/r37ie2fC8Amw3qUISe5DLGqd1jwWeSvA/Fg/
4DLSOaLa/TKoewQHdlxPj2em6GSCGHXDe5PWYvEaFvkhTjYrhBf//MBrC+gYhhsw
68Xy/Nvsz5rVnJZYEhgJbE3sGVSX15kxXvzSwoc5K/q3K7ktfMfaEPbeaGzM4I4Y
JnPwYF8G5Drs+oxJs7Yavh+Ey5KoJ3mE537huWWu05qEWHT9xOs4PIhcFvURlHO4
7xaL6r+IBk+A8k4ncI4DJTRYi1DFYQGe/6OnSQktULiwJToQhn5g8u/v9+39dlYr
HgTPI63Dmzg5C6vUieCbBWbO/WmzgKGYYrVh2vKfMoVB0ZBccr4ewmA5QOjmBzNn
hAVNfUDVxTWdkw6pFVT9DKZdNKebShu27KP0JvyPTri0aZpgNgOAqobnz7l60Wnv
xO9thzjZaioP0aVdprEgARSVkPRKTS5dbaqmcbRgLQ565jkxbYBCraJI7KAZRkPx
373HIc7hGHMBc39QkFYJ5tnrwklVhk2sujCyhQxjcYNhGLmysQXVxZG+o1NobzZO
I78hZuVS7APxwTiIctdDbP2PMVtdx3ol+2HJ147Rvk/snR9IaoDxjXcIJQ2pzsS3
WbAJOzLLSgxhs2uk/smmupV8qnG3KQHSitPZHlrY/lFcNgZaemhhtNjF/WmfGRb9
n0wMV0CIhkc9CoO2v1mAM9CxwGxLjNb9fzpB+fVLz4yn9Z2yBGyZxl9sUgGAt/19
CMRZ7BWt0idCUVP+sBJlHaKqjn64B4Gimj3JRXqtRBAvaXuCE1ZdGlBJ1mVlkTjB
nzT4YEPRKazD6mgpKK/Q7Q8RBZXtKu3ZAsGSjziQB0qjGXF11O8B1DluEhjC4/ea
YX4l+e4k54PEWIkU5NuRv04kcXRrjS3wG6GW5WbQNCiMRD264O3Pi+cSzC3oDAPv
nkTG6TaoRHJmndIvzhu6RIm31ndj4vzcG5o2eTTbozLEz6mbFPVZZRz01v0cvFEN
l0pqB7/4/qvguX9doQ0W7LBmXSDKAdHxoPSQuSrT9qN1jMVIa/FwCpmu654Russ7
oYAISTk36p9nXRceVzWD+x4+unQGknVIxzMxKXPOVenqP0Xqj/IUOr31p00wzY1g
1M8zgsnDlG8Sn2/l1O/L2D5s1cYDOLvh501ILQi0Ulp8HIZTRfHqGE/jhxLgtdTD
KRaT7OXgCgyEbfa6GMOn7dT20yaKWxJsgAJDC6Tyz8OaqMNx+1550nIZoVpuqSWR
Ji/ya+JL1IV+Cg4a81VDw2oWicVUSpiCawaLRfg62J5iPEX8EjwzqlWe8UcFUdel
D5QwfSM04AkXA2fdLwM9uoxWPZJEdOO+PKfh8Tcf4lJljvFtkGdQXW+6ouhtrKFQ
3dEjDNDfeOK+9iXRD2bUtp/KkFrBOHeTxhGDCWcYY0T9+PMq1eO69Z4KWV1iPCYI
QdeeFi34LBBhSN3Q/zBICai5vhXt08IoNW6GSgBz8xttRR/0MVMPNv7AbIMgWoCz
kHZ9cvssk08P7rNjQGNinMAcs3teKxaZ6BRyig2dKdB/Ta0pWClCQuo2vLHoO4j1
NtZYgA5L9izvgMe0z19ZV15kE1cUg2tgbB3bcDRDnDdxW36lVFo4I1LBLWF4Bkv0
mkDfJ92QWPBIiBnbg8JjKmHuzseaUxfCq+u6pnw6hjSKbyWYFmXVZP8ORZwbxKh6
070hcvvAiujeo+gsmWhJx2jFDRjTA9u5pon2tzwid4ziSFMdncDNeVYDVVtSMQrc
tYcjWUyUMnNw6CnR2V3REthT31pRWN5XC1zzc35h2E58dAeXdBtPiJioZGLY98yv
xUh2kzrkHB2o4fMHZGcneiDb3NDDwZgIDHKij5TNJSFqgKtz6RsnbD3iZRdzwGh2
7jWXYfZDN3nsqhSA10gx6VpFpmlsLst89gda+Mg3D07SDvgWZrHTszkTr/ciToWC
Hxq0MMbETOc/gM8zUtIHSv0LkqIQvbrKWdmIdz9jJVncVtSQHCNnObzYaFzs4f0V
H49lyrUGT1yOaK5IiVXFF5eZJEsnFOUra2YJnnxlWfdk/OMf4zul5VIJAXg4P8PL
bXFK/uoBEw2KP6Ka34WbL7Di4a8Xm5P/tGFWNF0lMyWwI4Iht5GpUom1Io8pNegv
688Po/kuVecWYO7/ovJgUoD4YRUZ/ks7a+0gEN3NYKTG599LQt/e8gJ+5D8tPcgO
89a9BAAUWqcbsNuF+bjwxmpqVSZfginO6QczBbH5WRW8bRHZw3rRKmaVzxkLJbVT
GC/grXQYzlUJieiqbmYxjEXQl+sZ4kKY+VBBGTNeLGTNAQnk9lYbNwnhawxYxkjV
9EJ5VGSb7ztmR4WFHb5GGy8FUou0EP6Qootn+tAVzcKEdWvpEOHMcybxPL0Io5xv
kmzNCV9hjROng313m2FWPvcdhoTURbeTr8Z5XlYWWQ78eU9VqN6LQ5zA+wQE1NeK
TBhxAv7ZqXJwpR6VACtkUsbHjNQ0TNBD94Gh7M28UY/qIFJH2Lk/+0we9HtEVo3F
YYKynqSDz2Xa4vgHoOgC0iwTUX0WspoQyLCtlzFiyClcwYKoL20xLZ49VBgN43Mr
EKpqQefv3Hxb1w+bzRezPMc+axScXNeAm3679WuGIgQsXMmaCZPtGadL5uoziAOU
mGJ/DFNuME8UNEjx4YguG7AsUrpsRUHrQs4NptXjKG4DwU0SOf4JcQN4zmZCy7w2
e4Sy2iSCRQ79jp8BC6Jlfb0zy9GITa1BsSxJfdEfgcoLTUawu5STYqCCjGxY4f/R
Wd5wLnz1d2UlH99PkpFTtQlx4w0UpIX8X/q2B4IY7q/G8RCkImAxDGnhkr4GwoRJ
HQ5IHLPoW0Pm3eHp87zUcwERwtMGjhrPL+JY7aP1RGnCpY5aX6a3/JbmtN7lmcta
GOlC522uMgoZ+/ZBwMbC7FLIQWDU2NhjgtjCw/XwiQrEqqz/A5Tp0NfIzOtSg10k
xJKtuBd0ZtLlOcbR6z+Nlf7LFYv0UByZ83CvPsSh7nKWUa5QhuUK9YPhD5n9sAx0
cSFgKd9aLrY9qmNWKpJTU5WdMvui1q/e2cCgc5QgVYnSV+YZ6aK6Tem4w77Zuecf
jVvPpSupEheWYujk8y+yujAnfxDmFg7XVBhMj1qBLfzCpeMgO/sbggRwXdMGFanQ
ywzqUYZVaRUpIkPBaR7sP8rDigigFSZrW3hvWmv8wxYmQ5fOFM7IIFBmcpk+YJk7
6X+GUvTXhW9joyWB9NlGb2fH2lQYEyNdcSlaZxJyJq70BAzCwxU1nsmBC5LJP8Kf
4u2upBcLUxXYCH+hmi/YscfFqN27wBcAZj/mAebeikuVzuAQR2RqHpAQ5Oa9uRDn
xMP6QtimtbIwl+X5m7GO6oBwDGgIai+EP+ML2hYl1AVfFjlk8h9lppm2qWs9xD3L
MTE7VVY04ugy7T5glhstrNMDzAZprr2UU+Wa7Unr11b+EwZfuaTUOQfd5M1Lbir6
zZRcvs+MDYw/90J3qFTcyWC+5L1DnPGvf74AS7UKaKcrJr5pZ9vizVv2ueR/jkve
fNCwlq6NuaCvsLkwqmdE0eReCQAXzJh4P2yZ16yaBPn/HnqsXU1Ixgwdj2Ygqmyf
k6pJesjVx5zrakR0oq6eIIOZlZkZ1W1pb5C/V/ZNTsImkYj/CYmCBTN/GjICJUq8
L/M47mniLznGperShu0yNIYIsjA6sLzFGONn2o1ci7G9gDxHUbRRfi7kyLHHtCJ/
EAHq0OmxExgj9CBHi+Ik9qquWsx+XKHNO/74h1m82WTe1n18Zdo0aVca6LUZ3RbD
gI5PvoYoS0euvw7GbJbZ6d0aJNUlMuChxwuH5JGAhTm8FR3majNeyUrz4YnsDzeB
vBBbNzwi88dMWRm5I7dsDwbdKW4QMRxBz7WF6dh6XX5nslol9Vbe79iWAQ/QntnW
HQ2w66KHiL2feLnVriEaGSQlNAdsdhk18kTD8vz3QRiKVT4wa/ifDPP/yaLTuL88
7wxbP80Bxlr7iOq8GFPALdUlRNac7vi4WyvTDncx08ajytFW2pl/pUfQuwRB7BOr
9igZFzt21wOthOlljpsP7id1iDi4bzHVqIZ4CoyvhaLkdFQFRzbpKpW85CFzylyv
gATNg0q7pHeIhvoxFSUSRtnGyDoY5pm2doy3bPW/uy0zrraqNOkL8IILoXjvACHp
bHuaYgCzk/AHE+xVaTdjlMRUBMbQLVJ5z3xnqNnUi41WwVIjmSvpXLSBHw5RtoM9
4eoFVK9YfZ9CHYoU8dlJBB08CulRF8GilHPnzOU6waGmfjHP63ITkCFOO5/VTOdi
BdeBGVxWgMjTsKrJ9084VmcVUXt34kI+lUdPufUyjpabyt6MGgb2FZxiamvohvXR
+ZfOEoUsfTpi9/94JrImxdGQD+mzjZAyjOK9sR7oyIRCIQK8Le9/s5UGW34POLDv
8MxLh11iLXUzwwc6Z42/ahSJP388d09t/+2SH1HtWObwl10A3+0q9HKFjMh1/NoB
HkQXgA08e49ZmpTo2dpeJSnJzU7LKO4ah16vooMlJ0B9CmHxBfA4ab3X61hiqB2C
F5hEIricpsSRZ8r8CmQoLCEBh15rg08sp743aUrexPu5pYDRBJfxeDi8J/ii5ZXF
scGazfNEkO21D6KK57jOenkzq0uwz9fr5vVlCHGXP8eHDr/ro64/waahJGsO4h9n
tX/TAh8yW/J80E8YhtJd3d38iwB3tp3I7SIWBBaRACdkDf0JjuoD3pTP9ncnQ7o9
sus6wqRjHJAc7iFbWbgVnnliYXYblWniTl1eSsKoTqzQhywbUdF7fxBp8FpWb/jb
ZvEVberEsSVZD1D2Tu+LZQBWMk21GcqLPS4AsDJMMHgaKOxUOhx/S1HeAh9i+P++
7S6rREVWzqmajxF0kJSYqILmFOPd4TnPbpsOteXIFneyKpAVB9V1LzCyu5eTWfdj
43mFXqv3uB35IbUQ6HKxkc2JYX7x7zxHVzhHtdw3HXeFQ4HXL+e6/8NZTv16nOXg
fZ/t3pgR9RJ/Tn9dUiWNDlK3Yyka651HWynGataXVtBvuDoS7+CPmnH5ncu7wWrU
5rH3pCxDdUQoPXZJwE51NV8LvJvvwHe6qczg/4oEGCqiRo3sMfnRK3kMr5I6z5yF
+cII6Ah9w/c7vo6+uB9T3L9fM/yYdTb4xQANL2iIRagdflZVUVsZLJozZNXG7j1X
6dmhIZEPFJFyPeA32nQ4C6K+QNjUv9HyunJRIBjTNs6W0W7A3Z0Ls+7WK6KklqKY
JgMrHdjUGnEm96xAzj7jD9OWD7ph36KaCdFqWa2WRo3/Qm3XeoVMo9jOYTskwCMS
jO7iivHX/9kQOqF5mKR/fEr3ioZPXTc0NwqTgufBZfm28v6zPzNX+sj8Cij/ha7Z
rnrUYMdhpNUbr92H/2WTL3+KZMmlAAWkcuCAnARprqr9dywof0ZzrBpIxz322yHK
kIWAjILgd4sl6pKXgghEGLhcLppicYUlIy9N/vlAEZL1hZNxloS/shbfQjfP0pMM
dkexvYoWqk4WXeqXM+Fh+AChWsMY5Pl/E9uVuZhWYegoVzmdReUOwII3kZErvfMv
qV0vFJhrsHbyY4/t1nElnxgvsaTDord5/b8X6brjs1EdfPR0upNcTScduT4x6jmx
frk3g2N+wFHki6eKkEdiTiIfL62BGYJX6Gkg5xS5XVjyJyTXBT1Z4wxFTOGbgPBg
zWxa2mIbFrEhfw+2yp/SW+1lByzIygAxxU6dCYFflyIj4earjf9FafhmUz7ERA6t
qQAFc/pf79JVIeJE+0fj9cnjqNAe2jnzj9ax51a05QKvm8e/N8E6qAUrlgd8gc2F
53jCcau6HZrbB/6kEhmqO7Ixbi8X1By8Log71yxA6YUAe1IuzlYnQujrR0OVwSek
jqLeeRg6cNHB/AA3rrDuf39eKaQjn8OthxZg1J77PwqUK754Iw8b/pi+BFyTS6R2
LPRguPUKfS4PE4zq09Wy+Qtn7A+q1g4vBREIiwESf9a+bLEx1/J9WxQCCg5ubqwq
3fX1UzvkW4VPN4ju6Ch54G6sDH6GvsZRf7Z0XGHRiDkVHuoqY2rM75gRO0PcrKTN
M6RfQiQgtt9IzO3ohEH49SfBsx6N7wvWsgbxEtS6BvuUeYTdv8g/QfA7GXF/QLW7
ezClkmxyYiLh+8wkj4b7SUadBNi5m+mOMcu92VjsevqEWy5KTtxw/ixKheKhCOgh
v9aBL1s0n2LBlfhBcpqkAVC5D+Cz4JnnFaZFNKrm3JdWnkakmFI7ett6AF19vOvi
Gl8xi1aFZy08e2AOwu1rug8BRvoFow5ql6W+A5rgBqj+NN4jnC/tVXqB3FYRwrhU
MNctGJcep8A7CYjHU1iVZW2ryKBT3PkJmzXfAC9F2/jBqeBtj87nikwPB+Mx7jcS
yzcEJBEihQnwp/dkpaKgF3ScZsA6os4Kme1KVTAKqfzUia5ZJ7xTJeSwTHxC1adG
NZku1sXXr6Y2Vn8C9Xl63DUGiJc+TjkPwCRx/M6bSWIXNjKfwgDXgyuKT68Lgpxw
MMsjA4SOGCKZcCNXiOVpTLCQoXn9aVv3oZiKOj6Y4qwUZlFhwHHSLdmausFAGt6S
EPmYg2jnGnjKbTX15XO67ywdDEOPovGpYIn3XkA477x81IqvIrVPzLR7SP6z3N9i
+vJFH2ozcj/3Q3KIS+a/PkHXsS/AH3xlxsV8/KBVnAlBUL/FBe6vHc+UOCz8ayGE
Q8YfS4t6dGO9bFUX+v0Ql5NnnvpxI/alXig5rrTFIju50DS7RR7FGjRgNBwWvJWr
Cg+QDRC5uofBWHi9SDWLxy3CvYGkvMwD0tY3r20pakn8leUb44UW6UKrq+Gns/Eb
ZdzNU4RI3j92Xt1KqNSN2DHP6GGkyMwkWf0UTmYQtmYTGwaBlb5OWEmolGCmu7B8
LmvB/erwJACLMhgchDrFwnxDzeUTu5n0D2qV3KrGt7ZxCItxPvvJk3Zmmcnn0MJs
gknLsaKEab3UVbI06Twi18couyb65HBIY0U9wQOIg7uVLdQwEPSsrKAwjiathN+0
mFTtaPWwDyRE8mzYKhMtpTikb/9HNU1Djp+0PxXifYfYr+0D5Fjzz0YG7phH0ATw
ljVhIuciWYuBAColmU2OgTqeRFO5H0gZhLFHZx2+gBkddu7jMSaIim9HQF4INyY1
N370nFOrfA0gmnkIOcEFW154Lcl+zj0lFKOP8jU/fJQHiHAeeKlrttcfpvCGurDg
2lq8zgZmikWmq88AnNECCtxY4y81Cg+3E4va3sJdWcfiqGcvbYPhppE3nwOHzlkE
MtVPStzNPEQrIG4ZwKsfL/SuM/fcg25/fh95b7OUo32Dz/gUuhMwH7+xGFS4d16E
wXFmVWBgifH0IXoQSYuOz8ylouGAuVEtSYiyJxtkDXU50IWnvCygfI67+sTESHWq
WaWDStvIwTEP3BUpPDjwzGaLHBxIZ1tw9SwbVJ0CVs/KrIdcVtpzIV9JP1MqLG+2
QsMnOy2D1vZQ0NPktd2cqIdg8kHLIlA8KULUQn5bRZRqzes+IdvTPMTBdWwGcfjA
DE/6Maun6Rmsl12fpG/vNidn/8nuqqlPLQ3O3WKAUcKDYA0y1sNtrCarJoZVY01C
jniij3aXfb23NBfeczzxF7WmSt1DKdWW0vRZRRPHOKjJoAsolzkwsihq2hAocXdi
WxiutgyxkziuQJJahTzt8VJjQ5fFTN5KFHj1btHoXoER2OM0rbsIyw5p+HMI1O9q
X2AKuvsv9eb8eFhyU5H2+3jcu5I9slM1GkeGMbQYD+YZl+cfHJqhr//35QKjFLc6
3GMwDMnmtt2JaVDxzxJ4+rESXfEu7DvHxccQtnoNZCHYiK3DwmC8/o+iwEHmyyX+
vajWc5kUtN47TYmrADYaC9hE6iQFPArafbWDM8GGGD3Z0GNJ32+iaHuNcXae8/I3
DmzRRhyNw0R8JK1uo3ONdtVNwNqXB2SCNQVFcSuZQgqiDpbh66unpZ2EyHn8Wz6r
s6NKnEl4XsFCDNFiYJk972pU6Rc3CTU0CHs+Iv6QFpqNWAWNgShkwX0w16Ame73/
UatqV3ecL8W8FFIDqZPoIRRqPlKnPTwbo98yXfuHWv18WvnZbJzjF9O7PZdP7YSE
6WqbAZuEXcySsf8a3ARAIs3pX45csWbetYYQeyRlFkCm6sPaZbON0p9VbNWpxY56
jUMxCwxAqTPdP12f3/4aQo7BWqXER4EKEEgYfU27e5ftdXSTdoqCeqkbwvFBY1US
wVklVTNYaC8j57gslSgbkXHfmsLXAWax+ZCWI+m+b4mp778X9Za8dXXtwoAL4yC2
rd29t6J9rKPSOSfCrrKqp/xTtZ7fAW8GFVcg3nMSzdwjwp5Ql3FxrWnCkkiNo3h3
xx25MJabocHGzitKGXZztBaSr+WKpQ2l5r8NauUm9FDsWT0kgKj6YYZxk/l/SX2Z
3jwgTA2nmWnc//RiI6r2iImy4CWhjwgEODlumHwljD8hPl18U4WHDqPZM/bCwfxV
oebPSw9HtA+CkD2iGwEflOGj8021GiOCIhW5ig749ozmGDXM52LIdmYrMgrZoPTQ
/K5t49OYf/+hwA6sSvuWgma5FTOTgH3kdVyY755H7vajZm8crUf0zDwFfbBhn6fU
VHklVS9VYF/bKuUn3MKILEYScxqVu5s+T7WBoOEcYiE6MrGZRSbeDCOCg1u7ff6d
khsSBpQxScKkIa7a/scI0Agq+pGaCIaWkRyzaWbnp/RnDDwS22rgZDVMMdIRBoPv
0h/QtQGBAvbjyat83DQx36W91qqWE/4qH7M7SBy51RpJcrGz6DZCdCHnWr5wc3fs
boBoDISzuk8uqM76PzyzN6yHPZ4IF8Qi2lgXM0ZalOXFCXIAfLS+eP7PSjY0oXHK
VlRgpM7bJK2eeQd/qpfDf5gNqhMKmV0DmPGgQvDOYtNR9WYchfBUGSwuPM5lHeQG
0w1v6/W+r1OAuxv9cKM+j7YojEFyOq4j9IqZsnP1IOdN9b1zElYdENdYHh+qr++X
j3OhAt8N/+w7A3I7ycjVX5jBl5mgsS8h28z+l9tRrnYYasW15DFOXrTMpOv/GTBk
9wE5hV5+896KMC9f5DFuLaM34dZUuT01TZOl0iK8itjq7FyIrfMCXDBV//oB+eqW
bXZuVThZzP2zG3LjrB6csV3JQpE/p/OVV7a0pPheF7rfXvJaaGHb2peH91lTUF/H
on2iRZbtryfflFbjRxLviHAYlCNGzqrHaOCkgcgKvm4kvWlBcuCgsnI+0W+kXe6F
i2bunJrFYD9vyBqAAVVD6NW3DXIPXI3AspPI8lMZ+jqk1Fyqzqdo2GmbxX1jJpk4
4+W3O4b34FSpuV5zecTppDkDEFtVyW7OTAy/qOMp+6ysSbv9LPGk7zanlj31P6tO
g4/ERwdETi2+zhmiiO6AVgJf/rXBl3aG+pGUkeWQdV9H4qwFDAcfo/d1+ZpxBZKp
X1E1FXzsLaQzvxPxZ+rS9tVCQLz14SUdMeTzOtkaeSJd+C0mkSeTbGGkf7GsAT1t
GpVWiZ5VHwVX9XtGe6XZydgKp7ZxBhH6qQiLp44H3BOcZOXmtzdgR85E3MRBLDPn
jkjYnig0xIwe0uQ4VH31mUBqhqK9GrZrnklKA9Pnvrs6BvKyboJNQNajjmDoAhkh
h78QS9xi2mZyRwUEkumniNsqos277rUArH83df/3Wew0buORyaEmMN0wPf8LvPbW
5pvgWcU2NWrCwQcQ58XjqoeQhpjnyKmpDe0um2n1tlOyDPZSGhFGRQIXmdcD3Mna
JS40na1XYRX75AAglADaq8pM0fyKfYIACZ98QzVNSKwLH6PLA4/C2rxGjhFqLEqT
+McfCx7/YYye74yS85DdKM6xPTvQo7JBXOXFhIt4BMWDsNot9ouf0jQAAe15mGqd
hE0VAj4EoD6hiPvy21aIxVlZQkisQhJcEtPuAH/Z3qteUyki16pDK+qP9mRGjnEe
goSxM4Z2L/eE9d0JlqSqvi/z4G4LSec3d5rPK+8mU1zISJ68ZcP0NUp4FmtwdA4T
4ayFfsQdPIhvzUk970BPtio0It/L9NW981w60cveH+KzxzWnVFsw1EVHnTqA8KXR
at9dJE1dxMMqA0bxHdOuheFWF9QtYopcOYpI/r8NasB2G44suAZHOnaV84B/ENDm
FOnhlxwhWgk90pw0Ep7qQn/ikG7Edre7X8D1pu8JmQktoEDmTWrferUEvR+p8ls7
CTkFDESrdWCKRWuIFfqlah6iZRk+A9StVDhGtSjaTcTb2oi9YNRAH/oB7y3zO6JO
G1CH/3bU8Hazt6Naz3+GLr8VAmOLQp7bqfLbFkLQUsM86ZapbJEXGuqn6mSVGSIY
O9/+4BaIVIANDQZt1ZY8XbsjPqwZDoTry/YmfHRWLPgZ1p1QkCLO8ED03Pbqbs/7
RqCIqTdowKWVQ3yYF5wZkFB++9IKj5G8X0LllsadFxEEATkhgsaSibsHjL4N6LPU
dWAEas/gaRK90DkO015ivcnUkj0cAiADlNaiPueQSY/2rrOpu0lMl4/7txhq5H7T
KdJT/rIuz/xkREoUqWfJzSu9d7wYz0qXnnSRw2oCdp0RomghP0pMqC8s3reLME0r
EUyoOWlh+mYik4q0hfMVo95KoHViMaZmGAHUTo43GwaxWUpkjyLN2T6Z6m5X9H6m
CVgdhkezObuqKKASeyhP+gJ8nk2jDqKcSHokWZvInuOvOkTwdjOTKwGfKNJzwo+M
D2Xbn5oivkVNUnzimGhXBXJ/3Z9SQHM4RNsJFTuHeCjXO7g2Nn2w36jAtwXltmM8
c5X+MC93TXRUa03s/SoSl4I+os2q9EraK40ZyHFq4+9dvmkFqOUFyCBXB03VbfIC
ZY8QvsrsMlsdaOk0fNIBuHhYLPbVhUqv52u+ryp88GgvSLWZE7H5kcPyLY2ux/A4
Ec7pUDF60eSCyfefXe4czaOtP/WE//pl3N5SIufO43Wt5GEEemDsOPRPdBIySpQ6
ZFy/VGT2+Db6+oEphoBbmsdXyNe0Ekdby4RDWwS7IC4hea4J1sjEzt77yl0R2+KP
bMmQs7kn5Uf4XGK9pHMbDAkut0Z1ooipz1wLiWQdxH75Y9h8vh3qHjN8+l/1s6tT
iqV1/xO49unjxWQc9OsMc2fpRG79E2xSOFT9OtOxbKpgZN2wm8eXUwZH4cMLsMnx
d0F5v7Gs7yxPCeYg9ABXzFa2+0P0g8tdk5WtqOtg/NvsBh7WmrE4WHh4WrK/41o1
9NNKgbztpROl49EtrT3Jrqke51QHYh/LRZwkTmHvgZwQo5Z33X44N7+kyuSQ5xy6
o9DDkiwvcDFhsurpUxI5tVI72CBDMim0+SFp4Gfvfqg1aDrc2vBUzFqn76o791ww
yzq5uZWXEs2UayDNv6KlMqW+GorTjOIQJxnYphNfNAYo+So8lvyH8muCf9m7O6AY
eo1S+n/BtTztDXo+5jl6ob9A5FbhYsQJ2prp7EYIHGBwwOEZPGhvGEONMOOeYq33
SwqSQEKDOVn5TpM5FPtYjJFdDOCBgwzFrohE1fPKZoG764Nd94Hdu8rDGhvPWaic
c1tramGNjRISXbTAlMUAuuQdgQ54qz4tom7iOun1XM2Cv/WXeHeuu4PPp4nyNjph
mB1dMBdIgHIIF5qoh6wCoetTYlV74ujMGe8lxcpDCa8PyS5YDhFp0WMYO42jKjGF
50Ohis0dHzsBpWYS+/JjRWOqdXpJgvW4NsnY+Mus5ES62tWjb+WPjIpTGcNicmoz
yl0+72brY5nOFJPnfhGiUPXbxSQbBP/Osgnm4TaBG4Nfd8W9W4JcA+O04hH4Uz4a
EY33eIDkf8wU/JNhTNXPGUjxIVlXMTuiX13sSGVsVOe7eLe1r/6FlKewmEL355Xi
wbiZ+8PfjmSKs+bhF1mj1hfibKQGAFk2KnBZwFF8VPtR8bFJaPLy3SNFRgSh4oam
boAurc+fRQPBH/7Dt0O78QF558xGPvMdP4F9HdayljPQc/Av6z6Qd0cnNNPH1J9r
d425/d38VNNHbV8X2uAI/kddsQtPTSHlNMAh2es+25riHiqhNbzrWgWRiIaNaNWb
RRt6rmUdebc21zLb3Ck2EwfLpoVzLCaqGUGPi6M4XoXvopyav6+oDC7VpCRqHJhs
wVHZPskgcF2yKaBJLm2FWAhxT8tQbCq/qXmObohDEoUZJZUeGaYcjWMOf/fCitdU
QTcDWsEt2w6xY0zQIR9QhpZkdh33wDMHu5gfSpwcaK7vsSYdJBBrtK5QvOs46ySf
uwwONYjaQGQc6JE/IlVtrIe06lkLvIKaWqtaGsuceL2TxeK7FMRzjvITPTQh49jT
UQWVN1Vcpyu6wTek3GMj2n7Ul8uL8mkhb+EXuxG62TSpLXMd5if5a59RdyWxvibt
TFlpxCbkpUlhi/IX7sal1q37k8l/L6BW40haTwRu1TVoH6Yzko47LTkl4PPFc8sv
g7IR8LaCE6Glv7f+/S1jCh/TRImW17MMRNfAYjObbLbxsghBtkAEz5enHWm1rx0g
5qlSq1+5glHvsXLPWJQBDh/B12Xunj3kNiG1nm7uHVaVderrJl6tx+Hbvuof8Cmt
zxZhYYDYZGC9TDuQmXTwlU/T9o+vU595sFq2jol6nZjriEIc3Qa+FK/+s4XDZNUY
GlV+/pBuecpcV0C9U7fsx/in7J1J6ioHjm7IdwbjKN6zWuCLeAEkEP6dJH5Q0Zuf
SyOXapcHG8RYJ/5tTb8Ds95wf7DUadopNvucgQJMOCuQC7M+ZAgwBSwc+6pXrgqo
ou5UYO0WZfMFpd1PSkp3P+vIvy+fT4ZbrAU1PP4piIkKOCAUbgiJfbK2uq+/1UR7
OLngNi3nvV/xfoA27/4rOdb/yYS7J9iQ+RI7Rjs1deL3IH3YjIs3ogJ1LVR9Kakv
8yd8Ibps9f6ZCub8rZtzX48TAiwsiMzlewWpuqDHdM1vYZsYThPeN3FevsV9rSMm
1QoXRSOapP+fyn5TS4gXtprZRH25zCJJj9PDXkh1W4sScd8VTAhe6KawVwp+UAHx
IJure/9ftrHLKVoUaKKdtphH6PO1lqR3VpHHK6SzcB/AmmvxBON5Uf7RcUbPQIYc
cg9lWv4aDxZSqN094cdjbKGP6F9WNz5WdBb7DadUc44HtcuCHiU3F1Z857wMz4Hz
iasCWp6bwFe0uTXS0qrxNz5UZ7tmjQemO+/Bma0j6VPvk0xB6lKxRsbLzAzVYmq9
1mp5hlhB1qsFYYhUYpcL79SAwfM/ShBS7MAW0b3c4dIwkW8cMix7iFT8HLZtYqal
qc2cHTFl02yQ15/1NQwkI8tj/RKb8boB88AlkD4r4bsx1rwgxsNI15D+j3PKpl1V
TY2yxRmRVWJATRxhizLN7UbziuSUe9nGQTjPE0Wv6eSkPbbQl0Yp259+tmmmapsB
663WgVkOL6OgghbnRXKYg1wn4nDy1kml0A1FStSpIpwgY5X7Q+Dt+RIKrngzPrQ0
RNp8B+uoJiuABoVZwd6wu/mY0lK0MTdXWMXRxALWrUQu88+E1MiWpmyefAIlC3r2
RHcyfdiGGhwqFTayhwhQsFT6sDVeldH0V7Zq8qZOTngWIhCyyQ3sNIxHeNVxD0ew
clMWPLIG4HgdwaCcUPOcSkLerWoayJh109Nfe5NyNS6NcR2ExC5WwCVCILzF7+3z
+622xBSVYVdbXyCfL2e0jikBgEgdbi058jcVfXCpyfUfBtHZ9eTuMfSnhHduAhmW
FaH3SwqKHZT2ORhufnOGDrm2TIEKXKjqhOs9zyxREfioDfnDWWhg9YZZ8dSem+U/
+xsoRZx4aoR5cR+DLf3QQ6dU2lF7fi3NHV3cEhqLg5oXcaeA8yjEs5IjOxHAzc7/
BksYb3iNfuK5+VibIF1Jt+NLCWWXZEWZZfI/rJepDBVrfoEpi3UwgS2aQ4361kKf
ncRVLmjBYYZZ/+hgKgIwg8VG6PmTo8ZhHh3N6mfOy0aMbI/8/x4p90QzcIDS8RfD
CSO1R2N62gk6eIEYaKjyh1kfUpqzeptqKbj3eNGyHQ8jfSoICMKcgQwcC3APx2Nu
WCBbjZtm46A5zn60BZM5P7wS/0zL7nN8J8SPZOEeLDmurKPrIpJmIhxnRnX7okSC
2EA7jhwFLrq25HhkqDT8PTPGmKO60D8XLFlvZ1vvtXR34/iAMmmD+p9o28Dt9kwl
0A0ShvcoU4Ui98aA6CVwoTVgGzjuL+oYHw8cA7+irTyom7gUcUpTKlb2PFJA219F
yzjQToHKUGr9DrmR7lD4pDNBXc/yAAI60Dry5w8CU0eAbzKmvRYSeFrYdHgTqGUo
RVBxKQNlT4zcsllCJOR04TpQGsAt8oUJ0X7T7YNdE5mKST15xyW/mzT+onVHOqX/
LZAwQ8OGtuWpmaiw8I5aKo9x5Kc45uq3qL52EsLswZMriEI43nGrMX6SyM1rw1AW
R1BTb6qqRmgCaA2Xhs1Cr+7CUbIR9tqzgeROI6IZaoyhdOVYUf3kp0XkawA86Sc3
8mk6lm2DiLD4vqSZSRWYqfBrdZJMT7qufq+xhzG046zXAjA68ywk/jxlnXqHfe8j
yAd+N7NfHCX+b26kl2NYRq9WiNnxyCvG+Dnb8nbGrapwhyMpcMAnugb6SK/seE65
R1Ba+7lcFwx8L3n6igA0MpHazODNKR/wl2Hxn8gLymK6OOMEDNwzBNdHLGgQDS6R
84Tbmi/Z2cTlI2bAQWy4tP2ytyJcAhoZIgQ0FJjW7QCd79jbgkyq4fJa5Tdjz1B7
L1ReQVQEE1dmkBTkj4xD4lXyfD6QRmc93eRls3TL1AH2Zwwu0glM7MbpGafoeTUb
fkbmqTKUOIpNBeq+0s5fu/lrmn0iALIdDxG0zS3i8MXprzvjCRbUOE9oMVkBCxk9
rAArxNDC8xDbHiSuaKHbUmXcwF3aDh8/XR+j9562PNf8b7OnnaEh0D/GEHD4Q2Iy
GpxB1Cy0izPc1JclbO4vhDlAEQAKIWu7WxdpX3aUlupKG3ljdcQ0zpb+ot9n6dc7
T7piOVyaHPfIWODx55CLBmdMNqMWesWAz0ihdALQUaMSqn93+e/dymctZ0walmyL
18+5+wiUBhrm5FuasnoeZa2Q39xorDOwiG322IHNgEnT2KMnLkOEVpOqgr5hpAFU
VJ5f5CicMJpCntfLMDThl8aCgBS/qz3E5KxNuR85cnDahKTiOeOSpVZyOEBLWXGP
SJYT13wYvYfmYPqKBKxmSHg2tswPtyQANm/11YAF6S4IJW5VkrwLcBFamRCzjsDo
T3kWyJ+OLPP3fcfYnvjGvyvjXASgDeb0stKODZsxAbPXQVtUmbn6Ak54G7yLM9co
2owTmzyILW8tu9L1L7qMKAVSNbC3M6yx2uNS8WiGGNuYLTiIjRXd4Ap0FXZW2c03
GpWWToSFBa6rhA5xPTJlZjw2i+8WeXIMSh2fjnYOY+TTmr/vNCH1YVuv0kHPKiRw
zAMkLMiw5iZvef/oFIAH/Yjzb+Knz3MOD/5u3N22S3pvocLv7D8dobGW21Agxbph
PmrOMrlXU6PWautFe/nZ7h/Rrqkycp6KI2Nel9pgc+F021bB8UJOX0nvuKkc8vfB
Z4vRpzOg/HbRTSELBBqdFyuopzhA/BwW2H2VOjSWdeE6T+3PpxQ1wNb13Rre6frx
EVxvzEmHKYB8ODPoADw+vftrUqrIm5Wzy09boiHxyiDNCcpV2P6NhJJeKKzFPLAi
/MulgpX0byukS3dSjHnhnl7Wl2peuZYpZT88d8SyUqVTZYZmVarbH5ybHdUetzta
VbS0ST/RAC7z9hX1EYcwfXp/uTZ9PpPxWw1fVenCgeDmUuCYZ9jDVSYRjBe1rUuB
OCGZZG/7fE6qKYjCtiDfJRwFSLMp1NB1ysNC0z28xmfcKnqb0ry9hf4CHTXiFL4U
gThdr5UaUuHwtYOZkuQnrsSMVUpJirMqELd23FeUwsB6UWuvkYa1O4F05hpErlGy
+FyTHK6zYCKnM+UWGib2O3mhQ7dIxmA1W58KlmxYYxo21kwPxsuwwCwmc2d0vUCE
PFRxeoPbLX1+56dnEu1BJk+3Qhw85r/gzqlJbMH+M8mCaATPhrg9rMIjAXX9cSe5
RkPMT4QFuiMEoFcb8JF4xtVfxlZ1eSsFXlIaz1hJDqkwR/anVrpJeS4dpUkInrMA
cRx4jczWKydkBwBw2+YJfNaDdsicNuH1/8lGnbtTzVGoRZmKMifnNItxwh5Qi/hR
W+SbGLROIiSfovhZ5/B/vuiH61Hng+R2BjuUq/BxUXxFoEJUoPzgfAuF7t1MN9L1
+2mpK7oIqet2tK5+OGHuUKZ9/ns6P+44p5rPO3UeftrsQx+jHY149VlDENopbOwb
XuLOfq/WntugF7f3FuYVabVOrw4isOv8yO3qfmrDXJkLFOiNl2d/4sUDXtJh3k/n
oPiTZIa5jK2HMKeIl77h72Mv00TvlcYi0BAVzVrdm3keAHTlSwRtc/kSfYThJtB6
TUq5Sk4dDkIdGCUAhDKKfBXg6b5pLy7nE6m3v3dJugeYuVTK/ajkgnSPZAFA8N6w
xRim7tjrrpshFKo4Klwyg0ERQxwBQc+t/IIPAG2legOsDkakkLltkxoO4hPpJ8AL
5BkXtawllfK+Jmm7HtzK72cG4Ajn0zJaFvlTOfvsCdx1/UkObiYcvpDNmjB27OQJ
yv0+6TeywF8RNlzfgb0D15Jw0Z0g8ynhoOgsBSHjGqJ6+VE2KoEYWx4LxljGt+zN
MlyCfc0R3g/SBvbavawucaDa4fdaoFIVXhwvYhv5k6xv8FyZtV6HtMn5+GOJn7Qf
4PWuMFWnfMYb8JDokOdswlSGyuGuownQThk0K8jWl3yUdtTYgY+yMLUgVb/7t21v
w1LvzeXuyhyaXksUvcTbAx3AFC7CH3feRK3/ElRil2upKDy8KvPbJ4ZOvL25mklI
SFfphVD80GrUp1w4l/8Ol6IkJFLjrrHdZzJdh1bLLCHXHrce4o9nTcIUzrfk4zQp
OaSkO+SNB3B0WmgW9gRYk/rnx9+zCKE2eqUV0o6pE44QOwIfJ4+17Xax1oKPS3a5
q4xxSyhv39RELWq4Cl6YnU/9ZdnPHC255JswJKyAFxtLGpJ4opZ8HDduQ56DdP9j
B+5IMJamRz1gPI1zXHyQJe9F52vytPb6K5pc4kdkNB0SAPDENOU19cs1qkgUkzmm
mXQBMR/rj0TZSCRUdVCX2SG81z4m2VKuOfRFP407IuR0KWnsFg19AI5XN1bCh0gS
OxJQE3orCMKLvEQiR2+8ZaG2N9uh6YQFj3zr7WIlvjdWoxvGdF26HZNMQ+6Y3Snt
QkH9RlKj2s62FY9LiG1Z4FarIi1YLn0JxMgdXjIMEIb99s4mqILfGxdbVq7uUjze
7E0ur1eRI+nxqfBldwY/D2SQR57K6hJPYrzRZznLb2FoQcv7BMJFJgN3dcqRqZuQ
GJOpon2WGnsCo2kwCIjtdnWoIcdPJn00U9wNOOSxgJcx2Ajajx/290qV2C1PdjxR
p8zrKTmjyZdn5HIrywiDN0eGjh/xQLPqvNeK2bHDpu3xOwode9eyU1ttRMcix8B6
IC34ivO8EKQnXFXtzvkFtZnqnx/TI9znX1e69Yq46Isj49pZIyn2qwRKGdoaAt9B
2cDpybG8PmHrHdxaJJr8bunX0H3NY90395HqawUbjtFhdDbsnX7Nvsp6JHBzK9Pb
XRrc/IvpADElInh/gohf97HIKSE2EXIeN4mez9pCEhB05cc9Y2IQOojkAkR+HyYL
Misp5iz1veNbWPtGYKoFEwngj85PE53guvJ1OD2DKBx4YnhV0V9JG91msJtLEqPN
+4H0DPaRDpWNpClbfqPcpxqknPtst/U4mkJKgCEFpUgTV6WM/xThBZo3Jzk7Q2+S
htJUjEbPA39TArdTzRA9Qkw5fSO6SmORy79ByfNNlRBecqjnGwj1QZlwgBQLr1us
/+88CIPRC7Wn6C12eTdWPnlekICnkyDXDdDf0x7mfeE9grlszmpUTPmD9BzHMHBA
lCCao9Zj0k/dO/BTQhazpIqEK5CZgYRTV5yetntukc9aB0eWh8VlDzIrQmejecNo
tbi3zM358MF4JvC18I7Rf7Uq+8+U71dPXIb9AjQt8+Ba3+efPi/F3yHZOCrH1TkG
tbdzZQfDsOe/6jgau8WfyJuZ3c1tamHhbXS+ySOIAlp5CaoBkNdI7TaglzS2soVm
mFqXjHoQ9WCPwig376r9ZVQ1GnY00xyoN7wP/Sy6uJqIoRRUhR/xQXxSAwilV5y7
zAzGr1dudqo5VN76cl8Ov94PSN/2HC8HrhMs4vmNj8XAvLwiFUHRdPBTkIbn7b30
traheXCZktUgREcqi7PYjERX28kwlNLLDOl1z9h2u1ySZPrKf+0BTduiFnzTusqY
R5O0HhmqKsptjbP43VIe9Zk1AeI8rwYegRW4fMNRo1y1kKPyOewfxkYan6GqXhlM
thq8wDT+Nu3aNtTcij8jXzVwwK3k0hzKVsuQ7lzbpBL7JX7YOUixRTMJxbIGuG0a
zxgoyG5a5mMNpcbzw1ddRG/hl+suHwVJNPScWFDSed8ewD52VBBxbv8/W7Pxw7e+
zZDeVo474iSpJOG9zTOR8fOdGEeQDYoiuIWdBfSj/xc2UHRV8Tn/sFyIxcZAvD33
67cPdH+kGxd/DzfBsUf3UlBazYAbrlm+A4DB45WVLAb0splEtQI10JTXahEpIkyi
XPbQimcJ+e4mVfDkcQNIGdlKFuZVAo9DgjlT7YvvwFdBny9r4TdL7TgeDd89i79C
DnwkKJq2Nlwy5QC7KP6UMy8s4U1QZZLLdTFvhszPS0f/Wdirw6pbzcA4cIDIXWVP
MvHYAk1gB3wi3q5K1pefNxt4UUDI2908SYcdoufG42808GaQB4ol3I0YZuhUj7ni
QwXp567NnhRJ7eu0gmGPvViXpwzbxNJuH7BaiVxCkf48xUyp16Z6E+t8t6ecVOWt
tPFUMcPppI7ZBuTpLal2WD3Q6WApDAFmlTjctygFIk7KRboC5ppGBlPfQ+gIKOhE
GEj0lxf/fKfV6itPi7ZpWw27g9Am7/pRTFroxAtFhZauOIhxjrL23gxkRwMoqlws
r6vNUnBmYJT/O8H3WaQMyp5LbJCg/jmPXAA1ZXQ5K6X6xTciSEcoYUuXYUrAIxwS
XSZxSTQsEKPMsAgG1CxVU1lfkJUmOmsVAxGr4zw0k2mN/jybTNj9NJyCImpE3KKp
abp1Gxl9YwAthOLmaRDfLR+814Hv8Ly56EVbmTg9EcOyXYe2lhTuZtyQns2x8y/L
RcmvGWyL/V89e4EfxVjMDoHK07m9oWl3Zl8Pq5ssqJsNPatbdGn6zacnu0TC96Xm
hyEKmT0ZtdEMNnJasoLo2aT3T2+f+FHN4ZsNF5a6YvpkpfO3ai1cWrfl/NvGd9Yu
5ghk2y6Lg51eqeZZyFALuWdOiIkYI9jdf1fdCUA836cCsGWXBHWPwI895Bgym5eH
Jocee88EFtvU6f8RGq6w5GLyerIZ6Dx4xxUkG4dxOovm7Lf6zrv7WXiIyChayHBd
mNs3sbpZDQccVEO0gpZ5a+quy8FuQZ9J/o/lRsjm7HRbDzo5Dydbs9JAmMbeWDUL
tPtvaa1ieMLOC2q2QDmz5yavtGUx20qoHNvKO91tb1K3SRgX8rJjSXvSJINxnYGM
Z+/Tj8KZNOA0xCNxSKkjYCcTX5eH7agJaVkx3axo61EgpdNr7POjRM+XVLmrKoM9
9NKtHAhmgXnA2q4ymctqYdnqkU1tVSTMvH9E90qvTPuVVxic5OEC2Ih3QUdjZ7WA
2fKKqcFJ0F3yhH9rALTJTcW4eN+ayLXtSr09TmSsdIkcysK+jVjefI5fjFkxeLGi
kADKUgQSLMc/K1wJh7/ZrpAsJvU04ehyVCBf8ZKDGBhN1f1etjeBoEliFyg42T6T
fIagzLmM0zn976zH3vBDJWgFHtvUdpVn73WkM5cpCVYeNa5SlY5nOCET/Xt/xJAa
rUWxWa7jCJrWDJYOmZHRAi4KafT+OseZqGsVAmhULVHe0ebjbDUUHia7799yie6e
8npiPgiF+LRvgnHTZd+CHTpAOBe3gsod4mlErC57GI9RYkDYGXtIEDaKhfRUX6jw
sf/sQ5b+K/pGkc4ZaxIrIqaMIBZvyAAD3hu9XztL7bXhYS7ccP71I2o+B+3avVMI
nkB8Zd4tFMIsqLyE8ALDeiumYe+ApiaBzP7p3Yr8d4bdzmP1HAH01wqnOHQV+Kaq
cwhFtPtYKisY3/zWIFgIL/t5AyT6peOuq5gknQZgfhBI/G+ZnyGZ/R7wee5kwoZd
PCPcpd2laor76gMo8hIerdx0hupho28NaZlu61b7ipX8Jev+cwk/FqG35giq0mMd
TMgQqwFOUqvaJsukwBrESpSpyxQIxtizaymypwC2IDlO0azS6miAoUcqiTNj4eS0
WGc8CSBXO8fFNKAsd9gUnwZsUBEalmU0BiLqvnSg2x5nBxS0xrcDktuQJVxtctvi
QJ1BIaw0D2KEyTqcgV64vXxc7G1bIzH1vGbO4TwjA0jcXZkomz03VXAchTNjT7XY
s2N63BBIEOcMzOLYhtphKSKJxPfUdFthB3LuaAABSY8Oxg77NEmNZIqqHEHXvFHJ
5YkM4iL9MIorswarrgKtyK3Qiy/tmn1Ml8jpTcETpoPhpOeQPYdAR5PthWi3VZEZ
S0ikXN5gqK7/zXufPIwRDPo1scZbtRr5q4SqSMCbMpAd4EEDWu6PEk63+GuMoMU5
nagMXAQc+kG9ebmD3BMP25wW8NP/JVZvcBXHSxF5R3BTplAsKUDfbB1e+Wq+9nD4
YP1dqtu55h7R0y2T/ckrISYDkqGjn1OboXf/qJ7trgTvutPxnEx9euQLwhBVAYFw
o7twPBg8WbZKoTLyxb7Bvh8/t9rTiVTUXowkPSk4BevZcoh5LWy1XkTc6URM8991
1PYy1wSJBaAKSiWLSShqeZAPOnif6h23DrrcfZ6XQoD5gV0B8Zghx3dyWVt2sWpe
RssoEWEwEbl/cuwoHzgsET+3dxe4tc6Wz7yuCU7lBu90u06sIKDrvQZIYH2wWtAK
kaNS/M2cX3aghh2RAIMFUhS8eSI17LSPaQrENccw8aaSLJG5/s+xG9X/JmcYo3MR
tJ1+E/NOdE90Ooefnw+j0nqR4wvLSHt0gzeviGYh2A2MwvrDYy0jt4vKAt1Ue30a
ovauV4vCcrN6MBZj9Hqr+P5/PUsfB9WfxHR++B6Gq00xibSE49Vp3K1PiAQs9m9b
MsY1oO/s4d1+QKOywksKIjQdiV0xVkWOiR795hl21yjRd7mfduIJYinobw9OSnx8
qq40jhWK4OnoqtKFILgujyQ6/EAT3ZmQ4BNke1yT2RV3zxsbSsPr4b/3Si4n6GHy
pe6qcsPFvQI/XsVez02oAg+ua6QuZlHEYO5RdtACAk7WVJ331e/MxAVaTil7j7TW
PsCtNU3DD6fjnJmOtx8zcj6DxojDMt55ygVwvcAmvw5qa+iQT96BmAzqznxnJynY
uBjKR8KyWqedOTherD3gJEIM5906iXnQi+bET2yOtT1aXqV1r3ts1Cr1qW4dzRMT
0+ZqAgaBVvxT9zS4hxiF4PU4FtO399lD75vbfj1WROYfZEhTkaI34XZAn0DT4Kuy
NwUWOOtLAPAjOFNgeBdzfjrioo+311LiUzBOrHZ4g6ZQDNrNw1LGPKxYe2G6yCzQ
G0dGFqi+88/wPHBq2mE/ginF4DRhduCFWoEIcSRjmG0f42dD97Cu5h0gUNTpMxC1
sEUDRzPUKoxxHvSwZV1M4ZsWxjGxUniwsN94NWZJE3h4mDZx6D0Sw6S85qC/t4Aq
kESs0qJT6jcS0XIBqCSrPNyKUiYdQ6RJdrqa5zl9UvDYT+JgNc+cj+O3jSR1mjkK
A0w59fM8JhzlGw7MsdIMDvDov2iYe/d1KLWVcTrddJI7Dn2OOPz6sDWr2owacV+2
Psh+QOwIqd97ivTltkteDo6kt7b0wrXL3CnC7ULFg5NVV2iusb70Bsu4WEf3Y6zi
WPnrX873lqkE1Jda6uhvCBmAbvfxfmE3eWpEtthC5vg4EW6hAwdkB1io0MbzRKFi
eBRlbwC0/MlOF3SNxfgvaklVbsJywxUJvcyaK9Cypg0HtLzLo+0CWEverIH0YhRC
RtaAqFnYC+dQMN+fmpJxsv8nfIQutxOT5zjqS5Kzy5Jn1nfqJOqT4iy/ta2qhTo/
EDcj7wellNfUMbcrNsUEgDI186Qh3FwSsdCnjHsnEwC+ERQcaQJXugL8M+NiwcoG
RVYi9OTYdVnL1C9Lm0hppEX1rwutqB0OG7pSEt1V5JaKHRk1v/1R9XQpx5Si2zjs
Bxde1QOr45aAzmUEu4ZVGad5JzkDv4c14MkA12ehQQG1MWkwsWpUlWWtJphJS5Zt
JpBWDJtfjuili/sZKwx4lRAgv2YGbc9PLr5ooiWII/HV8leWicGs1ac9doyOElRL
Ih0dgR6xkC/87CJhKYd+J2Fm450ZXAsuYEmSYUoLozBJWjxuZft5zSoDlnffdAI8
h2q33o9BVRQsNiaikMDYjyh+iUdGsB1L3BCEiifXMEWo6XRsZcYkKLiwGK2H+ne6
hQtsIwdGYVahGBVOot3bxVtDI3uzuiIbUNw///fR+LAIKn2M2MlJNCqnZXOJuZ9M
kSNwToGL+N8cTDRB53qfDNiPSx9H1PChlu3oSxzScoHzHK0tf/V4cGPxui2ELA0v
xYubVNc/Q0giPJDiVKf1KPaxxZQOOWN1tkqFrEX0ThULKZE/gjwV+95ITvPrQAHX
FnhezD9fe0o2swTdpn9a4XlM41nJsBDBYLBjP9qYbjtEK75ENJi3fTBS9taMtcDw
BCoJz5QwbGgMJOeTw1BpBOTj/z5yAWO5JrfBDTycDc09EAX/5y8+j+zSI7jPGWGL
i7NIJ8+ppSgpXhasrslfEX0OwzuK+WzKZ5cVWJejJu7LY0Pg46L191nwiZw0rBjw
AzEUONSD7Z0/VeMKJ4k/5iY9C11YEsHDMUzMkSzSn1BotTYiMYfAcunvr+TpV1WN
0bZIEj/ST6CF6OC8/hOR6MgIjIsEiumP8b8C4voIN+/0XWdLI8sb7xtfxNRlpu39
qEgeukTyWaTnzeWdGgkgccXH6UAhfcA6/96anX6fPOx1tEXfmZuovkZSBHatRmlU
I+7kJp1QSoNFF8lVa769TinkotxBOe+nGBNK556e4k9Lb2VD806Cd/1pTSw7j1Wm
z5kRlQIZjcgAhfkmNvD8HvPOlcxiPJGTiXtpV6RiTZcJq6dd6ESKGooKAR8lwPS0
MnjbZbD9rT8fT/e3Li8k1aD9UuLK7UTNvz/wVEe6tb0DpcrDSfGrK9bW6IikeOhf
SRJ1MhZVnFwVeO+v9MyrpGkRc0QQZmMG6qac4bVubiV8VAKhRPWBTyi4JKJFAUoJ
tQrjyFEocPBf/ZjaoHttLKR2wuvL0FPg4DxkEoj9zJUEGuy4mB+2h57XfofxLtYE
RZ7bhq4S7aGh8ZXNSb3EHnSQAY+SKgPgmm689uxkoi+4Fk18mW7vQntuujxaVJRr
2zu8s1SSca8XBw2eLe7G29TsJR74jqSMgOdDG7g2v6/gqisfO47MD1wJaYauhai8
PpqSSB4F5JCNq7CJMXaZPfrapC5ISCVOchQzMiRQIzhIIx1nbOwwTMVamD9jvoFp
wcYnQ4OKYXlO8XWP2ZyHMQeKLnGSpDGAOcPyPSAv9/jh5sxrS+RpAOp2M2tk4tE7
+AV7rDT3kBZKi5bIqv/YYTrBm9jpctLJSNMxkRP2tAYuhKMJTkxxuqQ9eM0zY8bQ
y1pEJ6kL6Pcj5P7RO3ub2jG2AGFuom7AyyVqKIkx0671Km0txZOwe86RVLbR/X/o
u+ot0XVCf3c9PXyVjUxSPGwi8TrJlsPpBvQX8zSVraSJgoGsTtNLTosIpNhDilAx
FFuSgjd2kK1qdI27sPLIoVppXR/MQZCqzG8NNIUBX5byXW792Um1gR48LiqJ0SOl
h3R90jiPnf2+oAqbPHJlqKX7O020Gzp6LtZ4AV+knK/oPJfW69+1L5/zimjIdKDo
+jnlDoPdG9u5p8w31MAgO6/sa/46RbBz53CRTIuQMmmejsn5TgfV2gnb8MAOOHFw
rhHfDbZ8vIgh5wsUkQ/9J2sqM2B3Rqlnd+KS8o6cQeivJWJZnxhf919sX5Tb0kEE
UcwS4xhO1rE45Q7M8At8P1jioJ9JonoUuMJGs0XVsgPCoPXYg2dSIzeAf/dxuKFU
za9pfgXHBausGO3vwAtaCHBt94ud0l4JHBmqRyn2V758qnZdfbX/zSjqfrXVZXpq
78eLdX8P6JA4Jtls6xF0vHWkuMolgFNRuCz6wBsswGh8fNalqA3E64udvux7d9m3
jl15uE5ssBHn1Xd5b7W26dM+nZ6nUTQVskMcDZ3bwVrDzMtRhT6Ms3jEMX8fzO9l
gZe8Hy2jTdh/Abn3l7IEdLbdbK6uq7qqFnlFBiUBx25g8gzJ/4CdbyhQZDQLm1uy
MmhHZLactUxq/SPlbFKIwC5rBJK+kZTXXmvgjZk7i/8bIkTujerxSPRxdXUrxREh
OkNjsNLkT4I3FidGyqT9Ihaw0B7NfupMSXfnSgbZKBmOF45oEH0okpIp3JbbIOnd
wAvWwczYnK7kkV6YngmCvHKA5g1CrFXMSTuQfJiW0TO+CqF3KiepGknbUFoGKumD
771fJSEzvz7gme2nfkx0RKIllkJ/USJjzsj8xBK94SHwvd9pco79+chxVGHmb2XT
FO/h5fmHrdHn0GjUVzqVTB4EU5t9eTzjZKmqU6W4JWhmGAsgjkDzruJZ4dKYxIfA
e3+qKJKDDL+D2ZvRGzrP76r2a5LVIEKfsYvEBotEMsRJeCeGVaucqpiyhrukXY5+
8WrNcMpvIhX6xlWKaq/rl6YLWvOvNrHg+1/HFXmk1x+AvFTGgQ0g1+9kmyXECIR2
EvLfVqcXKuxFPnvyLL6Io/0vlhFX57FDPbJxwCPT5MiZM/9H/PzcXw7rj4TI2p39
nh5EO1FGiWu4DDdmK5Uk0JGxP9sg3nFuFI+Chd0I4TSOrYWeeksuJD2LKwTiNG5q
tY/x2iNELSBEdjUdE6BLPlRz2stu929IZg7urtxMjTtByVyl/AUkZGf+qlDPUvhs
1CvT76KQxL8fjMFKR0YeeQkZ8TOsMHlz1AjHHs3EnXoeTwRcmWKUi8ImLiimbclQ
IIS4jMEfLOxn8QVJSIpootzV9HfB+BPbuF8dg35hj3L0exJA87FLFEcfSVomDR8n
EYWW94JvYi+r2A6Oxh7OyDLIfzCrI/6wAOBZcS6ugzmmrNBGjwCaZ+ae6NtupbvC
JIK62M0x+36FUj7buLl9XN6x5KlnpAtQkDanfOs6j8/V5DKTB4vxdjqIPfonZtbe
4SaVMmwE23MbTC5CfxvHXwmoYMvzWGCTIUN+iJedUUhtVlObNueaUT3qnGNdR0KK
xFNxiHxhvkveu2wEXSa8EfISzUKTeSaII9voOqAAP3s0siWm9pt7JjdDCS4GuyQf
YhbNdmGoSigC+qAUtiaLu5Mr7nBG+WIpencnhv5ryRB31HxUT89xNQf/jb71kIvJ
asdG9atUVpDm4GbB1a2HfpNz4QLnadmttFkMdgvwOk+yQvEYaVDcRC5QsFzsiVtb
EeDmCGx8X8PrPkro6BagLmTcGBKYHYGATYepuzDI3dIzUzl28MZZ4tX+nW1XCz7f
p+0OpAnDKB+4C2zwqn1YYGRcYYU1Ih7oHFOgGUs2HM2ObYHBNk9AZAK/iEeRscXF
xRZg02FaoH2XfFnExEAG2l6SA4mhFMN7VVOZIEIPbkVXOAjTVNrvLPv3afQZplgq
v2FUPU/vGF0pr6JQVLnNVsAed2DmD6XCvBbNbqR/Nc8r0/TC+5F+YLl4wVvushVs
AlsgJvbzf5s1PGlYHvK3WrdG7aDl2yk02I+RmHnocwhSxbC+PNiwnKGpcv97jetC
YJ9hKFJmk7NWnhZTdTHHahMQED1RV8NO/qUaVDyibTWWbZ0Y2IXj3HCtEEMLiJ8+
JwXahiNdKczxYcb+ZkS5GLm8Mx4uU9dqx1uLE1QnthS5Z3WLxdFVK8sQMB6jMyD3
tmAIyW/Jlnkzj3XuhDQSwwd3a+YDXvBmdVEBSMPcIWHB/pwWvH+1eIfGPCRZReBz
0d0iCMCicvZN6+p3IP2h9NOyuPwB3u76m/vSeJXlpL702OQC7d2iRIvGVOJn9A3o
W3sfaZzfZr5UC+bTqostj3XSKKP4xF9hufVtCvQQiE6Fx95+Odt+oISpOWKO+K3k
p4T72a5TYteki3SYQcAkc2A1S3nX6H8p07jUTrAs3ukFV0oucm3Vl2dgxxI6EVTR
WcJUdxEtONNCdSApo9kV2D/lW11UZmW2NMJwupjj0HnS38GXKTgPt23m2rq/vyVG
WMI/p7G4Duaaml4MH3OEHsv6Z3LTFkWqvlJMib+fASAsxw5SGv7IBOLOpEaYiO3d
XTdA8h0rSmWvbInidqcwNg2mEdkrVcpqb3TOqkyL6lhhQiwshqXmtJouDMNSqLi8
hJXJkBM8sOY1IX5dqAQG6Uk1Vd3Kd2lys8ahg7NLn+RpI6PcOoblbd9ZPE4HR1x4
3EbybiINhy4sHhx9Am7nYAdYwQmETh/mzMpMmbfDM/8/rPw3T2p1+NRYyc7ElMHU
Q5lidHtnEClaGtxRaFtTSEkgjcGZDiuEAXfi31sFtYg7nNuIgATwsnyXDPARx+My
g4+P2M8jj3hQLLfNrIwUXEnp3dphOBn2z3b3eA2+7/5J+Q6vlj3irXQFjSs2fbNc
e3IxDGydmNGSJnMFpszfhwJGFdxpBxqqqMoUy3gw/36+CodKPWBdaCaX/71UR+s/
4NARxwAAHsYQIwDji4j8RLoFzIGv6ShkjViOUFLLaPL3/GDCAAUYixnFSE/3HWDk
A9zB7NMqkVMX9AyqpiRbElrk1T2nlqkbjJcpqOr4ECC5pMUCDWN3Pe3wL5Yqu0PJ
IdqDua5f01g6PQvhajHlZ1cC8CpzyxGTnIiUToWxLfzyGg5wByeT5YQnuWJrP0s/
+5M6x+hwBp4hEMfIDXxtbVOQjs9+pQaPHque5pkgbD71PWc3g07AUSHeQreeKxqF
/pbulMR46tRTocTy2ajxOrHQrBIkreGO60ECDjeIM6S2/nmq2n8h7xNPEVD4BfIy
uesvoq1Du0Vzqu45UC/ijCuQneCbfvV+u2Lw0D/rb6yIWh0sJMGIiS7p+zRPiI7J
vbNmuDJZyekcQAjnekvsJlWD49Mhb277GxwxxghczOx/+ycvWym33cZNFjtM1Kn8
G6SPa498aHJn5O7V0OxPjYvPAxKq0bNrlMoJIzyKLuf89AlvH2VfUeneAi1jkvPv
BOor4iyqFBJu2hqd9o8LQ3ijaWjfIpkOKgMb9klG/5SADN1w4Ksza3QD/35oJr0e
zYQEhKOj7bayD7c8buDnu2NCrHxPQZhwSz80ts8gSbZC2LIQ/k+fTi1QvLLr3MKb
SEJIbhXOMdk1tWddp6dLwK8ZjPdGUKX0WxedyYlqV+jhsVHfFbGwOU2095vLdZbD
qInXac+6u+pSJVvi+qjhZThlsU0ct6pRx2Q0YQ0SwyGqf8trV4XBhf9FEYWHaMGs
+vWZ8h5+KkTMHcX+EbhmRPAs8qsZInaeb3gttm84zqWvF+i+5emfTUcM5IPCe+B2
iQDHHRuHKPrarZ6HfoEN0ketKYJ+uVfuTizZNecofx35GTgBIjgjqN9e+hGcUIue
ndWOmefMhHI3vxPtexRkY63SK3xW3bY6sonO0ic2yNiG/K+bq8OC8reamRGOfdAK
xaukV/MqtqGbwMAw3NIW5RoyszSRFuCg+4j02oPHwPgFudksucesV75JpSTd+at4
sJApduVWIkb7BRBHuATGrfbva/LsEXkZ/oR7uti4i3wHg5EWrdMRHoakOARl3vXq
g507v29O+9eKUaMcfinzPHdbnwkSyZRonq9kMnrWLyH8itjBil+SkVR2fc0qoNAt
aegTJZyaTo1T7hA7K/J3QkaLugStiXF3InS729y8mOmBTb5mMSgILjWVoAnFcF86
gNe1YZGTakSnl2zxT4oaJDif70T/Msk7JvZ2afvRL3t5fV/WJ/bjjo1KYapETEcC
PHV/7XO5EZ48anamqBq1d+LhpnuqdK2cN/wXchpG26N33p7ScgokW4zYeAsfcwL8
1HhwxmRmQYMkDD5gSQivNtvynOogH2o9nVallHjfjYijl/Tle9L2/VywHzoPUnUs
7pvwIW+Ys3HI5+zxOCRIuYPMsgg2uarY+UDpp42BgKVcIpYWZo0nusefmngroq8c
jFa3DVDPgPdjPw4zWW6rEWI/GRiUqB7+geiDO/DcXhlpoAm5kYpomx7Eo6qH27o6
RfW42mYx/bOCnvyi+gFO8yh6mTS8jxEk0m9TlF4LlSw7Da2DQ4/vlV+LqBRIWCV3
gdXl1gP2G+e8tdPL1eP0ACvCFfZ12nWiKh0ZLynEQVRXDrKKJOS3pAW46sEr8zDZ
Apuj04W2ZWJMxMhZd3+IMjCwnfI8+dFFLDf/s3F+B7NsbuUKUwf5P6iZQ7qgWYSy
ynAe9PSQ3TtOH1+y0Tm8pWpMeULblkojE2CZrp+CmulTzKGkZUTRi9e+mw2PUPtl
3BkMgZh2FMLB8UihgTFe3n0vGcAWyrN7Sli6almtPLNX1k+wO/EwB2v1IUhp41GX
4/VPdmcmRpPUpj6dS3Rwr/ktCUQcu+y64bmeLi3IA63zjeH8OFbPJOnldmCsoZ0S
u0oa7CALLYNl+7RRZ8evaVnxkdEzkpmhm5QS2VLjZaHterCsjayhNxMeYfOVlgks
A4WfKSEyuB2B2BdVRlqDRHzjuTieasMhWRGQZHoKIwNtnc6bLux+T37Qn8rQd9x7
17Lg2Gjx7+kRUKAmVQm3TdueO8tF45Ky+IVR/3vqGB2nhq5Wxr8p4AI4kXvz7wi0
2dPOR7B5AJ0oGFOkeAlLXSnUypz/tBQliGfvbQrqpvvEmyEYGQberMN2PvyDkk2I
I4PfcaAmm3sISAg/rFCdoOCCMbwNbxPbPARmH055sbGVAA3ROvi3gHMuXqqpV2FP
8jiMCBjcbXFdT2LroukUSSAHzEQ6v1lKHJPs0xN0uDmCVhFDemx4Y6l3t0seiQyl
w4BJaZRRByQLUMlOYK0XIbucjm8wyCGHzFdZ/bFUsqRL7VAfJH6+YtNGMjaNo3sN
l+nDMJQEEGZmWfWC/wHYxnxXvz37v1uXdK6qlK5Hoo0sdZgtUPrySXqtDo3N6qAx
pF+FmsBt6LeCD0YSCIZsDMacRlJ15ezJSZl0sdfkbKYlXAyzX+H1u6G7NhZ0V8/S
MCY4aSFNXLWDJSM2VSUHh+VfZHAPV878B8lUxd4PGoyGC2RwFUKhOWCHGM+xOdF6
yRehW9yPXumgaJ9sdNPMMkwGq8MxPQUN8nGLd2KiBSEorn8e0gyOHGiQnsBqilL6
KjvkR63HiuypAzB5nMEAhFEtLjLWEh0KeKNhac4nKLkLm3H0NMopFpNFIRJuFukt
UZKzgtu8/BpqJ61zgTTTkOoya02gr/IOnsj3EDnaqrbYsAjPgezF4ivV5rWCjmpd
JZm00vuAxRCP67ZYF/6YhEszPh4HMiFYCkEzgsUG9B7O2untCpRZNWTjahdPR1iV
sDHWrJ5moGtMOLfl+Y7iw84aLqmKI0IiAgKdb4avzjDK4hNuCbt3dq20xBtoFcnc
SXKZARXhX+9ATEgg0n0yvPQl+i1hGw9Ser8AnZm/sZsdUUKCEH2muXpJiDVqrFPs
pRuKEWWhs4zZNRhekQLe4ZBkZ1DQdBFky8gatWyx49DXkUwzOHr5ohMKuhuAMbCO
0z8dFyB/xdGlxyXVwRiYo7JW1/OL42g4dqSbmIumV9dKM4MFcuEKPDIjuUSeu5au
Xz3qBlfOu0yrYSgNC+92+nXzTI9VegmYuzs8yfBDCt14de9NH5IUW+dODYLFNWpJ
RQ2zeG01M73KY8GoZYbQnlnYIEsGYrJmMcWiocH0BYttGaqSF8uGtDeNYpG/KCIE
g9WrOOt8C5s0NbZoI/2nV8Fo3hzSSGzvm/MrbEGXpnmSm7tPyp3h1/bJRonnRfmG
isnBgauRYJ9ejiplfTQYiGaAnImV54Te8YXytDodwrfrESBRj6sUzgMXVc/QElGU
3GtKGGssweBWIoT/oloZH2JNMW/rO9LfyoaHJjgN7vXKTpwvHMQuYVMtdO3U64Or
vxTS9MM7qydMx04ZysuHHdfwRD0CFpY4T9b6yILS/srIDKjMofAvSX4PX7AEWvcH
j2MI3nvHKHC+28EXOZsjwAl+eQU4NXM9s1lvACLWsD0HR4gHDu2kGCP/ziBLpKtf
Mi59fgftVRZB7Lzro58SaRSTBOX0sW+RPn5lGf121IFLxaX2OBrTrk4jdIu0k9t+
5ptO819DI1mMUKp1a2mvU8aoPRl3cctzSWpbTw6LUYldl5GLh/g6tmcAzvnzVzz8
Z+Zc+fo+FPUgCgK60jWffXuEQoaaONHW0slDAC/P+athZCDRVnkXh6eYc3rJUq1a
8C4dN/QbD66rpScjdI9CWPTpn5lkXZpsQnWYYxvMat+eCxMGpeAQKN2SB4dtj7lV
xMGTt9T6UBtjy0Dlazea3NSb1RgLaa9GmTCM+72HN2xNyI5qnXczqb3NmSOZnUxJ
y4tB437Kkn419b3AJ7zDE5LVaLHoof5qh7JIQcYomBXfXWJ8JI7uWuZ22j/64IVF
zth8F4Z5RRPx6rnTAXxj8/DGPgW+VhxBwNgcOH27xNNx1TLHZOEIxdju5kObyVEy
bt2X5RVa8jvBgXoupijNQULsHJSdiNAHMx+e+aB4a0CefRqN0tnjDC528opAwG/2
G5NH/n0muI8t9sBdBF0RaSqWAWdwskSVq6KEG4pIHKBcUA3HbpnuZgVGNbAiip9W
I5LrIfL3Gzs9TNtdvqsz58Y9exaOz+FGeKj92LTPf/s+880rarOW/ftpsJkmk01d
BA2yWQG+DjrzOahKjo87IymoMtCUwpj3S6YGFdhcUH65ZVv1f4ltXW2LQelpIwJG
jigN+Ky73roNNKMCHGJeOfDjl8rrIB1xyVEcenLhEu9p0E/tS4J89qEh30L0HJzo
4iA5ZgqjE75pi4yn74sMxXK4Y37fA9r1PHQrGbgokMYj0cTeoAyjPNDVTEd23lCW
4DfPwl6AKP6eFB3H4O0Tq/dxp7bLjpQz4dMl9pXtH33iF4rpqCFJewb1gD1a1TuM
olQaIgBXZUyLT9o3qKb9Kq7OPlLuqJnTBQotvz5EKv344w0PVjY+dQQVBqkbnWS3
L6oVfc9K7CkETrmiXVSZpJ5iiTHVonbXjFWuuSsDkA0UPg0NMZ2cx1knX8mpJJdg
LjOOiX77t8qpVEYI6V4sw9JDa0IyOkzo2AabjC0RBnYtkoCxNgYxinME7Rv5Y0+j
/g9etTjGArmocDai1i6gaE32Zf/Qg5kKhTEFuvZNeUYCsuIWLI4fzzXjS+MYkvsX
Yse61rQN+3aEhiKefoZe0m5RwMBLsXqW/ejpdv5ql5uAzp4m2r+TgwvEBLiy6NjO
4S8h5u1lYRMqQX3OTui40Wol3ToZzrQWQCrGfeijoadHLqoyJPj5kMA9d2XTvvsT
nZ7e2cQO6MrasMZC7GRjwGQ2DENl4n+S8QsYjwQHluB7ucN6qzv4g180XmZSaR7K
ed5eE3Cn9aQjJ+DMTsA7pq5XiGW6GscVwOr7rDF3eGcmfPm5Y/bjgaFAcI9/LGE3
d5Y1OLvj+zGhhn0KlgXdf7/Z7LKNiHgnjBGVgt/2HGeHop3VT3fwcUcBaDrRhB6M
sgmcW4o9TpfUApPB0rvWds+k6h0EshnyXREj+01i4gSnoE3iYSEeVTKC6nWREQJg
hjj+JV9XOdJDyAfHgvu/C8vjbfO0jSBCXd2h70XJrHJ9o7K6jHGsXTz1CBvfZ5VH
ELtU9AwOUtSuVmzEAv6fvLfS/kU8T+8ja4pyaHs7h72OUhfn3ShP2r+scM0qgh0+
VxKVejHMYqe+JArOlrPr2s/vGh5qa1arm7VMRF4jlydc5Xh2CtNTNNAj4cGlEgRr
z6fNuGiZu/w7oJHsHkgHmBs4s0yB+g+WeJuIHVeBx8N5LLDicAHzXBZlWG6fQvX1
/ikiDK+wsIBypuX77U9+Vvk/4GVysgOuUdIymhO+ouPjx+N7Z6Eb8xFVKGZ3QPa8
6dPK/pFII9zvVpWxm3jhKEszgwLFhEG+/zYhiasbeWsan5/jnfkEX2TSOkEsw+pl
AZ0DH2etF2C7nWJ/8OVvFOOBGlu+q1fUwVm1HU5ODbBJeQw95Rw+kOE889NDOknY
6rky6rU/olF9a9i6rL96cVjumQ3DGec44dgtOM1SFh76ymcoiVnbjZyTZwWnd40O
8lFWTOA13/5V85qzceYpe+t0/Z3HpCdDv0cSsn92vLHVDO4vDwBwiDEj9hrwXYdX
CpzLho9FAh2H4Nul56FDon4LTy1fdQyXNZ3m5VoagypBqvsb0CRciaoMQIGBRiKY
hojidwrze7cWflizkz5zzy67aojmjfPioKkfMcygL/UEp82zmyApE6EE/f8J4G8B
5+kQSxx/oanRygniNHP5ixPz/PP2AURR/a89am3rIk5G18Bq+6hrCcoEkDtkhCWS
aOiQe9u2zGu9ImridBBxiddRvkCCLzwPKWSBO3FI/92hYW5gPDVsBhNbnUvXQfid
Kpe6ro/KyLX++KUtJko+kZ7h6EM7tnZwf3lmpWC2DdHtB46Ff4Bud7YKZjqBSR4V
bCgDvr+I7iLQgLufKru18ANxzgG5ey0lAAVZeG96ALpXpe6RBJt2MncDMaLjSB0x
4PCxosdQx0FPQbtbwKkw6BTx+tnuSJw60eZ77n51/Ywr4Fg4wq4czfccUM8+uAJl
ZeWVPkVyWu7DnVcarrcdVc2ruSl025vssCHqmfVcMDq0CmOJrVyYae2PAsrxGlRQ
jN26cASUyx5gk5ksmfoSqxf6uU9JQLp7+DYTM9LuWWvgVjo5RiJxkeieQb40SSTE
124bHa/01ve+O7f/qm8iASl7tn0hPKanlY2a2WnPM2/g8atTqnsOCKqfUgaR+H8z
+nC2iiC+egBGeRarno/EsGd+M/ey4QbAmIvfFERr+LfXJhm2LSiIX3W+z9qTxgcP
sc1IGlezInv9WXgCbZ+qriIjDLwwjjO2rOd5BZFDLSf2rNxw2CZFmCzuFEQIlg9g
/2iFKS9mcKpIkjuGyv2S2P7IvQ0sO7bmHNTslzwoD1y3SssQYh/iRNHsAwRquDEV
u63CroyNnoULKaVZE1e6lD55OzEwSl1Rccf50yGT5MelRXi5mw5Sh/jmys77Ba76
jNb0GtfY1/xrYpV1FXc5WvShOLoRogTGgA7YYh1RfeDLr38/zNJShAgglCEHwKQP
GaiSM0WTxM5lRT1FcNftF+eVjLeHGTaGKwxtGcZrQhxeHA8Z4/yPuKc9IP11spsr
RYcHsTT4JCPD/GHzElqCDh5RNS6DK7Gn3iKpohAPv7SQixlfKZVdbzgBJnRTFQWf
qNdgi/NPehZIljVSE0gWWUTbQ4ZbptQYwYVCEg5jCBa1h3QnUCAdKSuyW1pZzvKp
ecZ75pY7dpGQlxgDEwqa5PDt5HX8Tm/XB60EpsXXeLtgILoZo9RLKKY8TiLFtuBs
4Px+QezC9QN1b8HjErCk4LOON2ASrbwTEJgCBtFwZClonZovugxdKf2DSCQPERx3
UJ6z+I/Ptb1mQIBANSiAG2dFUAaqHEnksHBssSkMkmXljn5hAcZ0GQ3gq5kiUOyS
EzLndubv/3rfbBgCd2LRG/tNcBrB/V1Zb51r2yjvvmFUwC4J7A6HooCnPojRPYdH
QpFCwglBhJuiFP0MCjj4qeZXvfiYDh8tNqqPWWUnuyX7G1/mj02hmBABwvUCBaSs
Nrh4e+PQ/wLKPCZlpUPGhmsVIJ/0fMMv2ulNxT5qtQOvN04MwgK5Wo3IUiDDXreF
GUXgMTPqJhtI0fUso1ptydRuhoCv06Q316XDgbfrdXQSq6jpJMoOCwCucExX72fx
ezqAoP66wQ5Ro0U6gEr6ablIxMEIWcraarJKZo23ti/tIBpNWTOa8qiMkkm/L/GT
4GAcpRxxg/OMJVzNGtx2Gh2SBs7RcqgpbyRxW9wqKNN0738WLDpcSD7aGnqxm5ZZ
PEzbI203J/88LMUPkmWDM6zyjXF89HZB0aygIfMxMl2OrCiQx/q0AXuK1AKe37E7
r3jqGbM76preY+QTCyWw+NiPX3QtMbGitMAoEkUcQ16Dsxy15/XgsaS0YZmvXu2Z
g1MrG24O5e1jnIm7F8c1+EKWKqjbWB8d7T9N2QZ21UcPAJO00rBeVNUgmERNicFV
IKMzj7itdvU38TwJMQRMQ0dOUye49dysdpYn2hbED1dQOK2czrSc6nZGUp+8t7vz
BocFGlUtxkLe67REbnWdafMCaw/MSJ9YUbMh10aqJSTMWkmzhW+cYjSlyvhPPLZb
ZasVOtFnR1KLryRq6N3ErBlBT/SjO3ufsq13+swkdsNcF1Gq2fJEpdwLKprFzeC8
qaPwHmZ2i6RCORh0ubL13sZALnnr9tdnLIanFwmJKsStGTJoyGhBHIU9bmdBGS1U
jFwGRzituMNd13Qmhmj9YrXZXvWUPcg4uyhNiDYYRpfY9dycey/OGm8o2BFLk6O0
61H7w7I18uAkalfWXCQygatlj8v26461o7ZPpxlwrRkypEbAEj3k36tZBegqRvXf
NLZIqAgzNZvk8u3GfmV/QpKf3jTy5QImBmmvmVJqmZAXMZ6ZrW5CYWvAb+U5B6OO
8b8POz13mknNQGaHpR5qRZtifwtOsSO6Ne9n9RN5QFH7VH+FD92bSUVhltte5E/n
yv//B5L87J3gm9lMX1KwhT8FeCkvxK+IelvO4WMvmAdsiJ9ONTWxoWvp/zSnX0R7
JEX3Ag/WsKf0Jc6unE5tKyVEJIH6e81Fyx7wxbMtCjFLFkp8cm57b9BqMWfFpsdM
jgYVsKg9TiGD4+LDNCSXaYjj93cERF47VwJPaT1kodu92SPDtFedCDHZb7qub1gm
M1oNAj5HCiDj43EOTItwSSBmM+Es8FlbIXyXA3U0mWJH6utJIaeie6+qhwrVyeqt
GbLWXtrQj+cOoMlCDk5sBEaBhUJ61KrrOz+6wTFPQFF1/y65q7tfhN8GDqRPMair
WIKekoGVC8JLyp+RjGlU2yx2FxKwsdhsOoR3l63lWXTZV+4cjL/UWCJKbKvEE6r+
TbQzkkw3nKGC+3wu6zRmAMH6l/iJyHGDR9xtiC2Ic4jy2MR011w+eCeXl8+EO3xT
dit8QsxOyweqU+ocfWSqlQuZF57i+btob5SWK/tm7isUZChtVDF40afhUnLJvTRo
K4NAnKQ7M1NF2CEazKGhecROCSkWkhJcr9FBAejf2v0RBAzgfsKCuMNof225CGTP
2/VrMXWlj3TVrohr253PVEhwXLXkxsYYCkkvcH1aZoWCKZoiE+vQbz7iPBzF5rRT
rf2ikziUSMf/jMyLPRx7dyrwNtqNa+cXNTK5XSUb59sG9NoYopWfI2QNof0z6Lqo
S0xu7R2JJO6MJe86OZwSlZznyGoIf0TgkLA4OX+lKTjpqKaxwEgNCJHi7G+iTzRz
gEec2JgnC4cdiC1bnHoUY6PdchrhlG4IilLZoR4FIDIxAHcD3kIjOhiG37y3QPyn
PFlGbD4HOJeMtnSPQJDzPWGTuLKSrghEahQaTh+3yX/iDv7QLyZz7bfTY3EnKPdf
FnqLFqFG6k79tZGkVeUpnJHQqlQcBAzjfyrE69/R80QdTWD+RAXb+foGlOQDL8Y9
k5MRQ5jyp9SbN2NRVxyaG+K7LvkKF6hc0EQtVNwyueXMl4w7i59kRvNZ32XE0E5E
tdjPBxkeYuxgNt3cqiNWBc13gf0vv44uSY6h1bl/kxCTZYEwV+oS/b3xU2QHyhLS
FvSwQS751FLrGuubba+Vc2Oy55vGOgMMYh1yjc/nJn3U5Lm+74WZWpgpMqnql5vz
iOX+4YH5/BrXIdyFEtbeuN+B/iMUx406Y8b4M9nGfyQIMMdtt209I1TTBRPkaozu
KwH/HmbilufKjqbRnBzhqjX1IfMyq5Q23FyaxoXOWP+0AVXcaiWy9cigwoifh4/0
0RoKppEgd/aSZBTFW3yRBrVWz18rSon+pTPOwNddYiBZQk22R//2LvVo4QhYcAMK
BPpuGUb7ajyDK7Wc+awMpvuusAqNKkFCOYeiki7z9XilkyUuciu+NB9+3BjL3Muz
jZVaK/e3LVXu40rqm6qYlCoiwuB+7wgehAIwoq/hGYW7HFMlimc+xV+47F/LpijM
Ii8cJJQFZ2nu8Dp3MNq6Q+nZg7QaotCnuISuY1UuXkwAERhA4JOcez5F4O3ty2S/
NeBqTf0YaVTGXx07YRzTEnVtjBQv8MOsLsomJSV109DmKxjIRPQtv/zfYHgCVnwS
pRPEoMvGzf0QT+aF8ATbFnuu/jNd2SkICVXAyoPJthUDtnm07h1VoibKCCnFWma0
bSP5tl5zbi0hbIpcYZmWq+tZWQaiN1qcWeQRktzwsQMXR0QIHqtXy7OMbga3LIar
REzOM439La02JPV1gAKHfCOwXvtwrGQWS+Iv8rSpKqQ5tbdQVocm9o2xsE84sQat
HLnc16s8HaRLYcCFuPGnXYP+Nl1zorI3CiMt/cE7SDYNQdWyDCMl62creOdM+gtp
3DSa+mUO6FWQDHkWRj2McXvvi4BKJ1CCKzggZQ8H2NX+S9d3bli4P3BqNeR8tfqA
/MQsgKdRYgyv0iZgQ6+y4QXzgT4crL3d2doPtMg4x5TZ4iIqsbukE2VEa9DsEAnE
QWzvhN6rZEzzcx49gnwnU7rMoauntAh10Y9XFH/tXZv7n5C3zNRjbJGOcVV++igB
S9ZoH1PWzGT32+LXSCi471Q24PfFtR/ZKrowfCrFn/afzC6PtSGGAPzdyapIFS31
IehZnzsXsyHzpFbRCMkJCj+ay7AKIa19x0ySOHt2ztH8mN7ZVYE/MRR1LSfIK4G4
VIDPenLgyhWV32hpNy4wpBSu4/XbedMmrLG8zm4/3HyG8pqBU1zefesX1sNyNL2n
GRPpFo2pAXNB15TzmsK6kUAGFWiSkvcoxzlaPs/ReUGIsz6tSW5P6iZuZlynjdOa
881R6RIS9tng0PAzqdLNF6zTBrqLN06ZSi4CkdAgFUHPzkp+Ob5VcWgikxhmBT/l
m4kVt2PPYhoEsTiKnQjcsmtkVgA6BEU7zEWNcXewZpRY1HZowM01FhkNBNBQIjUC
HlanygKyJZjPfgIwupG52PJXmxOr1RP2EmcwHXvWRU7Rvz0tP4/XYOGRDi7pWXd3
Ln8/VqCQhmBJlWTHFL6BlselNdnABJqgHTzgh1v+LW9BHrncLxUy9jtJWEYHx5sP
xistq3GEJEjOCvx8o259G/5GBHDMtoKh2XtVeL0KyeX3qlt5jGRkcg0VIoTo7yV4
TZRDq1PuaCWjzrj+9jy1T9QhxOsjGeVOPGBHcwWRG6feZBqZKXhvl/JA5bdqGA8H
tks5xinkBmoExIoU4dkZROWeCCVry61QO0yQaQQnC5oCmRs4sVLvbgN2ej3KmZRg
z9ATTuV7RU6he4GqghbTu1WT3M6U+JPs3tcB1x3l/EtQe6Z5x+d8HSqUrWNyZgsM
C1tMin6I4X0JYGJKmAWwKnLgXGU/Y1Nlehb7sfp2C+95Q2o2IfaX36pVUhuQa9Zd
3YxyVFy2alUNPSPlRHeEfPE1yuVE0s7vc6mXrCjsEikQK95wCMn0955lj846tWbF
rFALliTihJWmEZqy2I5fHf61A6DoaVs8ejatO4lXdxPMveV0+rt/v19NvUAb5OgJ
GPElNsk2PnHtkHDTSOI9QQ09z8Cs4/8P2AZM6dUtLMNQCtWVx/v9SFIEJgLs12Pc
XL7VJySuuoA3EiEbXIcPWCfob+pjZtVPIWWIS6mFr83KAZmOinnyheK4gJ9viJVO
xebAJRHMAQCnLYcFFsnW0oLFJeMao6i48t5+uKw2+kET3UuYLspCQ+H2EkMvGoTF
8gUAknOr2/zd0J4l968oIizPqCWrBMyhpQLN8WeOw1YgNjTqulP80VIAzJ3+6om1
QWh1hqq0IMbqDsqicALWqOLvTDGwnFvuRwbY9XJD7so5KaZyTTc15jz/6oNvOJdY
7Ou7JeqvXAMzRmcZNEaAOJBX26EmrkNX+i5GtSRH+7Wy0wgJ3UuuFGz9wlYIGYCM
HxhI9/mTJgea1QxZGVGKI1N2lzGoqqyHhv5WKL3PiVAeC5JAHHnfi5A7v2VxxCoY
O5DhqP+LmoQUVx7vu9Hv7jcvx7nH3kXqnGdbJl8YctixQuRWxlIrudIIRX9InAnZ
2k0KQ/J4+XzomQZLGmserfln4kXhJCEYuOiFy9hElrr5Ca7OJBPw3IrWzXMiNvdM
fU5Z61DhKzcFgEZR+unpVX+/Iqv28HSjspMaw0zbH2RQCLhx0aG4cnJWEJ5ADCLB
5ADiEANPy55Ku+Ho9DeOCiA5LGXjs6slrHe0BPFq8L4s8NL7m/WA0rd0MXYkphtI
9i2r44b6n1Fh6i0Sr7cD2vm+vE9XbNYOv6tXBFc3lgKrPy0ZkMZIwomQzPxCVpwT
C9THVzRjNkVJuHXVjvKpwKX9heZSzq/PVMwYsFBq0RRLDLrVYlZi1xWKQCbGV5jM
utHLnafaWZuB5+dzfqOuMjIVqMFjL7vLhMPIy0Imb/fpVIazRVLfKOgfTOd5fYy3
eVQQpo/3zFfUd/ka5Oa5ly8xlEPb+kiIEQYVxDcyajisffkXRq5SgKl1FkL+Lvg9
lTvo8hu48sa+z4UdQsXxGRB36EsWU8329sLwepHnU7EQSufYBOR/uGDzxA4s1CJp
/Dmgn05bYwvvkiIKl//P5YLZ/XS88Hjwb/s11/h0BpOByyCUK5Z1ddT0VpbkOUpu
vJUMXXFNVOq9U5GVxF8/Wy3yBOhlo2wVkWAOvYNlHqJIGwOZe3VRD2yEDZsbEvHG
YlFi5VTNV9Yl6B6zFCFW/PchueUsNwaYJqrpXozhVPEyErK5mkILMKFSjPHCaF26
Y1SCB/BIOXlKN/01eXR2EUUEVnWNx5l8RYv3lUs0k5HVaPihYdsXis4/+Ny3TCZi
tdVK43UElVh3t5BsKIEgwDx/lT7mD9iJK9X4aZlz3c3Zv5awpp8P2dZ07oXJb6V/
HhPtkVWoPDeZBZCWk0qlUXOHVIDavFYwV09KfN1+yGVScfgWooFTpYcgjUAF/sWR
aftHubX+sTijIYXEgnbRTfWShQ1af3iRMnls2Yz68jA1btOcMRDSLck4iaUcsedy
xfA8PIBFEqwsgEYNvrSHBrdH8rsEJ5J18dN6L6hPTLrdi39CQCEO4QoOT5ShfDVL
nM+y58E2a7I8HDn+vqq5IDPdiCP43P9cWDS7e9xlMWzS2JDovsjgpdehzbPzfx6f
tNLmmq7pDKelYAyCvqw+378IpbnMBRIBvg+AvQHj5PeXgxR+WLAM5YL04nLifkAq
h21ByOHLd1cnWbcleTCbEEpRiK51w7A059+fNr4wjp73OU7iFvsY+tuVTxCqCyu3
4n8iW3hp0sBwzRRq643L+eQfWgx0rhF9rk3vYziQ5GDj+4TGqmNDnK66sIOKR1Fp
RivIx74hKQyMka3z5uWbTWqHUKfxjDy3bwsjd1+dJXVaIqem85qrYHg9O2i7TF44
JwOszPm/DV+8VpTMrGMur4e85IoJDrxftH+ZVsX936CnC4Ip1lLgd1Bi7qrHUw7T
WnpPsiZmSmCU6ZEzC0Q3gocdn/Pgc/Fp0/jbwtwm/iN6er4ttYS+SdrJC/C2oCmw
oMf5f7Dxit5uafnohS15eJamlTB/YMG6loV6isiRDMoz2Y8XSVQ61JoYHYi0bImn
CjLwY7SU07leFw/Bo3WLBPp3fB8QKVbgF21kKC+hWCLiDC6nGibcasVBREkA0tFP
7cj+rforFXWfwJnGCvFhvEGnoXt26zQzd773isxPkudRVDll/yBRL3HI0HhA3/eN
PIgxPg5Um/27EIpZUW4aJnZocnQtZhSqHNgPyXgkPGh7RfrX/gIKmqlt2NrfBxUV
9B6Lm7fNmyhIUSnnjFtatJrceO2xxxXttxtTYP+uojtJApgBijNurgrQw2gc+GI3
13mMQzZKD/VwBooi+Wj/henQW/Q5oeQUVmM6eU07yrRnHpSwU3EIE9GU+h0tsu/G
QK6S3IKE4gy+4OznNzIwu9bZeI4qmTn40W+jEaGF7darrXMYLyN4/04eMiC7rwdy
Zc4gLPNgC8WYizSIxwN4JIhMzMhMpAq/1OtucVgocFAk/WARuGApn8r5O6SSvkC4
jkliTgBkb8VIrFWe+O/QXovORn1N8bV1ezDXzAKcK7cyBUY+gJQmLbXIA8Woke9w
o6VsxWRsuaIhskR2a8ynuu19BRH74baKdpDbYJO6ngh5z1u134FfPWdX4Yv0zbM1
17lt0E+Mac/Met3dxT+V4NOnB9cTklDYUnBnS9YRpvyJktbF5fVJAB/FGgpN4Mew
H9mvucyPWGp9Mdy282Jyg9YSLIjF8L3RHucZsvlLjZeNuRP+/J0q3u4C+iAYmsV/
v1q09VeEQ00GLz/Q5H3ac7xQuxwxEp1OZWcKlRwHC681OfA9Cvtox33/ddzHVUYG
B+xPjHm3Ic1+fbyrmFMug2+0GR01vuNwpfYAwEwSCwD+j8Fu9Fr/NKG21KYb8QRJ
8LoNtzpaeYQRR7bjKAAE5OesfztA0d0RYBXTN66RBuCquP7ofyB4nAuyepD5waBU
ggAW7lR9H6MX95poQxQwIjGE6/eKzW8N9YomVJO0aClk3AYh43S8jiHYrhid5NEj
GwerFb/vnZoM9IR4QQlumzYkkrRNivytHo1jiqoCGAUHw47tY2hoiaG0CavmadBG
xJeByMAbN2gTdPIc8g0tN07zOpDF5eUqafI4v+dYCsB6C3shfYQY5PCho4Yi1d64
VMDcrjbD3NoAgyUkHWsj8bKMtr4aIhlBcjpF800v/TniI0B7qmLH13VUEJydvdrh
3P7EZ9+8In1zZ+Lnqad93EWgsBA4av898yDJEg/NXAD8bpnsF5CqIQho6oBEZhag
44yOdfUSpkV/fAd+2db3YAe/qTM2MfguIQVAaqMRU8KSxY+0ohpxTUnYF285JzGR
So3w+jYXZ7nKk0L3f1B/quBRxAb0LJlpiTbJBNAbMY0104DLE8b+CDDMvVCuD6eB
EZ2Q6xOhDzu6810fhh3+Uy51AynWQqhFHgqQacBSgBstsaNuZ8GMKyw7fh/32aHv
17Mym+jRq2oJx9WjJrOtmteuZzejknyMaNMnT9cRtJrBqhBTmSpI/8Dehf0ihvgI
R2LqBJazdy7OkAiJobvTac/06xfzQvFawrsD4lqHV8gfWph6raaR7HtOM80GVr00
kzAzHy5mbyVIatVQ9acIlE606i5eEKCCuinVSPtbqPKvzfNO77tJ5jdw+eldBiyi
k728afqo6HreghXDKQ8o/QlDbXSmywGnG8pE7W62hrOat2n7p8Oa0gF9deyBoThb
fi+oTZFk3yXlr+CoXWE00ERTI3lty5iPbo4WTySgcANLyHXxP+vdKrEaIMbhCF0E
kRXDKB2Ot4jlBLFZfYgpm1nubxRvckLrWhw6yNfPfO9eecT2Ged5lq95npQzvNbq
GUMoMf5id1MW7O/AZAeWQdl8DfBohImz8pyA46kc+qeJRAgC94OqIF4AQ1pCcoRH
d5Jw9yk2SqDw3k3W2Q4KlPfef/yJSjG3hnS/GTGmdKfPLtkpxSxNtZymxM6RylSG
SqbN/2dkZhw+H5ZZ9i93lqdy3YEPYY6/fIRiIddZcHVg4/Rrf8e9Q7kMEVTkuLQh
PQ40lTfc9Yu2PQT+pCWv/za8Bh4Iq15lcE8SSNE/CXb1UwGxKwB2vhcvtPqcKCDO
WAhoHE6yNWsRwZ/pb18ctMERv/0FVWDG82iYOIPow1oAdmsWGSUoqjCi5r+FotJD
FguoaJgpsYMWPw/z/U6na17aGzmIT2VyZt2L+xrY7jXcwcjhIX5w6nOoVrVHboYc
SSicoFGZdD9SSivCM7eVB5eV1MZH0qEGhOp6rLzzkb8+u073QOINmi2Qy/s68jI9
OLFfDV/ARLflHxUQMKRYN+EA2WIXRKKUoEh3tf+frAabPhG2XcdWegWiq4KqBCmW
hdwOTWGPSZBfzMvtsc9dhOBsZS7lKa28efHTfQdj20ypBX8wucT+Urp03QTnoS/g
4oKq19ALsT4WugBOZMx0Jx3eZUwtyUWINn0kgkbmJLQc4BGn6v9ZhdsxC3PyCcAY
FrOgvXsnXZoJ+kMAj/1YfjJKSzbE4sSPEL/iuWa8twWFbseWxWDkS2QcC/kIfrQn
pSXMApK5pOKRfPQFjkWbvLo/QjqKslWV6lLAZ3p3n8i6buKyt4g5/ekKUkiDV0BN
vKCIPMcCYFL2K+SKVc/C6pxdXKk8TP8aI1Xghuk8EvFXepd0ONBYUPfkP2WSjx57
Gx/FdK0iy4EJoiF9lGTbg9cZCAYKzc0fAnB+WcS0mpSsA0DX8gujKTf2HMvZ96nx
jnusP5V2H+VMHYWUzMCr4IMVivRUjOW1asTuw+ANwySwE2kv+jHWGf8TVo4LOg2k
j6vmBckBjHfAX2+dpZeVpdhZe7N4rjCIFAgkbVC4M7+XDgOK3ELFqXP8ck1WxP73
s+RivT7kvkHPvjD/7BBYqqMa/pcFm5lrnkC9iXirmOmUSuuZsveCSTThD5NR2g0I
kqSZs7qmvqkw3qnztYQ5fr90UkVYR86eSRCRLyZo+cqk9ouOQMBA3VNO1ci1bofV
Ru3LsqP3bk/SCbotJt+SKrwFPcM9NPFpD6afKbLI+iBLMUg0DLYpKI4+/Q/R4RBi
CEbTQcY3IkFuu64TLCYjeQKKaWaeKH0lxwIcxNB0yHtwz6GJxnLOw67hhYE9VYfY
OW4inWaHV9nRAdA+AiRGfN8esEicu/WKJT/ZR85t6eXEg+Y2Xps4++XSRcc/6Xpe
FZkbduTsmjiLbbFGUYuUT/Bddos1N+dbtfb2KZ2qMTl/sbYz2fRb60w9TAh0PtFA
z3T9scMM9Uv6+u+Jo23e9wx+ybiJpjuWGPeLDtQNtH84QHJxTwEzQoyw7RahsOfg
/CbeXOCqDyCw6H9as+fMyZ3Dqh/afXX0VzsjxmGB1P78UUqfPJBQtfH7OX9EOUYY
0arJBnxovPW5bnCddWANOvYYbdWg3/v4ZBXZnYn/Y1t2ywV1oE+AxQjstDXBnfXp
ia/R6Rbw3v2ZqnV9hwK0n7EBxST+EEdulmyxZjLJ/EjAFxWHt5lS/P+juDRXCAIT
K1IFweF0kRNCR2ITCLb4PoVMcLvfuxZAKxDP94hppr8+nWGdDADl78BDQiZYqtZU
yV2g2G0cF3Bh0XwHYGf3lRANqnEiJA/49p5Ycir5qzFL4NNjg+MlxDW34/WYa101
wqUjvm0ibrovc9D7UTcrQ0HduYYGQOrQ9/9blMLWRT9q/M17b7LD8MwpxLtC0VXJ
PGAELRjgLx+3JZuU36JsDpDlv8PDdlhNjJzIyBEOF8H2uCUZzv1cJ53/dShbjmq9
eSvLbkHPgSdu4BwaBaSkrC9Qy7XDJ/Q5+SrksSCBV+lS4zTSAHV9hMbDdMBqWWzA
xl7sp/q0JcySA04wh3v6lt0Lfe+PvGTMtIWDhUcPYvR+WfKfAQ+nPNR+fYf6BeYy
E+2h50q67EP5RVDX1iHBdXFSYAmLAODT3iKn4jh8+OslIds668xeFIirAtlnDzp/
2Ap7dKft9J7psx+cDJBHhXD0bHzCbgvYwXNmRI1pJvOnXwWj6E3JqzVS9piUimRC
ZTuFHLAW9T04xWMtdwFeRNPb3BEwwPBMA/ToVcc9WxqxzRjcTwuHO0JdOstn3GqK
uMtaPDh8q1BLM8Ulrk0bsmBuytAOLJ+kXtYAidS7LwrZqhvO1x5rnE1ssxOS/N+B
a1msHv5DkkPyvo0KacA6txXphkYNjbIzMcVtLoW2uDxE9K08ugUjjRdj6wyyuyA3
gXCAVeS9qDYg6FBioUobMrcGjcMYKaBuQ4PEiFjaoXJ20G3K/Lj0PfbiDQsrywYo
haObhvwE9dZFGYfV+WThx/1sRdYOXt/JW+0ETBNRtTfyirgAg2ysPyhBNV95cewn
0eZ4Iw/NF4wzSKgQedXT561IUkDEU0RJaA82qo+ZoSkeAGhgQwRd9AhFwFrhPzEk
tQq8ah5h3NGlFKbR+arkP71wn0o4hSdLUIScZC2BdwALRaRwlsqahQgSVeIEIyGI
PTTJwaXhyANBkT8PaFu/+OfwdOCebIqGX02oJc1UIRhYKgYjHq3YxvC3gFBt5Pen
SyU4zhQm/F0/RUmSFn+5vOmh7G7fV7PH2i0Ao+0Pel3TE2HrWyyl/X6lXSEZE4nI
fqTMUUI1UnelqFSAYMa3zFatb+f30pSWXf87zkXV9OUqZoLD4oG8RBo9k5h/LEPn
/LuPRtmfLHHVpfCt0VrpLHIvXssmT4q0qHUcIqoHyiEowlboEcw6H0jMEmkyGruQ
h3YewwzZCQvNxoaIe684qdHllPBUmsvHkzLow3jR6dklj6uHmzUmBNQ+O+g1WEbV
KDAqvAo70i0ApYwg6801w/9OPOXfZJu0Z0+T3PraK8xfGtJEGxMPivKuYhtrxDRc
6GDlNwoxg7wpOVZCHgDeojm6bn6raykTQLpVScfDwjwB4veIAQkgecJgbX9k7oOI
zw17Mj6zGJ1i6qq3eNInhMHKzcjPAK9LWQ7obUZYPtALuqqf2hs4bpaK4GC3l7/T
lTU4G9nOfyTxBM0vIlAaf3yC9Gu9sl6/fKbcP9OMLbfRI7nLKzWxm0LR0UhOrlGD
rmSGqFaiS7D2akIpHgpTUJ91WNYF4Vc/RPys/9oRaPi3+i7TKiOlbVGqAqRdNkrI
eC9XwOnXNuBwQR0lp+QnbrzkYxxU+cK8yzkzMdYscYxS/8fHfSfkoV1+oel3iiuD
xYctFu7qSsFYXDbID5OEl+Z3cnweUcCi7GdRGEUaKIndb3N1zU6+uMnyCLy3pdOE
/OCWQiVkxsM39BpTKNMGa819iPIEYMtBs9b0xEk8M2POB0EzUTYXRNZ6Z4dAAve4
jKqbmaKGOYErV4hr/k/rVAujNboQ8DewGhatOUEEdS1TCQVfxFdZgWpC2syZqR8W
FFYLuZNNiY/8mpkDEg9VJStI+Iq8b41xb56nBTIsD9Gj2Tw94tyGJduh0xHaCqZM
X1F56qeBF85ZDyBkYIEnpMIy3O/vYwAs4nOHJtUWn3fYazsQ6im8ZhFEKkSNdn48
xxx+R36ERH/UKjPENdunJhfrk0Mh3DjCOz46NodIuTosRxTrKv7XpuKP8vAqHRx+
DByTNaeZv0RKg6cSy6/FXaqO186/VuW0Sy67i+aduoUalp4zW/8kPraDlM4Rlqhn
2mVmxV1dztVRwaMwHc/HUYPBa1KI3sLzmir/T92APg1Y34QD+byJVw+TfFHXAKpP
o4vfI5PyCIs1QYx88CH81G/bEoRDOkpNKbV0/dt/YeBf0GBnCwprLIkNhxwiW9N/
dHVYyEna/5lUO7wJ60e0mQi2tIslpSUwONDrerbNPHxroDKH243+sY7/ThIF7Kok
NP73eXZlTuZCThqQSl5wzFKJzmvmDIpasjYX1U5Cng3h4PBnA3je/rVb0/qHTIiF
eOGUg3LQvKUd0mprNUEGjR/pnq3h2tAmYXTzMUBbKb3wOM/izSHsRrDGEP9lFOvB
Vxb++oACs8enf473VHC1Zpdb+LmLzHwa8+9CPdOtZodbjp1997rbUcCRoFcEn1YZ
Eo7n0nysPbIA8EMTfW0/2tLVn0OpR/qVzqTRkgVa9ahVNgvPbTT4CkVmco+gn6aM
7/ydD+8C2n6IGgDKTAuuP/48ivmNpMzwgqglwtJNGvwLZn9TBLNLJUzLlKwNrneY
BhVX1B8j0pgm3x6PeXKmOd8uDS3oPZWbHo0KarptJbaSbS5KZME3S+kyWmXI9600
XwbafKlA4N2k3ZLGqrqW8YlWXPWQLYdizpWhE5H3hGERObXidMPngcgXbijPXlax
czDPBh4o8HdY4c76foUU+kbs3JjVgW1Eux8GrBOEu4Xv/U1OFhgNo1+J2To4Z7FM
bXGJHTb9QOTkJB5CzY3IrehApBKarW4c9ebTDheq6Aqy/crQmLbfEXB1U7gjarLO
RCxBagsQalgjJqyvnmx820ABNelo6ar44C4wed2+Jdg9ZsCooiJSt5zWVvxrrbwN
jq5dj40l7AAN1SAWQ7/9FMFyeKnIu5v+uNAzoq+oOKsOAIcw3p6u9791N0vmY8FF
I+S0xoJWyxI6Ik5MXPrZqFHiNZ5XliWCWyQkb3D3an0QyEBc/NbKC9x2mEO2Tveh
grnvOKs2zLctiqb0TR9KmQt6Bi3n8XQzIyOFFRFpIrCruA9cGRRHpY1yMySRLJlD
Rb6PEVQRyDGx9NZyBMxX5+TU6DFpzM4tkeflsrQ0pC6Co/d5QpT5Xr3H9ySARxfw
asA8cIRL2oSnsEAloKFsk9j0f7/Uf25eN6+cgiD0fKVLm/dl5bWq+EAf6iiyFqer
XSPze7sBDRR9hDYp5PLAinJPvu5jxkfMetGJv6mSxkPTiXYyNHNTBMGsENdjr2re
bU3ZnDYoiJit6KqJcxcfVIQ4doC66Yh/iXifo/mhDjNV/gWMYxb0oMlRlnbRvMO3
7Npwrq5XkUQYVimWvLpZYBWq2Qj2sut3Q1UQclqeDztlBXzThulP5VW8siMoyV87
HltfTwwiOV+/xpZSPVzO+YXh+vPfgswKqgl52SHtmEFsz8JxfBkYMs+PxRaXRlwC
iNn4IoY802x92PgOT01hxpVXyArSSPEcyB3JmCsLVHsi/yAEHGW12a800b1QdM+N
OFueW/c0+gGibeItZXHlBc+Bhwtw7LxiXolcAptLN+T/eCfNC9sqWZ9IdR3Lg4Xi
78JCsOQJUgF9chQbcApB18BzznQflqzZNkiF2vBCcoCSKKonAeqLsnarGRnm4x2y
egs01CcBGy2wxNumZalrl2ThKaRdNjcYw1wln/Ey8qBVg3eObEiC6D1MLZwmMdJd
EVtG2Ut1wzCfoS/h3cqUFlk1pSJAJDECZSY2rVSbHO3BP2Xyr7wWCD/jvbuIDFvs
1cqCLg9NYCddSuvHlvuTEzg8lOzGx50+Qet8UbAhQTeBZVyTVSPcwAsbh3onuckt
mEiniotRGzEa7s1PrJ/BjDz4yq3SxkaTidIUjcuFTD6rFFU3v/twWOx1Se0+IhI5
M+4YAYamYcHzZ4T3nJFfAj7pM5uVseLJpoa159V9wGMQHoBLEaMXcJh//MaCo19B
AP9nBXRdsYe8YJ+LhhEJ50XbkqX7FZup1mLFi96qwAWm5uOfwkFKOHsxTYMiI7Z1
BpjmSmgA3rExseicGyc1yyF1k59YafCFU34gYMisBJOoKfhpa1tre7y0ABC+Ij44
q6AO8ifHw/x8ZqVVqqi7BGy06EBIDizbdCuMj126TsDR7sfk/vWzo477JZx/LLKn
xrrEfPJpNPJ70TRXZDbrPOGv5YGCRes9QnJJozFUl5i0r6yrEHp7amSG6wFJSi+i
unXDgkYuOPjN8bcterpff37zgeZV/8LJe9bX9wvEDWbwrEzcmjdtHyMxC8G5v7Qr
351SRN6IO7pqC/5hFwuOqnTgPRDNIc+I+60Nsj05Vinu2L4Mr6lBAa0kvgtyGjDx
DkHoIaeNtrBf6pShPmxdNrYCmU2/5RuunkVtOHokO8x2Mk7FuTQXBozWlxEu/Ivu
RqKScSo3WUxqhfCj4QZH67DNwq5bLlJUOAXCTS22/nUX1v3M+JeoDFHMnBWTC8oe
sr9lTVqY0g8RhRGqPvGd5UFBZTOYv1X/R8M0FqzwKsHHkPu5xrIHZQOyYN6SH84Q
sLCMStPDyhpDHiSxLtnyS8nMiEUPz/mAKRWhfz/ouS+LtfORMnYSM772z+Hd6b7z
1kzQGsXBFQ+xryuZGzV0QLwUcNMs4IK4bnOUHLPTuHFOuMf94pvY7w5kG9uIX8ps
M6pwfXwW0zB0xe8psRfG9N9NgdhZ/LBd8zqZ0VPGrRuRBjh0DfxatYxne/T+v+VD
Fo+e5ZlZ5w+ftvX4pxUY1wKuVvBQJELXyE6J9Eaq1J4a7Sb2gda0JF/y4nLNf5um
i1/BrdTNg32AqUWEnXZcIGAazDgJZEzVnLstJCNEN4E337AT6trmh+51lQgUX5G6
+g8XbpKSiXEVReqU3dhZwGRggVYxLTqejw/5E/520T3kS4SrrmU8swdf3tSBMZJb
L0seFchh/EhuO2CzCgWJAsW0h3zOyCByzOVT+KQh/3aXPT7TKcRKCUmaUw1Q0tyN
VKlSPol7KaEvgo+aEMBQcJRbuBDbogkQzWaIFOLVzR/1yFCBWF8HoHOIZBqqEKU6
iAXL0PF9tkNqBWHJhnESTAcrcubbLvIboMJCwH4NPR4rdAd0GjevH2MLV/usyuhs
Al3Ob23X9PIGDhlLdh0YwSynC8zqxryPvyyAPj7JTDyasekWXiNXuLz8xFwttToM
Lxv9Z0gyI3b14G0zfk9RZxpAXh7TwLsWDHz+HgdB0USse3tLu5ZxvxcQV7VRET+N
cQFZreYwki1XvQBc/vy6pCItLyEy/0jwRshNtlA+/M+kVH8i4uIMr2ZbJKlMsdax
l52YzM90hM6uamcOjuBu5l5DmJ/3K4C7kOPTAycQBmMewwMI1vHCpPr5ENIRKGog
AnJe5kPyVXmzEJikBjEvIJzylnuS7AIigbNjQAtW80DqDKaftd4sROjon6Y1BHut
kLp09yvXGAbuxfyPac8f9BRRxGRAUqJWZctgi72352/tjhQJhNNzMtavv1F/G+Pw
7TtjSskQ+T7CRwxaeuFV7mplRvIPDTlS8Z5sd5UaZwN3v5W+A9YnT0pHs8N/4ILx
9SCibeh72c7XThp9VFkxbg4fq8m9QibzXe7SguTBApczex/pX7HFuhogoQ+PS50m
uL1wJ7f61Pf6nbRaiFBYhHjE2sQ4cSwYZp+Qe5+fN3mtfEzpGELNV8S3ultvs883
p9MTnbP4DaBkPjJUp/LQ2F+jvJE581n4F+m7K4IXx8oukQxF9ckMtH/FpqokCDdE
FNPRm5YoUgmWCTkKjlVnbSSz4AklmbAX+78d9ngmcLU+je63dGiymeI27aoraiR5
XEh/XB41ac4FboaU9uKrYko+aENLI9eU7n2SCJYf2KGiPAH+cc2IgmFueKDjGkXA
DKceODS1yCJ6LZDuPYpPLJb/7QXwsO785MbYQ/c2ShqUT5FFV5yhC5aqZSRGjWvu
AZmKFn8e39wY6/UitBwGIJDvV402ji1MqTckWi/BsFQs6RpWrF3S4O4O3IXkWaVo
deJmVB3v5O0J/2DErFY6N7tesRkRWGY1shs4mEtbDFVFiMmjkVzAf3r3tK0BBj4p
jy5p7K8oKgLfMs8YWCBKXXKQJhRZySCaq0ewOm5ZceYZ7hwaUYR6Gzswl3D7bGcB
NaAeAtsNDNK9bdbLfasqvpTrMn4EXxhfOPjTl5F+bXGOoLLyENgUIqtzR6ZtJHbj
6HTrkBStBw4H9a01mHIN13sx61tYkWC37mWFo+9S6M4fQIIWqat3TNzxHs3ib0zD
ByyW8DMQEYR7w3OelgkVSLdQ9EnfXXFIAPZ/LQkAH5jhaJz+pyDMMqEKAVuJSRvT
F7B46ZwxH/E++ogs138bhukTT5EEK80QLzphRbubiWLJJMipoSeOA1ibCYhaYjBt
w24xsyRJm2n3b8ojll1BfM4rs0rzkTdOQGduUyHz2HtYZzyb6OZTLe0MXdv8LGim
InTyQivRx5r1JJilik463NkL7iw/0BW8uzD4zE6jgSsrJvG0GMnbCkhsEA+EhHvE
Qi9heshFrG/j733ImP6vwdZxEz+KRrkNTgKs/uc8BJLsiT6WwBlodENupKk0BIsN
F+GkBI1D7scOC7jUUe2F6Rd3ZR/n8QaCIVlalhFNct1NOt6nn6VxWdcKZQofA2UH
sDRyLxDJp0rRjj31A394rqnWnr3x7niXGiv4kH8a756Qia7MqWsoRkh283n/79PZ
ypyt+R8pF0GTL4zFfb4WufTjr7TWJ5pFKNnnOfFHcydNA4Zu/OSfT9e4L59vcip0
eLEcbrzA5Z/c8IFluPE0Nz73acrYLEoDpgq3p9h7kxAJE+SuV6KI8bW/cEBcFAAY
Uwls5f0a4BlkXq0QCbry1dkygXdNtYaADD/quZ7meVesi8pq23mP1+MHsHWYDzju
OqQ/1L/yJAaH5E5jOqIsZaWVEJuE04ahOWU7HASJQXATTv34xkmxoWLPxfJgRMts
aU40y//4lsxe8ickAzwMdG4i+9Coju8JH6pl3+xpUVC0WtQ2Ra3rQD60DTkTXIeG
a40UQFqBNC4f3AWwlg4fwBztiRvU1KZ6W8QHK8hpJM2X9fxJkr0DpERJ3OIiBMkU
wN6xG+VocJ0zF81V7g7CqF0vtQZsqlAxfSVQNgG1uC/iVsxSQEmmDsK57RVlwWdD
IehnnmKRjux4m7f+3MT57uLk+FdtdP7ynDp9y1mjB6MsJX3TsVqxXjE60eEGRJ+J
ED2cTzJKvvV4x87mm7a/3QsrfmTpHfxGIb7LZ1cx7qQnc1Ufsg/LhNZ/SVVsaeg7
UXDWiNwN7hkG/EWIP/0vDE74E7BGJcMM1vYON1Z33nsFu5DPxpvPvJrXFtI+9Yem
eV5zbd5A1lncb6EuvtAC+p2R7OfSizuszXxbHWHq2StgiPB1xd85r3YtHpIsiT/x
92NucvlM7qcTFe7Pn96D7yEskA7TlUyrahTBI+9N9DxaSZYnLeqwf/yzZf+RN9KB
q/q2EezXVeIeHKXzJrrT192nZHuZnSOoY/GBtsxsMXuBtfrvJXrVd9igsT7d/7hK
CB4vq0evm9EWFqoSIuhYGFobGPN1ACOvYiPU5aWGxkAy4OlMpZcNH0sVZiFRbQGu
4TePP6TtnalaoGkpWchF2SHmHaO61OHNsvzhxORGU/wst19iiU+paXAeAnsFtSZt
zg7vojh0XU3oQ0be1J0Dx8BYjRlPbt70z33Tvrf9++unx47eROvUgKEe/RaY7MRp
VZ+d1l0htv5RDX2ZOzIvpAzXROmyBmWKpOCcUEdhEIrS01pghzCnVp5eNUvciWFA
jDZjGzesynn7+t3B8KCjDnhDtoIUVwg5vjRYeFr7s0ceXU0NLx39Q/HaOtU2J8Pk
J/e9BEcB38mfVtDBFwbGiegG5ALMVznQQF8qr6m4VX0SrOG8KJhsZa2aZXBNCXFC
sWTDus4noorz3+EJjGuWuqhOGSLoUi1h28RHnwtTthSqDM/tQaIdvcO+niFve5R5
g1y2TGkgl9UP449i4KEb+BNtFXyeniHh+fvVPdqtA8Rcjvx6KbahjDDsnZWxLxBc
hgaV6wb06WP1xZZVATpH5n5CRsrqF1n8e19/3PUh92NpjErx6ziDzXfMnZskk3N1
9r9DynM+b8ZLAMlygkGeq5vImwmAT9iaJ9JDKFhSKWC5MnPcyBeEEJeom1/o8sao
ACZ8JTqjt5KVcQVabTgDeEiA8YqBeUtpMy1whDacxihgqqB23DjM4lQw7AmeURBF
VHSwv7286mP/+P+8FX2IpQDc8UmrpQbIRht/i4HTdr7iyWyMdTZX9dpazw4TQ3gh
0SGpOfG/XqPHk/M0/9rj8+UKl4EQgki1YQdrCsDMq1IaFFoPHfe1upnIuvDGMX0s
NLqyX4afq0r2D7XzYqejwQk0UiOntqAg7mvlywuuPdgCTlzt+HVDYrcd6k32By2Z
PkWkf2itphsmItrp51dhz4BTGzKpO21S14vvFP3SJc5i4DimncLtA6bs4PCvb9Q6
6UA9GzWnlUf7m9kQQrUo75vUDcMmIf7Xpweva2oVnatHIvagjvPASjleAKPYRHjc
RK+7cHfYLyu6BZLMpMfB1F+mvEZROjEC0aGpSx2yhfvLgtgQHtM4f83M0msW7H0d
2POM7ML5FrZGW4p9+Tb2cD+c5rYLzIPFf4cXc8NIGXAuyr5NL821Gh0Dlef8CHQj
E3y/uX550SpfY4O5558KyG/w/rJEg87d8gQ9P0knARwh4S9Bc12BK3f6BCzKFaK+
PbwGoO52WjZ+UWnM4EUzU/cggbWnRmrTQcCzWrnhcaanc9AiuQBwGz1dHSo/iM91
KLu2/0uuOa9YnNKEn/ZJWny7XB5lyiorJZS4qGOzLViNCdpAH6YnDdkkKD/5po97
u/d/iV3xn3FZZnA/H2MqHkNY5LxoJ5jmluwJVJjJA+UddMxGbBjldIGeNrNFrTjC
mNlzET5OAS8XCHFkI4e9J4QGqVYP6hVTi94wQzoBS58RGDktLAWm5LPb6Dhi4y7q
1iwBWuYtySdeXtQSIlumWKm5klqf2Vq4jrfIZkIjsoP0bKqNe+lF2utB+ostuLd1
HGWPivX/Xk/EZvIpERpe92B7DqZBl/Vt49Qxbrqo6xt5KRl08rEeqh8IjGDVK+K2
+GW0WTBM4wD+ONggrppd4WJGWiT8+ja4QP2MoV7Frn20ivSbKXTPrOAskV8Xzcj7
qNsBS0uger/a4oKm7RA8TB4L1V+P3PzFxKrup+71bnR2qEhL0/Lge3va/3lBx+kw
Rp9V4rq1PaJoqvgB/9tGv0IgUR3e+lcskAYfHnfzZZ1zWT17r3P3cdRk5CQ+Fc8W
Pk5oHFKRFLYMTkehe+ca13GWSGwgV3J403R10Yb/XCeJ8k2M+vC+iZ35wT+IHeUD
rO6DbYwJeozWlOVdRDjH3gESBYvwh0FhwcF9ID0cMn8GQWf7s1vkbkI3rJ3aMo65
/p9DCyLYc5jEo2KXoLzQ1uDR9dCj7pHDS22XuskySTVYkSI+Xks84dh+EBCoxU5y
4unGYnf5RkAv3AHe9IfvLUbyBoP7o8QeNZvI4cT4MK0iuTkBtj+yQ+s8L+lqExDE
W0v6X2wx18jd7myDeC+UQYEVXDlkpS4ZfE8xzBcFv1/FIZUGvw4weCKIr2JyR684
/zk3iT/9quDRn6g5b4C1O2jS92lY2T6l11ni2tw7iBtXB1qUg8aKyVUUDgWNOWpT
Sh4dkmQnLtIGj22fFpDljwLaEAAFL7mOxfNGUiuUA3NRQwaG985MRBY9QI5EBSkh
7O0DRpRqOywOzSxb9JUlaCRJeJlMGNNuBs5qrhMoYLA+vU8H8Ohz9Fp/pE5Pth/h
lC2tF0KqgJmaTXC7fADrDAGPegLTcKFEBtwET5vyQysozBOdsu7fe7vZ+3ezc3ro
3b0JQkFzZISSg/PQzLhdqyToEBWFApjwIr7B8aEL7uHj3hogGgwXZUIGk9UZn4DO
/q7vsbFsKxtXtI6SCI2LyC2P+6V5uSCbhdHahufz/AX1zQAITnGGr1MkfB0eZ1Ag
+ZJh+UQKpGVLXhzU0cvZoMJY5hntPa4a8oczWwKvqGzR0Yb7YT5Actz7DZZukn1T
nvUxm6xzhKdir0KU1DR1ceXvI1kX60Nb47t2zI+xWNZzu5ilo3uKZixnhNWRZ/kp
SXqQ2zQDx5RFLB7AjRSzlNLvt43OpoAjih1em57nest8tegrazoMEscO/IKBjiPg
JffOc/5KuMzI5G2jLRHR8L8o0QRBD5ia7vTxXgCgiRP/R/Faca5S8rKvJnJGxzgT
HI2x3lTEnpEu9J0QrGIVjScQhh99pfLLjyVFgDs03XzzNPyHeOwnZj6n2cTs2GmP
nQgSF765++cRIFZ9O0gv4ncelENUIiTNauGL/R5FhdH4mfxWpxkqG9fxzdJR3WV3
aBeUCvIIOjzcHtVGSiGqdcQuH7WJE/iyVVyc3W2FrWZNwq47nMfo83oAHOJC6n0h
03v44O6MTPPlb2N0z/UHBVH1mOenNoAmCCVVnMX+zVNLoijcww/XuWS44mybvIWN
QL+TQC7BI1+Q+Fq7rz6lK2R6a/MiiWUGzCRz8qdp9u4ZS3HYGgyQYR5qycZQ2fcZ
LI0NJ0BuzxVlhYBbTpxMziwLTwhmbqEX2fXFDkeFYBAikATxn9deHMjfrVKPHRu+
ROJT7eFD8mhWTOMPOfa1laKB+1fUdEsLEArv7afZyJMzGWndC1s+/TNoR6tm0JxT
fwb0Lwk5ZBC7fUtZTHZ3LoW91PkPkZhP9zuvoAm23DAMP3CepGw6BldZR0IW1zSA
/Dyn/ouYfxFd7JOZMiOgJ+Hx+yYp5mxIyDfdUJPSD2RfYoP/DjAsityj7eNSalr5
lFzqYcafrOW3qf3bB88mVTBQtN1aY3fQ/149agr5TnSSv3Gc6oC1bNsZKYufWXO0
fUpH48y5ISWlGOYo9IrLBSLAhvLtTKd9/aUyjW9/DrRsdPU6Pi7N1UZzVTw5WXXJ
okPSf4XVWcSlsYHILwUwf6cGPanCwKppVMrDGQvx6hnvqdl18qRaBHbQo2JtJtLL
lGinEidDOdtsy+Skx7X/tphZ2fyjdWP1mbeFRYO80gnKjjZKqOfdRAcx5OJucTnm
xQLB3uBf/4j0Hys2ZnJ7Y22xIybuDqUDQmlIybkUd3PjiCgKNfaEju/Zwxz9k6//
ubTkBfEa4dOLXwy0xN1dwG8BbRJ7idFz7M+X/TMy4R2Iv4ahmtpPwJkzb7raOKTE
QO/0pKl7ieb5RLaR95lkoMDdRVKJfIBT3UhkQp2o1WKZlIdDeJqQ3V4qSQ3/ANZE
LXFD8yQJY6uC+KiUuXXzrp0FVKR7boFrClQKYPWPQfIt+UQwXxv7IMXkrMyInDoR
A1PFA5rkatOa9542TTqtNaCq2d4NvjI5dAy4aFIw6cVTyOPZ7r/7jX1IFHAfvrhD
ZwL3tcyIQQ/o6Akl2aIiAK3+OoFSpFc+HIT0wYEVdvgRH8Eoh0QuY43iCkmbJDWR
MnKspYYhxz7/xPVrRdv+658kvLoMailR1fLzqoifzVv43s4+nodLAm2hhOBxstwu
dNi2tg3EpaogRPz91faVWyNCEEdyqFW0lU24tv6e59Z0U6BpyeGKrLxzvXw8Oxx/
J1tH2BJD8j7+au3apFsVEkrTWIJkuvSXwt68bT8/5hBze3RGuwNJowH/qz/oSVQZ
tVN8/olUekzZr+/WhAnz9MWN6JovAndMjPQdSlXatjiBp9JQbNdPTsoQz4gQNl7V
T+EakPkndEBeb8XBGVcvFnjuvnBxhVlkdXoYwXsESET7NZSTL7BH6lCgtL/yrLDk
yqHHNoUFJ2ogxIiea1yMn1KQe2vt8g0FLfA9TE2dPPQbGFZJ7PaWo0fb3YcxmEWd
xWpNS143lqLt8+fW7m8ryPMgTGqF+N3bUnj9CKlg1a8hCjriMRNE2j0WWnqbut+z
RRHOc3JrQ62egH2saZQJpGp6DxlsV2V6BDjQWhtETlM1q9T5hRmY3Y0aEV9bn0q3
VpRtFywxgFs8hFevy2rpzf+Akajzr9ycB5OUI79UeALaTYglt66S+WLDybaeiJnr
ysnXL5CRvxcdTq2iImJVD/gpgJCwCFzZOLzwM30CA0v6uTQucJ50uEksepcEIxB2
Dd5xAuaf5NPCs6/DDXJVJIsC1VQLJqacT++fsxc/7wFAYsGFa0wDP1AG5R+kUJ5B
if4iF3+qjjfBgvmuBX9c6A1yyKiD1ckdfdsF5eqfC30xs1c4J7iAyhQ8K2pvsHlY
xWEz7y+N4028ji4vD3tzxKfG8nOMUTDTs9j4V137tFKAAE4FWQonfmCeASZOS0wF
lzaCOQ+Wy4bjYMVBeI2xSCkgk01LVVkp2oj46TiErzM8EBdQksTtSN7wQ7pTRYKQ
+R85G3eIscnkvDg/U+RUzbtprFR/WVTRcdqGRVfcr6W+A71+uJp7kWdjktcAvk8S
pp4AzVKqKIVEA5Xkrq03QII7K/u7THLaDm566Cp7cBkCQ0vUrX/FSXPT568lRok4
b/cszINLa1GV9CPw0ZSnLjtzqZjjoO5xWz+HkeDLz4AsgLaJwyaVMRF0rEJirDBG
woBfHk6lIzjg8uCppB/gvyrG/6h2vquVU/nginbf1GIjk1up3bqf06LfaEmLUdS8
LvYwgg6zXZHeFGl4PaD90Amgm0ueAypOCZp56bq0yZ8sZfoJpeqVSLbqo7t+RuY2
GD/SKMjpJiL5qiDp8iXHM7ujGsaifbQQAPQDSNbhxfI3uivL5iMPgYsbzOVs1l/c
cst8SKTOGPtk1Mt0wmG3UEb3qt16Kq4ju283EWoTXuEJzEuI4Ff1IZWT2CEsVENc
H2zurDtDq2IeuYeSh/E7okCgbwc9TSAtisFqpPYQqD48c3A4mdw9P335dTTGsajh
JCdy113v11Y/Ob/E9Ffg1r0oV+NNBuD0TJWqX1atwA4ViyEHfp8if2ZD7h60cL30
J5BIGUJf4hH0dgRCSBV3C6ZsxsddIeVHfCqcbQ3c1Xxhgb0vF/3ZrWmhMkb4CzTC
/tLOPXZJWT2MihY69/ppTm/xTfnsMk6frp4pcPQo8Bk717vr1HtEyk4QYupdm2rl
iDSa0T2SmgYslLpEzHAElpVpNMcwHRTB8H1RmqNyp40Fm8SlHqVDyO/RGbXnhZJT
sgRVYqscnjFKnouITlyEyBwEJ/joiTePx1m77KjjJkQaibZp5zBWVnMKXdXExhlb
qcBP8MPI5/M79XKdp9blHlKRu9gyScM1Bl/VWt8+DvM0BWURNbBUStWkk2+tHpjQ
JZNsHUHr2v6panQra0WY09tcB3g1suHfbYZcbgTMv+wQ1EXim3vOumT4nFrRpoxN
nqxnMLdK94P18vQ6X4bCyYyuaO3ovI0uovAJf3YKKI5vJtrPpCciEPgCn/v4ucyX
xhuSVfE0uoPJ6SosrNEFaDMOn1AEeHWYW+W13CJcb2Xu+l/nCRiJ+S2y8SGiWvgm
V/myoKLrZITcapngFVOhYIN4rbPFbBUsoAckO1+HkiDnw41ntm64AiAfiqg+PXa8
MuuwCTwyxZzq1IBi49yUzrx3KM2bi66w37dxs/fC5scc6b1a7g7BbnRTtUovNbYP
w00OHv5a/1F+YiIXH7fpWXMN0Obbxry1kaKXSiP+UTtyjq7m1VP/Z3ZDMFon+7fc
zckk1sWpA2A2xQe/Ju5YlD5hQlQ7xjCXF3YBhfwy1Vrupv/FkR2vUeBsKaRGqPbT
XFao7OpSJ4sIEBV28IElSZmIunCLqTOmP9g6qW4IUINcDL00TbEG6+gR7cFjuDp7
20VIfwEkTzakqooH6j1iihLtMnR2dLsCyOAUYbBh5oXi8N+0i1e3aX2IZZM9YQ2+
n+nF0ILGB8hnkQ0AIX5zEPzqUZZOYHkyc+5oPMou1UR2WCookLPGkbAGl8ii550T
FArwdMeunAu0hfJrcZciNEoHANkUXBbHbN0JWwFegGBxYl4gSnNNfN6oZoXvHq4B
WzOSjiXbE7y7QxhXRJu9daxqQYBNLh7SzNcRMC3sHqI8X7mi49qxNthaW0t1Paje
LlnKNInZgNgkby8cl6u02sJQhnPq2j5P1l+2zgqIM46LsXILBk6+BlZTyOZK24jS
oppVer2w9vXIquqU8PXuUY/2mpu9rkq5sLbCR8pOFOtVrqJziuAgZ4JqJVHCPqnU
dRqxSSSN86sLxANoSyRER4UFLChoXa27NRazHB2fhF1pAegeFPyaxIcpiJahffs2
z9tE8x/GaA6Mby0JolvXZfCP5FXsKgZSJO83q2GQGR8m7lVUFJI9ZCj38+HDzh+1
B3JhK1qZY2qSdfo0j2vIpVKMAetcYr5LmBPfkqXAfObV3cegtpJ/CojKSWbp7LmM
leHwX6JEMpsiATx6eU4otqvuWf/Xd3CBSDw5Wq7klQolykApiqgYmvUn/RAwSzot
wT+1QfRmobUnn1i+Qzm3gvaFJmosPXFysW0+o/sVNtkMypGv+nAtmEOSX1a9uSOH
CHiCOrxxu9L3XQMEycWKIKNS0UxVV99E2UpEQYnfopZLu0nY2gVCg1NAVy7TJODn
adYwXUPkqrJLLYf8bn2G3bzMZuPnqrw6sw7ttJkvO/BSw2qwGauaCYt6/ug/9VnO
vpGHJJzJUDAUbhlyjMTcH5OBK3+aXWkCFpXX1XLpJcI88cd2Bpnv/d4QfYXD/Fdf
Tftzdf1jJTtH0JRFgDqLWYg/nFO11B6aEIuuwcnCt7o8ZTMgn/ZMmS3tSw3kHG8D
Pikx6SaFWOvbEQf3Ap0asIq3nFPTbITl1YJ6KdSH9JSS8eO+03Pa56UFzCkt30tu
cXSjGrqdLLa3RkWJv1p44pmVRYqKIO1a9O5RuMF4xJRknuA6MW3Z0Y6GLWoZOhbP
z6DfHFxYKM2pjmYdwWvDTYQEuoC4mx70T2QDUHgcYl+OZX6TKZkZVV6kN/gPpOAE
n1myUBMo4l8hZ1OLE18F+Mup1alVujDLeHLmEVN8g357f2PA580nA7Yxkop7GIUf
LMcdyBm5dE2i/Gm9gUpYrwJqvNZkFq4Exft2ibq1re3NE/J13AT5CFAKVtyVRsp4
sdVroZKNqZbXlPGYEM1XyynXCw74+sXj7lhW+/9TfcSDLvUVIpu2sk+ITf5JtLnu
nEwMDG4KMbaEKxPBZyRj9Pqj8GgYCuLzh6dNb8EA6CcfOaUMuWNIll8dkkshpoOX
ow65leCPZn4hd1WTcDlwsWafZGPXLLNZaAMSV3H6ivMJQuOLy1VjsbfY3uR7Tvm3
B7lWgaeNoJbN47NvBfdQHF3EqHlOyDo4/iOWHtt8jwNL6XUnseV/EgAxiqCFuxW6
eL8Ts4UFeXx5mB4ThazHq4Z8SYMtneqX4huARLRTbwqrw7D2hDt147BVr9HsVzEg
gf6cX5aXy4GLAvqJkULl8DPy4MWNGyL459tFWUtEcLsRKnFmOuvWeR76WamTdBwW
xHy4besy/9cyiQ678J2EIg0K86/lrdX0vKGj8u5mat0FE9Y6RKEYv0O9LxixqWrL
GzOknGFcb9hsECmlMUao/V8wtrwaaqdU+j/eVl+HLxVAs0GIHEzYcZHnOhVtcQQ2
jQMaIMhW5Qlt4XYSt/enHT+yqmi8MB01NtGVH+8OcFOeAg9CE3U0XjBhymv4k32P
5C21c4hJGOXpo1crK9T/5YL0sp8kbjLOj839kEe+vjfA/tBYlO0uv2YjchO+P5Ch
LZK2TOff3N7GimCrTjehCIycShxAW6W/+XgoyppIlhvPM6Pz8H/2BZA3mkOMDZpa
1PwSiBTLvHUVIlG6ivtv3N2akU3WRgZQSbLuUPIgybzstZF6HmnfPqk//BDdJukB
hcllUgg1xuRYmDfEjG7nHYlbvZ06V5ZIT+iFLPH5+xr/i6EsqcqtwSz3iNzNiEgl
bQz1gjMVj1eNfH6amb2bglVb+RRGfuasu9u6rHAYfzphKRGMaLbtG1dWcNNidp9J
Lkp1ZCyGS+OWskyVm/J3lYWFmBMv74xvDRuJZcPRo/f6QqTCf/tOfbmC01KgD5Sn
h9Sc1IyC4JJGC1qFAJ9zOZXFxOQiRWoPU9lXbSouCZKQjT2jeUWzAt2WfYQeplYr
2KJA2MxAaTmbS2NJNTO/YpFVri3ZecBtcz0B/fMqZ3MHPKcU/lNoWvO88r76/OGN
SR7z3QLvpGbpKKLDXxBMIxPsS/9J/g5W/Em462nKge48PB+C+Zmrww4uYPQfnEM9
X7veo6yQZNoIVQo/R32WrOh3EuEs3NQ2YKShAQCQhiq/PMIKajsUk9v0aiHSfwQF
j5+qSkLyJPo8qtSP7T4o3Qi2zh7lUMuL/mUVjKOl415S3E8yvsKKmwvEWR09JIP/
8DS+v+ldY6c/8BgKDjfBMdI6p3TstISkGQbYl+svD1vu7YeT4m6RvNdCicZkjozE
TMYEUDFA5BcItOo55uqU4qcE3ZJDoIN+BplftVxWKF8uHk9+5CFt1YKIQ9/yO9Ex
Mt+M5lwgvt2JHgtHLvK7MQbxHt688FhQPN9chL50UXe/uCofVk/C3NnBtw9LMHl3
nW6Ud2LUZHbdP7DYU/a1Z46qQbwtLFZVEFIY7E8kNM3wzubuBUbgdjpTnCnfHFqI
6oKU3nzOuAJO+AptpZ9N0wGyCc6B7sjjCOVMTyi597vDmKtp36Nl8PYXUlv/NpPR
Bg8t8Wrw5u4ULxOs7hVakgiOs2ThXt11shAT8sWx0K9ixypPzRiRKMznhkpNe6KW
jJ2d6qKWBbIMpaUvGh9qN+yzaUT/JoN+pQBz9fLD+irx/RPY2XhkWe9dLfymUbF8
x3lSgvVmuB5sBjzJGLReeIgbGVc4Zs9A2ZJkc/2Y5IExndZKOgA7qGej4mg/rhau
nsI7XcE9KU1YjzeKlytoXE40Bt/PpWpzMMo9A5DJpwkifToyqKYsNTHVSS9F98Vi
s81r03PUyVXb3N5kL/TcmNXo4li0QmeYsFhidAt6s0Oej4PZYvs+NLj5hOdBm269
7Ljx6+1+9co5p11tNpaIyerrhrz69A9ny4djIEzUPASywDODUO/Thx/Wj/QsuqkM
d8j6qIJK8RKFGab2X9F7ZH4NLypvGYSwCH75OVcKzrF8GVCR7cfjL4TvlO5xqQni
hA5t2vonybE55yJqkBapVzfH/s+kn8n75lcupKanELnutDW7ZYkmleiANoLRozTv
IUwC9nrgRTW9TRt2gqdpi1JGYKG2GaZ4kZBRHZ2eB/+hrmE/Yelv8PlmRA9tt2W6
CEfEwTjPOJFEFrrmLEawsjUYbRDVJMe+hoKMtIa2lGnAuUv3d8keZ3CpD5h3HIiq
0bLPvKfU31Qb9ePapGNmMcMwWHCuRSYwEV8Z9pTkOosHRtZREDXWzsusOUXtE/fv
RnmUna15wqAQXV7vQhjlqJ5XJVK9VWTAxAGSljXiTmEI5p0gCFzlR7Kf9uaFBegZ
EL4dwmIcTucbUPv2IJ0UvI0xYQbxwVWnpCwcb0u+mJy1AjwhgHDXRFcAnwrFetwx
PzVAixgiPb75yr6pr/NPe/J054Z7Tt9lcpstC17ZRfZLRLC/mYDv9QwcZReypJZD
xLS3gJoIldmnKx8dJIu0prel4I20wxudlDxMHPPzf4Lho02mRyfrN5Z0ByW/GYSm
JYvSHjXfaiDemXPh1z/0IKuyFt353z8l3Osfyh89I2RvchrxIandnY5gZzm9i0C5
3fUWBOaPGPNJ8PHSaqc4yhS9Nl+NjHGMufd4OE3491in556FaVjIocnnUbYk0YT0
hP8F1bXS1caeJj30semUPSDilompDPV2XCe/pLADT7eP2ZvmTgypQCkw6c1HUHEA
m0VJbz0ujic4ACSAVkAIioU/tSkChnGn9NfQaFZxPokt4dOl/LxKV7xNqncTgRzO
PTD8gFCgfbdHqppdBjmnLVOT5jwDg9tTjhEX38lpj2J49avSw/nnVB+IYhAdtz0i
ZAyqDn26MgAYp+ITEhH7LNzmNzc/fo2tm7cElTSvIy6M4RWOlgpy6VoXOzyn2Gxt
JroiWzsF9yT+/9QNZLpl1NLOT1B12QuuCIPOGHpWTAVwFIWhb4qtj2ZChLRGtxaW
6ZHd+qov90QsjCTG4LFpZ0zLoyWnrHCouzJSKgIxfoPxE2DpVhnHVf3SlkwpTdKb
bYz1oadc/fM/0yt1nXOk42IYvIc0yWZ+q9xh5pIyoK1Pf/Wfum3e5JPWtOo/B7fM
kwaeQXFf5UtZIA4Bg5CdKBp4YH9UOggo6eq1AL1bTNvRldxas/dUXdf36Bm7nJN4
u4chscCLSJQlp5RbwXkSDrUiOcugUMBCXlRMkEZ23RajWOUiW61VENFGhjXIAgqo
9He4SOpvBmxuEjIVZdfrXq1O6GZZNK5kwLPtmm5cmAhNdcPsgMpI5kzUOfBGJ67e
ZjVg1vGX8iaMdNsgIFfeK8W7k3TzZaPpIJjWI+cH3eRDHWjlCcYZbFwKdETw+CPA
vZCYjXlRKQQt7hRhu/NwfuWtPfkvkMlHKA/3qKuZkSqsIeq381c10Z19kEENujzD
Tgwg1g9zgg5ZLKu7lP57xw+oggnXAK8vfX29uJfp44SPWVSHriApCbHJv9ZtPUdp
1hFSAor+CMhtk/CbG8EdBHnmw4lMlDCrFi41zwD/G19hG9jRi5j9z3Jx5PMF1IoY
VZQPNJ6lpBsGvHLZJqOXxzd9/iWbvRvD7bEPLbeoziep3j7zP2WDCAKKDjVKW922
sv9jnNruJK2nhVPhHp0FmZtJ7gxLUsbPDLD+N+ahSxZ7bkrW/STU8gv3pV0b8fW4
ifTS2gfsnx0jxY2RFrZEltKH9ZMpgimkGU/E2JULfaNAqejXu6Un/Y/J1xZkQyub
UPazZZqknrD/g3AREFK2YNPd7Y98bc9kmIYOzk1mUhE/eyqcaDERV3ZkwBur3zpy
262XqKQoi+w/oOZJcgA4c74BZj5kKbbjuYMnYGYYmYPJHEUFThnNgFXkbkNUkLE2
G1TdTpnUR21M6gvQ1zPNrt+WN5Z6DLM3xE/HTKpChxj2ejM6zYYCnY8wi91QQjEm
z4O887FMpHaCznTc91LPRk4X5WeWcUWX9zUY/5+/UrYA542npwC67oQ4jYJywD3B
M5RLZ+NYUyVxT2yropI3D0sH5Zyt0Zn3nLzlOw/iHaFeYvbWP2WW5qy68G6tJCtP
RxxXlNoW8Qa+tDhuP7nwJsTAi0uZTiKJguCzuKBIkT3N2tCEKB94cEfEkEtzECiG
6PPHZ3nD2D1acBN6lh5+DyGc/PwodFPhGznXIrgx9khTN/rW5Df7AUMhAVR8mjJp
6InEmn49g3JhuXCdE4k/CwSt6OPU7XS5FfNIbWj9QKK/GszYb28sN4INcuwMFmkV
pM+StDmbv+zf7hzWOjYg/WYPQ+qvbzMKJK1oObsP4JpO2TSbHTlklGZM8hLjG7gJ
qWiJk7BblRxkMAAA3S/GW6VFTgCIGsPEr3fFGaP3Z01joJO8LcuHh4iBIq8cGant
11YnSbmvK5KssU/1HCsZpf94vYCCzW3/aDZFIwzaeJ1W+IxC7+2pce4TcEv5MVaB
Ef9IAGM41+kaBB4unk9pRKi7hdoaU0ZYtCgNc32RPEq4w1dQJkoIpLqaqL/b1U40
sAbQyXiMMwITDYcBLHnD41BdNNBqI+W+CYnKDLvq/8t0YvLcOYsSVczAx5UfPzzN
sA5Yer2zQU4bN9E7t6LXiDzoEvYyMlxzdGULcIEWn8lvFY2VGjVG9hRufE1AGmfx
d1Sux9R/5w8UbI3OqXP3VZ9BoK9If3FqGyD6FDaRu8jX6LDPXXZDz69oHV4WWk6N
hsGx/pN9DTcbjo7pSzXHNRCrrnypqKnwh7AXAGuJmkrhl3bjoFFLJW01lfPvERHR
6MWMseT1qMg6H9GkWKD96Jn8VzwR9EVPXWYCZlQgPf0sltpwvhwWrxmmSN6Xg8It
u56VXR/wgJ+nmbKu0beXwgYPfRgo0x81Z8l3TmoaLl2n0CeXQNNc5DrzbSYhWfXM
+gxdVOSm0sOgQ1FIxyUNUjx6ux/DGQMZYjVapgA1c3s6QO7g3SE4aZVxXW5aJZtD
OdJUQfaiHwcTRw3eGzbe5O1fLR4yv2OzTOk6f2/IKrVpTaNlKc7fxWUtF0QljcC+
UMyAej+pFlHgkWnIg8zeFeAiiI5AFwU+QMYWs6GjuP1jXyU/zqk/W3XFvntJgGjn
qspvIhjzDv8rgP1rNG9DGLXIUz7icduGnUSFNYgi6yrKI5Jg7BNpbWD9w1wl5EMp
wOuyOnvHnXGkD7tJFDunzD0JcZ5ckUOCo4AnZJdwRZQLGWk7x9aKOt7HHyufx8ss
JUTKyewz3icdeQOmHSUEzMalcmD4/f6PZ2dac71QMJl9q5rUCEzo6AabYmbRfNp8
fJWNe/I5j7DHLHvvXliajUARi934K9cHBFdX/iO3MfuyNfUP/mq6lTdEY8dKAP7j
BndQ5PO6dnHerJ6+NU1XWYEQR1mxF0j18nDQTtx4kFXwAigX32dr5V8+rYdpSfj5
7iHA4jNZONPwh+Hj+V/+I0MGp9JtpPrFdbhVMK+jGMIdMz5c9p4lgd8vY/TVeVl0
CQDngNGTRZnQYghK86JvU7a6t/+4CVwc+UQ6c3oPjTWIkY+wTHMik/No3PWfrXpe
TNsWRxP/2jYqvPkcD9i2uohfcX4Z6dVxMmLvzqsquLyr1MMb60i4DZP3gXcYymb8
fTewjmAjmTZkBRKdskJyzfGxDBgis73cZgDFCVGSel6wy3zy5TXjcOkD75sdABx+
Sb4JOz2mMdggz66GfG7VGZyZC5IbGdIkkl+953d0cc2LOuWr/EOEYPMKcvh5Ut7i
8GE72LfayaoW8dBm+Qur7feN9fh7rpkIPWMICk3v+1Cm0rJLD2/N2pQcxGEB3RG+
FrAGACmqfJx9nuwrrOOwPr9W7M4y8FwH8Jvu06NjFBAT/5j1dwajNndYO6IvWiOt
FQ3hMvDC6GMJBnP1/+Ct/AR+/gY+v3oslWBDhhOmpBrxZ6ht67OaSdIgPSryAot4
1YjUqgDi/beb8bl9/3sPGXmg3XR4N70Ib9p+8aDho/1NV/gYd8EHjZjYe3qpPJTs
iGx8Q/g1gpwOAm7+KkZ4ZgcRMWpZmH6jDHZIFgrAsNUZC9mzJTUylbpjIn0bIAKj
n/A9i9dySX95OUz6dEJvHR/NVJyDnANAAsdEuPDUdURPqEIHMpfCOGQGH/FhmTgH
zH/n7+ztQLkNx3kU87lHSD5xBhnFkFxYr0kRq4R6PdyK6eDyBkKSNdbN8AzCHB62
cypY0qOklxWqgqc9z/+CBhsJmcGw6ZWOyM1Wf2DymlELmc+O9/IuPs4N9JyIXg9Y
+oXzBLuY1Oy93dqu/+LTmUHTLFGKh3TdEaF0j/dfJFvBvQUgA6vjhefbiB++KXZx
mCfeRTq3r0KudRWwN+WN8xkw462sel2T3lB6X98Ko/G3xR2Yrdxv+ovGFZugLXpG
jYvTquA7c5i0eVvkxc+wxD14hy2DCvzYMm+2SDyimsq7vPTN3OzA5eoWJEe9gisN
OareqAShu9Rlqu26WS2zVdpdoFcyqsCfCDKwOoo0HdT1PcDV0pgopTKFFC5uGF2w
L80J6Q/YrKpLVyIXyFSNvYj5TFtb1eaYP2b0X0WAM5II6k33gK0/7RLwppWOfRd7
wTpx00IajMyoBJiiKcPpB46F0oapwqmRQDmtFENHlA+d8eoJcrIx6JnzoLuTk63j
9k2ywe8hntY1t3vVndZi24kn5RpkFxaiVLZxalDO/JfS4vVxHPFoVouF9THnCuv7
OGFlZ7ZReClF58ZPxMCAjBfmHDx/GM7Rgbth4iPoOaOUOfEEkJ4i77WDP4FmjyyL
1YsBw7iD11Mo94OZcE0YtWBHT3QaipmZ1JaM8qcHHuqyAnGJxFR7QfzJUxH31rfQ
80tf3/hOncwTwlKsXYgYavMphpIiP4GBHPqmXfH76tIn6qdkn/V/27o9GdcGrStG
MQ+hEmlue6AhUiTphyEeHIE8tST+Awes+FpaRXjb6i3gwc/NxDykKQrBsO7nGAc8
ekNyl6j/fl0iD5twxZSGaDvdnvICGIyRRTekKjbbOPVC4nV9gRyeSEN6QOgUA+0K
PFWktq3SJ/XaamKW+8tpkJeTqdWS8fisEje05aUqppGJaK9xgiN06bvWhcgDkIch
eeENxSgOwa9giwGG+U21keKxc+aZmoqQdC9S295XmHfcnGrYBM6EK0DnW9BpMlQ5
/sW35zPIkPl9/8xO553qQ0nr0wgMwc4qZmKmm6WQVmoR/7kIVum4Pxsi70D0//uL
5WGh1oGJ7FXpDhld2V94XXguW3VdyqOdaDKa2vXIUsLesdk/AMvH3QSBFi169qIE
Ii4iWx2pmFLWFFgIqzRt4unqNeqVO2oV7vY+F1zVE/SIDwnVG/JjziqG46Gwomy8
EoEnFyhmawSiz4XYpVE6zGaJuN+4HX8nv8q+tEiXK2czwW12SqFwJl4/KbsZR0tL
6Y8XT7LeH69PtiJssOgk72euju7MvNR7I4ATGXEZEoK5F4kpoFIH0/xw54pKCf5O
h+U7heV4JlduiPOge7FOebnQkfkqNAskvW4CbgKEG/PhQTdBDJG7UTFLF1OokZHm
adXaH6TIeCdLqSSfa4eljKVCgUkvh1HO5jmkOTQ+C1t3sCabRaDwsz83uvtuMqlg
zjRzolIOifuYRCPLFFPAQobuObEZ7eVky81zG3kRXP7pruApicAFJAM1rA8/m9Vw
ET/7h9ikaPUh8xA8dIWLmHaeDgFemxEmJbsFVB6/Y+W9te4O6rzgMfwizY2jGmIh
Os0rQhKJvsX7ARvqt1N2gLwNWjWwtvtWYmqyHFgPE5+odWRvHisbzdIZTfMH5xfN
pyblOpLKbBLjaGxZghPiXtqPXmzX1VbW4pYKOgVRavFeEvgfaGp02589kyeakIXl
2NbvscCzXlAzrcOHs3zA9aapOoiHzX6Zd2OsPfYVJq/uM5SmG021UWoCJ4Noct7O
JhNaJuTw54Hj36+ZfdCoMGdHg06ErZe9tho1aGq0nfuQYTO8iQWcJ3IcvdAp1LfN
LCrdZVORPKyi5mnaNL18z9fb2BPVzO5Z+b89Q2koKskpt2b3Z/bQTEk9BfKx/Gta
EYelkqbV9ROQTMHhKl1VHQxbPbRMOYciey9DBAtTplVaQ+i7ue+aT3nSKVPfgPaZ
Ww1e5OS+dMjunjufn6EDIV0n3+1uH4SF0LVREzr01dOeJlHgV8moG1qMP9KwAArV
6b1T6KdThDXgv16N1R9Afw93TJ7IJUOhL8k9WzioywJQ61xzGY5BJg5MNJ4Jn4KM
PKN+XbDblxwwBojm6FvQqWUuc3mUc49Vy6oRMf1mPMdbmtoxQT3YC1aTpCnn9x5Q
itRMr4qfloik19DYXnpJiKkD1Znk+oG/xsy6Jab7dJ/cXn+rXoDONKzffosD/uIG
F8+Brd2M5VhETjaKAXWNrYl+GWewCcQvORSlxQd9HRiM9bKl/R4MKgiWXaqcixEX
ib5lxjLAi3aQ3fsMWvV5fVO097IzodpZdvGHuvLJQ1jBARvBrL6okvd9+vhJCCdG
Zo609Y3AmN1lgLFyWX3NQCck9kCNL6oRXepHmHQ5vauXjZ7INnAXO6JNLQ0NDlo/
7XTkgftChWt5eHGhLih3bkz2Wt5tQJ39+/G8y18zBClYJz88gMdqegD25FTbGglp
e+Ljh8j7w9XWiioNvl97EJvjJd00dXJq0JqaKs+doe3NNJygpLh+XRZaab3Pgqda
DqUEkvVY9z/dB1cvYRnoSc8KoL1pVRkqTPcawd0r89ZTyRr4lo4JU9aYEVI46Ndw
OyDqtenReCkPMzGj2ESvutfxIFVEQKs6fvAnnNk2LrT8sopSLR8VldXLpL3etSMM
Ma4jsGLYWvZ77C4cDyq/LU3Dn91evsmsKF6ZxuwpBbI72HLEPXIQ85JhBWb3D+Hl
vJaj/fvZW1XcgXzXl1LuArLbs53NtEQUoxlAZP5SQ9G+9XmdxN5IfZ0QO8u15KRv
dyQ0cHuj0mBsmHPAKhBmWNOXaWRbHEVqfCWA5iK536xinsaD1dm/NH833HjrNYRG
NgRPz2WUIZnA+mRLSdC3U0xZPzCQnzmlsWDP+FodOEcCELWLZDqYohxE8UvKiiLE
0lZS+qO3x+mQZBSJe1/Zglsm6wgI8tJNU9Op5OpdyDW7Bnjhb5M+MNo1RpJcnTDo
X5ajQI25eIOtHLW+Kuf1KltEfGn8MQA4zsVdUed3N5IgLLiPrJSAGGJgpHXuam0c
xxZo/kZCo9Lx3FDGHlTCJ14lpkjeIUv1MoyTRCvC6oCk8+W61Tn2LDieemxA26uJ
tZkdXAE+C0eMtnXSEdKsXU844dVEZ3BEjQQWlZtcUQiz6+ea6zfeFlh4jMU32yH2
OWjlvc+DjxX4mqQJ9U987Y5EAJ3p6p/pDmV3S/ao+h1KIhYmVDq5eXOozWw7lbpx
MbMho9tY5auUMzMKW8pUPGUaltVOjPIycaW4QIXFjkhr2kwMoIGkaHCM5s8GnZmD
P5WbGK5NmL+kxusVuexemu/zceO3xCL82HkUnVM7v8YOukMcmJEAyxbvKjwfHOaT
cF+ian/cXGZaBpMFHvjtdYZgjWtE2Pdkr3VXlPzFlCYuDj4w3cCi69Ns7eRHklMb
ERCJupOde/PO2TNxFYAXXAOf9rXktH85N23xxAqvq6NclxzSAAnZIS0vsdY90Lye
uszlvftxrvPRuoFP1LBy5WhU1G6iMoFK5v+UATGN3iYs4LEaXpgwhITM0+AnczlE
4pwQqOr9YFYNguDNNRXr7PC8xNtWST/ihLyFScel4poWHNX6fnJK9XmbQylfjCVO
/huZBQSufdhw7FGJwhOXuM+M1Pa592OrjWpNcjxW4qOwrfvs0rmumwqykRSM0xWN
N1cjfxK5fyZvPYSSUI5HDeC68AjLPsdRPO2+YjvnssRAuweMi+41H9rlQdkAxJ2J
fSO8merL0sZ0PmKWOhOi0+Afn824bUVVs/8adbFYgdvfpkmkREwvmi5EvA6GMVFi
ELOTsuRcUmS4eGODNQom8HhTUii/B5ocV73lI7TuJbRJe2fKVA9WgSgOA53EXz6k
Ybuuca+2XtOPTzWUcaovb/TkF+QV6nyzSOnYP578D79JxnzHGIPrKyMXvxRdBlKX
8PjYJYFZfiGIsKH6xF4TyoDMEaVwhilemWImuj8fngSRNQVG8ghEFkWRVNFDgAse
AS2uOydkGhxqAX5vwovtxSaXVVEE/4144Iykyk2fIGfMH+229BfWa8xYlw8DhLfO
F2uA+AiIgUeQtBhgZtVATtjVnjCBJtWTiek6z79NfxX1zetjw+rwn9K2ouj26ziB
NNIgIrajUpsZqpY2BhEClsTY/7YWCiPWn9JzWEn6EGF/5spsoqEUmKYLVa/8P7Y8
V339+fMdNblu7PUGhC+Jto/d5K0T+MoAYG2Jq50LoDhKxOX8e6klkhIB8VZofEUA
PKQN5Fci9Xvq+sNGxKRvVVAWmJRgKLjtjolrUp+8NjoczXSYVRewQIToB1xcFCwD
EWMO305KQmVag5+rii6LNUXWkVWPcTyzAZT6bSK8naYkVNkpk8G4ro2iTkl/rKvn
kDG1XnC7zEKAX1Hu57awJpwiOMLdoZvsNwaWGdjatVW66FpaEIavX/kgsu/PKIuh
JmUZmlD6z2hdXbisBohey2V7nUAviSW3MIQ+52J3hy63d8Kyqr8CigdQxERb46Aj
sqQdRpcoDS+9DyaCqLiFEtJn41ehqb07nrpz7YOS19qzB9r10M/vzaEvsjiquoAy
s+aouOcVSBo1ooSPY3bR4wh89dW7WnHq1STyDEeRj2eac4QUkI2sKLdrOs6RnxW/
IuFK0F1yYjuSo+uduCBjwKbsZTL7SwE9092ywt5Ljv2aE9XFlzd/0vO1nohRyyva
83uYfDBNZI1wdKAj7aCJQREgS9SIvQVdy70RJL2qTVmM5IcJYpHE/qSOTPos3OvF
/hReRYVNgD4HSvJOozIgbqnDJZqo5GYDPHHUIZ8dw3shI7CO9+xRvffOb6Oc/dLM
KXELIGtrbF/ZwKQbSVKJIYHJLuMFBFO8UsX441reHqgXv87WC0fOV5/5IKMS8ENL
8ooXRC9hxcpPsHZeulLxHIge27shQG4tI7Stw9xomOLxSFL1OcLg6gX83BBipLyF
Tran9RlpX5GKr8H0D5u91RdlrxFN+3iAYG+igRO/L5KzOtRBIl1w+BbvmfC0oCQ/
vyRjgVnC6s1tCUewDwD6OyRLmZbLZ81h/ES+3e6TJ+YN/4ZrHoQ99KVHn078TRnd
pRTJLoGJn16hOafrkvlQB9TVRDmSkfmbB56CCwPUDnBy/vfni1V+AuInhjcNtZbn
b6B5v5uhB0Gpkp/ALZwJ4FmQuTCBiLjgiBUb2dZ2IFOpV58A4ns0hs/dww53T2DZ
n4ObMiS0tZBCKcO0eOCys40zOF+4BunRfbIkroSAXKmq3K4JFt83oungESo8IXYC
VYKsnuf9JymQ2alUzB00j7enHtJVG4QvWFMMjY2tkfTPzJZ3tVO3uPBl40mNMzLa
a0EkG+cr0ZScUvG1KHx0NfrhM448/Qu1HOnfhGcU/b/8B3lc+Bsr/4fKyMGPRlci
gfpHn+Q7hF/fsE+a1WicAJ8EBLksjONf3LCYEtfofxzTTTQ7fyXil1QofTeBJKwr
V2S7YhtOKdzLp1KKB1c8D6tit4dmWusbzVQgrW/gGYwzNcnHxY4z0CC+WmuuiOZr
Nsir/ECSyx/bXVmz99aq/yqwF9e7NSs0mjztj5hMRPkvK/5aLhY86zLy/+PErFpf
0tUHBFKtSJ/mPr2lYEf/rWAUUP5ioTiXDkf6PCgJGBhQplmXvY+0mBiVUvQ7V4Jo
lcxocZ6HTLaJ0lyqgpvESqWR7WRrAby0KOBIaanR+sQrD3iQnMNue4ZVgFixzt41
nEXut2a/Huf2Pcnz+WEi9/NHAs++leqrJbziobAcm2C/ZbV/bN4VbJWGMu9ju5nz
2BAvUKc6YNRAU3X+A03/dUqQtml/Nz7Taam6j6UxDw/mr1Zcw5eKbWOUgbmN7N3n
Gzlu5h9p/VVmA6kRXNVhK5NhTrGUiWCEOWbQ0g0/MEjGbTKgzuLoLwHwWOfE4MhX
L0XWhB00mchbt7+d7FFILCH8YiBBG/gpp6VU2zjPXc+1y01jjmsj6BzBou029dSO
2lSR2x7Qst7lRzPGKyJXXxJVxaJPgcIByi9MibIoke6MIwE3TTAGHZ9JLGSO3YNj
WhrCGGu0wVArkOx5rg6LBOJkn6V6aLHexgfEh8f9MJzGORqaKF363T3C1yvyph0/
9orL5fs8VweQV9ykJGZHPKClCDtUgrx24cu54ojQq56umriFt5W5RudTRPHW1f0Z
uRGHRVdv6JWjxZpeiAYcwleaASev6l2MPSv9M+FwLbtJMIalLnuxX+Fs4U2Bi3DW
oILivupVLRZsBTLce2kf6LqeB+RRFC1l8Gdg04DpXzEhtxm5Bu47Onm1OmsqzcmK
weML+xKHbccOf3ntqMjBT2YKsm9j0o+qPwq89S4EljcyfEK5LzW7tMxgwpDw9LGs
Aqe1xEC9/S/tbkpNexChWAlwXRdQ94OTSGViMa/SHLPN2cjAukUiEgr21tOUgNd2
CYIymAqIP6fYmORtIez6ZW1hkYKzF5JLnebJ9cCyJbY5r6jdu5zLLad7+KTAQbgs
T6tj0vyt1alVRG9FSSBK/B8XHnxXXwTpN+RIq+ZfoRYJD3ImOT66I6vJi6XO8hl+
2dx+qMHWxXF5CF+CuHzP6vDbzaL6mQjh3743AaY4ju4pK7MU7QU2YXpcO7OfyP0q
cvvmlXq3UozWtQMiMmcojsqbsAnA3WA7ognY+WvHgOsaiwOKjnpsBHzgGmBXiwVp
XHQhnEHluRH8oCxdE7K/cDJVtcYwgyeBe32e1HccINqeceu6PWGEVJDxgtBETFnH
Df5IZjbNCF0MGC0tojndUan+XSldrIBJyU2pRLFT+SvnywX41x3FJo4+M2VPNWzF
zAT7UnTQaNJh+H23jcvBsrr8KDhyQyl6fUgAmUzJ+ihedDK3m7o/Ezz2qpU+qxx5
fO739/SJ+kJsnD5JYUIzQ2CoO7PCoY4/SGUoD3nWAnlxOsyLqImcSkbNe1U1GwKR
STh1CLIEdxulbQeRmGwodkiYuj+TquCnCVlOBavnPFKktrpIMjIbkIiYWGTckRCb
7xfOLIJF6IJBFkq130qslmz+ZYkJpZl2LcYHjUFecve1pPG7oOimcjtp8A9kkNGa
a3Wdz49NrrRncY1r6hTSm6Qis2ZQpm7l6ASX6I12pr6tHYdlB/P2G53dEV0zm53v
JOz3+8JO+8y7e2gxRUXKMAykArVVOy2pdSQ858uFS7VfjeuFxDXKvkR3Ebo7qiE9
GkSXInLRNOtcY7L+qvfXYyecjgwMsrcXNFOptAuZjxoZIz9CIQE4fjDXCFA7Ek3P
bsihWXZVnoQEPIa9/26FAkSq/JnR8YEnLdLf/wg14HWeWCHn/gNUczATwB/3Ifv8
/UJ06WJ91i6ethbTgPpaQ+qgT9sZIws9j9uQN9K/ubK0ysaR5qGQhe2gY5iZavDE
NRP0+GI+bafJAkr2b4buTde1F8WInzEhu/eq2wMdOR+nOjttUlxFlGCZZ5cDvn3f
93hRRUf5+VgtywI2LEICdCddvqhvCTaggZmej/+EQdIuJKxjez9QzkAPZG2R58I5
8yh6kGBXZBuxl79GpcbAcUsgwb/7oNcJzmCQ8kgansnezXpiBjYmf4GqSPSmbfNb
2uh7XzxOiUEm+K0RlTvs/g3zGwBBKWgRjUHiTOSe8xs/NA/Knb0ZrUFiuDKtaEdG
KKFTM4yQMj/QzMXRkD8I9mHSsv7rKma4Hbe6osL/+vu+JazlCUrV7h3yUy7hbGQE
prjnOceqcTeo7lqWZzOCirC92vJX2e5tpvTWB8iOzAWrooiA9VU38Z3jgL5T1Mqy
RB0LxveoK+FGvX3jZucPwMsBy+td8FUlLF+C6ttnJ3H89KCMNbkVvzyL6bWqHP/B
KKtiFhX2qViDKPAfWIp6q3JqvgedwTN3ckfrA7BCIyOgfKhX8YCpc5S5iUYm5RXF
ljFLzffIHxULi5TgbdtG1Fkmcu+hOyvNcA1vokO9xVpS70BaoIxjzTYRhiRF2m9i
tsSQAaIRxGBfzdoDEa9+YED6f2y0urVVodKLPbb2MCdYg5Fh2HDyFl0LqQsyig/7
EYUKw87Dac/0mHGpqv/3Ix4xjUMIEzBwlAnkrelnKmmy6SO8rchVodMiYLFGnXc7
/Cdm2/3RxV+pPrSplRanP7qhl0OR0vtXg5msj5LIYCAEQrgwcwpf2yq/fZOPZlOX
sY2ePGB3lVSPMX+lOSmDK+bWGPB/chFXxd8aax0Laamubo1C9qP6u1zg5Ahj353T
c39482UnMjzepUm18/1q0pSMNtHrsVQECdHFlGp5wEcCCOUDibWM6mEodLjIHtf9
RRPpz2ZYdJiTfQUxPd6Dg7blNdTTEq35FCQoSsXD9dYSRv0zTHDnd/g0LBGNO0iq
4DCbIhCdF3eRqQRxHDYpwX8qqk8/cEF/sJPJNO6kckFDozejdGoivFXdYxtfHsmR
+WnMbUtLgKesHhJOfMtsfZ2SyS5BZ2/1q5mgrWmqBnOWHoxKH/cWCOzwCnrZNMQc
98LhyfhqBgz5xmVoGAnO3qFpHII9G9I556yb7ky6QFzHzKOAMsDqzsZi5kw66Ryv
/V1GswRZzkUbmEJki3j9kcQxO0BwdRl4Q4FAuT5fyfbv7DjfnA6t+vjeTEs49u2T
Es5opl69Zx9MZelR+YaCRPAGXWufOVooxpzHIKKDUHIGo2YXiGEj1OtqlbdN2/TL
dCD8PJUfIgkqkvugBOkao6FBk7FOeujvrWiU/m0/cA2hyHwFCdl8Fj6XDs0DZU03
w1mlpflH7farSijdK6Gp34T+m2hH2B5JJQU+GDMysuyqChDT4ofaZCn3SoewGNd5
+NTh5GuKmH3N88PmXS1L/fYqPF6TcP3j76pdawd7bz/7K6+WXp/JyGe/3hYAXMZr
VVayCOBFXy7k29vpe3T3q63BrkyY60BJSSFOzwCWMDIroB4ftGDQ2njVjX84ecDq
U/mwxJeuI4dWz+3upfHu8L5rd+9Y+6L23S2GTRqfVde9rP471gGXXGxnyaoS2Ry5
J6zWvP+85CFsX01C6iiZy9zhFvy5XmcEzsNaYye9iRFhY25mbRGhI0bIjrEMwaFw
zBChkHg+92EMKlkmvudAuBQsvU/bxOaKvWy07VMmZ2UWaS6nzeYqvZaJ8GG0uZJj
l/nloLcCKYIm4kEeU/hjmaU7Xb251/k5zF2uH7kuztxvUC76wDrd3Zv5WI8LHxla
QQtzyTZoiGt9BR1ySAx0bhgkFy4+aqpxuhK5zdCbRznrAxJiB7NmceOSa5NjFkjR
2UHYIcN1O2oyjNs+ouMt/ckpmfqDsXmO+U0xRVcDB2EhXb3iHwHi6YRjtsbWcY4O
5xpCcE3h+3SYoy2x7tjOeFCAusjlCz8Jdqi7Lbc96p3qSD968W5Yhmx7hwZvGSFE
cA3p+ULG3BbGTm8faxwuCvF3Qo4wEp3pAYG7FcGi38WQxrd8RStyerZLCDdC4eej
O0eIXwl1c8DWcYaEUaecX90OhI+z7pmn2MHTK8zl307CPK24+/ufz6J736S3ACO/
cYnVBGtoxhmn/nmsW+3SMMfySsihLo9NCpi5D9qR2WsOv+SKdwewYdXJXoe3BRBb
nb4VelxC4TYb/ivPLAzYu8/t6udWXxr+lfCf3epOS/DXSEedF2wuz80SrCKWksyy
RyEZPaRAMa/R7CEWqxqqn6O3s1nG6VubBAUZj6WUhdhUP8hgFIy0LqGbTEwDc+3V
Xb2PbTtFu+WBu3v0gcwkX8sKBwzCSbFVQcrm8UeGatuEFUvVj6Vc+FogNXd7KYg2
yW1IzQD5wCPls0MngXHeBZepaF3HszHCUyNvf7whZntdJ0HMjqz3SbgT6cJHWRn4
kulXL/zc+6Th/b/nLKugKaDQZYEulqXk1uKsdJwfb3qkyKSt1qUlsCyvhC9v5KNx
gg5J0dF3RiXAC52HNB6t4uz6Tc1DfwvGLQ5y3keQPDmIXgt+yiV+L+osf9Ey8RQ/
ikzHWV5Ibh/ooRtFm6hVVKTzi4f6hIL+imwhZlxRTetDFUm6bd86+arkEDkMZ6I5
qBW362zlRapQpKBQSraem75Bnn1jPaECHrYo82X5pNYZbmHZBxuBCUSn3R/RuBuU
BXUnBYVX7GGyr2Dk5hrDiSEU7IsdFpP2X8+HgIwzuqAYQBf4NDeewZWhvWKZZDBA
h4mhpq6k0HqF3kfPqDqJ5d8Umj7quunfp2gQZ8kFdsZgtrciVZjmx46/26vJsHGf
3gF82Rb6UKdnGwJZODMYZpy9CW6TEQsLC3xJxEnBRxrUhew+yXaF+0X8kzz876nr
bAV2rDJAeUbdat5D0Rbuxf8hV0K/Gc8c7JlXpl4plYpzyYz74DOQB1eA4Mfs85CV
BaYXbyH+Rb+kdL+s1s08Ktvrq4HfHDLVezW31KeCDa/uudc7OlTKJqtYg/nXc0Qn
etRsHoTQ7sueGbKPVNSc3GJ33IJFm/TxZoORn40RCWWhUq9QAP/8NQF0JHXm75WT
k0DX2AOjqtGyJwBz35Ql7vQNA/LD5AYO1vc0OQInFAwR98vae/4qDA3dAp+l9p+q
XZUrpBSulOcwVdfwr1qUTIJu1UJPqg47xFee1Gqm8VMqPSdfqkIpN+xJtuPBIXh8
OLTUPIBLJHsSmDY0ja9MBpN726Ee7wRnVvYo4/+KQEvoE0i8V3kk30UT5fZMeAHn
9CiOSgehFX3XsOMJKhC7ydHlpidBwSZNncT/kICnditz6ygiUly7gB0Aa4d3hXar
rCso2VRHvviEpELWr1Zd5x8tqgAL9qRFJsymK7I7qAuycXwU9ffGUUMLHHrrwBMj
mXtEh9bBV0kNN3GHTDF4ZE1Rg/DmTIWNMPlf85PUbEaaUYOPjPsLgAyuzoLQTtb1
KSP7VJ+crDQGMq/6JJUC0/bk3rd9VJLaqR8e0Ex9ZyApoK7CXgbVC+LxGV9n4cIo
oUPboL4vI/flndbOps8AVxOoxg/aZpwmE09r3SMLR9Bj8+Hzjbx+v1jH1FdDwEAf
pRACNXWV5dFRAFIlFgq3APrMLsdBCofIVvdByvZhk6EN3qJTEP94JDc8LHiUtcsR
bG24f7QIcPXM71PVkhEuFpKqO3C+vZTh8faEESDPOT2pm/wMoHGi2XSmtmulpIy/
wbvJZYDYjKdtswGR5BaeT3cUWmzzsU6FOGULDAOmjkOkdKdFwY2eSwCzXTR6Xm7/
IAdvzXjBdrCj/kNp1arLwVDDKgan7eaps95AXWUV/JQb65+QxMSYWLwramFR+e/B
u24fBCiiL5xFxpMPYbx5zKNYEI1VDrb2J8orJe2wYJ8siF8TJr+MV+H8AFn12TMw
AUo6611g+IAOyQ+FA0/qKgv6EbLjtQtCIFROpfwxbJ1vlEuluy+nQkg7vaQKTbBj
PLHLbM4jCbJ8QWeVvKi5tiDuXVnBNgG1eySU++g6jwMLBuTpc8lDNgYw/JwaMv6k
8WHhBBBw/d8E00i9Wz/0BU5ADVVArfKEJp2PaDX8OVRe9lqqsqpn2pu6qW9fXYQd
oqJ+/BQElr//vIoWVx7Lbzd6aNIkaBMWW8AitFhLZTBJvGOmtNQEc/W8gATmgPXv
SijuZQhM/hsjJlg0aI0jN7wgIu0f9bM/lqXk/84euczc8Ugx3xbgEucSz9VwJrc0
aH6tHBWBPunGJ5qRBVEfHdIByStgaDVdj525qLWKt4tdDRAYb1YX9lCUtLsZ2mVI
QfsHVyKOdPlIAedQ3i2C2cV9f0HfwElP7jfXaefywpXA7bk3kjb2jn02byAf7jeX
sBiGbi16YoH9De+nYn2ugSYdOj5CJ/xjKr0LdK/ajoL2pAnATpFc0bzXIjRDK66Y
YQlYtLLc4n/JCFh6ygbrFqI9OPoDfr8TyRN73B89sA6d7EBBUMNb1AZpQof58RKF
TwWVO7koL6tCYtI21NfpAEKqloiFV8yVcNtBR/bl2OwTqoxjhfBijz+rUnWywnMy
tj+XPGv3rqm6ChabsZ/TqqtVxihlYs4X1Xp+KL1L9M9PoNmiOnJkESqifvZ93pbd
22l1IrdSktOyvel11EzrZ5TZQAkDOLMO1AwPibLkM0Z1ScAdQTfwbS6mdR8Uups7
g07T5LraCo2LeFMyTurHspHEMoptLYY9SoobAOzdjLtcqU1cc2ZnKZu0vFzkR6Vl
kQ8+CMeGMRHG0WA2Spz6oUDh7DVxFKuLkYNql2Crx8iy9ZoaGXlgxNCXtU8m6c/5
gNVitLv5S8w63s3jufoqJGFocH9pvxs8rxH8wHeKDB13Oij5djpd/UMKgScyaCat
iVR6wEYqr1RTqGcSf8aPGE2wJLali+VbBz11LJJXMxv4nh62UUjUP5c7HE2CAIAy
f78NB/PmFhZ3kbw1YkkdGYNNEyMONIEgs2jzUL4QqJTw+q0f28qoTICHsqOtrlPv
xoplNYfoj1+bcoPvBx66d1aicJmihwJSJPlyTvor+6MCB2qi5WFpJh3SS0jxF9RK
Xdxa3GdxPD425oTzAVf2O9RC6phJrWxs8mmyKGOYU1zAz9txPOFaGd1Ra8Ig6QIL
RCRyX/yLzny41PR/8fsXYSgSGK18QODBfuXQo/HEDY/NCuJgV2hQArbJAHzxcBla
0Z3BI11+cIOUpgQVdca6N99YTVGSkFNGvpbt96+Y1k7bEfmrGgaz9idQDHNbC/YY
mAM/4bTP5ml6lpar0eZUwN9KS/8vrCN53vLmCRgrOMJ5yBpQducKafbsofVovXiX
ci/k5AaONe5f5aBVicLGkuQYRWm6e1/Gsx1zhz9LQdC1kjOqZSEcrqSvvcUCPmBZ
Xl8xuCjWwl66yzTJJYqteDcsN7Z6TEnYkpwwTkhkWHCe2O4pAGka0E25EsGibZWS
QoxcxMyoDi9n7CWGH/Kawgr+aB3t6SQ9ySG/l+apPkhN/fx1Wfn5c4bPBc8fR+dr
EwLCLuV0OhxF64U3ufz1xeNi6FkjU8UN7gK+xel6QmCWQ44Sqcvul+6zKWVFPvHi
NEJrlnWmYZvA59K36CU9kEFizp7PktkAO6nNAlxfRpIfaDZ3Z0PB3sHIsSRww/Z6
MOjmRIxjwmUFcgsl5Anmn49jWP8uLGDv2WStYKn3tL23zoD7hqhpIkghMpLfGiO8
j+5BDNAeVfLr7/IHDNWkNXqAY3R2Q31Cc1iT+iIzRhkDk05qeWK/HArmnBwrlxiK
G5QSUjsKiqVH25kZMiVQagkU1syJz31kDZ2xA34DAHs6zrOA15RH7ydVvFTH8jE8
ure0oNBpz8++TY8vzu1+OeSbwU1ac9jBxmVteMPbJmznoRZmtPFZq5hSbyHty+L2
Y/MBvpM23L295AW4XLn8OuKC7SDvTK3zqlilzLGEZ+49riwYZknEWZVN/TLHCm6K
rl+uC24+dD0xvYDPH+BbfyIUYGYc+d8kYcOxghQCn6KqUgbhfVdyOuKhjnYG2J2F
c+oLmfuOVotHdSyg+nUuLExjBQuVglaHdWkQOkbKRKJb7fiC733bDjiXz45a60ZW
Wn0RPIw3pyVK9bCJkGH2rDokxqVp06uHpaADBsM2CVvfLYSCnqdCm5OjFZiM9M3q
eHLkNbbogpGR+hplzEZnsnsI60ZMrhDnzkgdeAXL8n0RlAo1q36syxSHvB8aUi6e
mo426oauvVKilxGVq+XaG837zjDYc6ToK3Sb17B2CcdFbB5FoYmxMXSc1FqBklAG
ed5Xzs8AKnlav2R1/O1VV8T1SNOYSrQEk9aw57KVCcOGyPP/oZFJnjjM+K3AvkDH
xPT5nAwPMUURL1Ynm/dZtOxQ7/nHyKrZsrlr4QCnNMTfozKfIlyOgyL5GPeGVqrC
INoiHsi+V2R+C3ld9e7S7v/LuUK/oZ7/MWZgV3Prk7CA+Pwn872AYzZp2oN6euvC
PkIOsTWY7hns7vUKdf2rOaqOK5I2VVeCTi+7MXusVbI3uO0adU3ONL9RJCmIrBRf
Ejd2q6/MP8DsEriA2MbWzEodLvL2RvAb+SkmrwvL5E6SLZOAa6/iJLudp2O/opWZ
meIszeC506AAKPqD1O3emkOltKdkU5+0A9PXcA+RL1heavVf+7QM2DM0lBYPwewe
sopn7hdUVRXREZJBgwohxM5jQsDLrjY8O+1VQX5qQ33brbXJG0KDGVIHJMkRG7O2
aY+EIz12vdal7ufOYX0Ivt7ELhwfrzWTIwcmI69lsq2UbIEnbl81giSPTR9UCF0L
/UjOF0Z6Q87l14MThTntqwWoXa17ioCBLa3ZifWuwloXyTli2xsQIckwcrwVLzn1
EYBFnWlXxVCFLm4/pNpBcE62lq5QIwQX9ofsnASJyTHuXhAceSkvn+WK2IMTdqFy
Kll49ZDVnNiTFYZ49QhBo701DyK3HbU7FCSPI2LqeVr2IjE/FkrHqUjXxqgV78x5
/IcuGg1fsjWh3uPkiil0gImwVPItZXQ/QLMWUuVHJ0ulRHY05Lf1wmkKJq3AIMfz
Z00jvf132Zyw3ms1qrWb8SYJfE/tPzkYaMPQWqk/7iELnkJ5M6DApDbyJxSc/2xF
yXhCGYaFethQ2+1SfqUQ1yy/23Cex7ZzkneGZgAWwQOLQ37coa78WRanP61WvmxA
IQd/mOx+iSg2U5E8/lHg9XwMJHICCvwaXdQla2LT3UtWb9E08kOYiTa34Z2NTSv6
WODjkm6p0aR5r1CKQWRGy8v4mWt8hzxy0RyShcOItqEIPGPJWTue6dxb+2Z/ftxg
DhZTED+f91ju3EIKC5QXOmKj8T2EmHOLki+5Msdo9EAuUjm0w4fccxQnD3QGEvn2
O4yXh++bLefthWYTW5APMWChwJN/MSmTr4mkcCNe/2jvMr752YeZuv65LdRGe8OP
MP5vE1rPSNorKYJvq1a7dksDgAcp1PgvmzVc3u8d7lpgRVVUKDoCQdlSyTo8xjJE
DX4vxUMLZ0c5KcQ48jsIEhbyKWMudVe9/Shd1dDiQdsylXY/ZQYLi80Et41Mz5F6
mT8vcAs4z+6mBO4Ul507zf1rWpUBmn6f/ihVULKAtjs1EbcR4CXCW8jusiGoKNKh
S7/rCznDeCi4ObHY7R8BF1xYief8lve1Fqy9uyCw0gQhUwkjI2RR96S2ddkoGC1U
lbbfkVmS87DqzbU5SnR2H7LkW6YPvwpLxgElw2l/v9X7Y68eofY1u78r3Wo6e599
IOtdEMzbJvi7kHB5LJKwSnWiN7MYblYlgogj5i+Rq9xekjQVdKxwIwdtWWTOlNCA
fO/0P6QBIurFbP8QIy/IDazJgDWKHNRVra+qbFL6FQYVGHz+q2Qxrf4fkG/hd7ar
6Bmgq/fyPlx0Ku8LJ13MCekK7vLpfjEiRyrWwyet6+B0wN5FVwM0phkNhS5LZk9n
3lltg6TSm9lTRyrdEdUJgRvCEScQDc3BYlxe+FG9g34nY0eEo3AGBVcEfhj6uLN1
kZAk4OEPvSbiiHh9KtQmxpBM96MiMOeBmgzg1tjSsbM4odnbBPEG+LVKIabo836D
tpxEOOm4qWtDkV4DK/mHo/2o/1hZ+jhIM/A6zvwXp4fSFSYDe/hJMQuXOR2kxiwE
46t2AFyXdhwhQYkWtHF4+tfe3z+KV8w6E9sXprrScKfcWcyq5EuRj/e2Y5fNhTGR
xP+1LMtdME4Vxz4Fy9Z8ct9fGTZ03TDtnNB3wpUPjEZfC03S+T4VO5/VfWP1jNay
LmthVHGawSEfQWhPxDL1mQNevegJRCfX4sSKVbD1h2IN365zABW1/fQJepb6O99l
CDYo172VKvchpeRfDTS7PrFz3cIV6xkuUf5+IgM9+4r6qS5cR2w3YdebSPaoIBZx
Ya8phdsr8JTKGacgmxsv1lg92NFwTRqXsQrgGIU9XbMKzJlIF+u/3AGbNSamxwEN
ge53znsxlRpIFTCCrfFvZPdNopwsWdufUamSmzwcfAw4vQYTFCf4aagHAlJY+D/o
TD4SUXZqELFqOqQOUiM4EsXWN9YHk62MM+SuteQd7io7b1KWqh88JE6CLYltpg/7
Uttm2D3LvIs+/SepzgNGpQTw4SuBQaYGWbP8T2gnEN4aMu4p73KdUfCXmMJVY/xV
P/KX9+rReR4YN1krc9KVMvqvz4WcxYYRPkJI+y2M/mo9dZf6FRhJD1TMuRMwmXJ4
r/ie3ZXIvE7IojSHbsyvJ4THfboPVko3aTj0y5hnO2cmIrviNvqakzSfZs2x0vbr
ofTlVqoBBTG/yzaxK6+OPX8ZwDAkgtYMQkKdHS+EyHwkQODcn/zxSXvwaM+pS1ny
LIgeKQA0xkF82P2jBENjJT+4bn/V/GF7nj+KOKte76AB3fXxDhhQiFYyXHX/NW70
c5FWP9qjR4l95eIdT+itpC5JafwuvtQz8FqoTTX3ble7nssjmM2m1TtfgU1pK2eD
DksuXEdQ79uteQ+9xnVvn6DtOPvBbk3oMEbDZB1m/AwARk2DRC42QyyzOEbQdRic
8sCaUEXqFcbbiTpCj2FkIHNAABuawH4uG+jgcs/RIAahDHFKlSXYZofZrho1G8bt
ZIVoN9ty/TyX0R9PvvfC+zTH9Yz/Yw0Bf4vlkDi+Fm4fe2J06G+06BjlATeFHgKp
TOlwkL8zG0nt4KqIbmG9stJJW8QKHzHhBLJVEQoM5luW1+j+ugsS0usLg8K5l6Mt
hVMJi9xEHm9sQ9URuhjSnX4Fk8TmPFah6tzp/hh+Pwm/TU+6VWxeLirMMXDxYmuu
KsvEQDbtn2XjvJJXh3i/vh2dssAXltVkxRpYdiULp9TlqYi63QNILWRKIIIBlnHk
9c2XaSpPhetd6eFmtlctIGYTKFpuypNWd1tWOty1iwM/z0j8rFVTpFl5CCc+0ui5
zMGp0b/P3zQgR0Ur/Z/eO1IE4BRSAjETyWau8O0Vj5OX9VdJc7WRCMF2DTOLMF3z
xMc3mmXi6AIQleeVvtPNaY5zcXKU0T2/1fkc4Cmc3iHlxhppZD1R/BelkVkqhr1w
71GSZZkE4JX7UXJ4gFcqdebuEAj7TcJSbUTWjeQRrQL9py2qcObuwt4tfOXm6n64
4zcMFoaMYm2gMTgqhwA8uiMv6w2ck9lcgjniCs1wbqZej/J/Jv81tLcf8RYS1isW
QJUA2shCBF8UeIYWy7RWz0emZeAv3i2uCGNaTYPvkMmoUvbE6zMkSsWO1wGldUQD
QrL0kxBIHnju3Pv0WncROZTp4bmwx9VBe9mOYYsRiBDMtUAdrZgIb6yxG3kjp4TP
kmi9MXuKOYiD4L4elqFViI6GyNx8aH3YjumIsiLzcbU6HhQfxKa/p5vfkvpDthf+
MVLOeWlLqP+3Sa76LMU3906mcQkihUeHW9v7+byiUkgikPI0RiZrT5lGn4A1ABkj
IF7ra63MYoKTWZU3uC7aFPHj7QoCVdpdAOXPZd3y5HfsnvhDBBokqHICEfSm0z4G
PgbaoS1OG9wxgLUfi2Z8r5LDNqnYh2x9oaeS+mDCdJZ1x89GFBsSSLRo2xZlqopB
Dz6Vwf/mtP7pr5tIGLgKAEJrXKcQ57Pif8ro17fXTXs8GY4bg7hCvpsAaOKl6ORp
W8yB+WdnjayOSB0j19a/15F4FNMgYIQjgi12HrlFnhaZ3knYLhDH1N2g6i8VbmOb
E5em6SThVsGnfTSZrXv1saeiC7/TlzE7ujTFBWgc9DFQmP1zuq4v0rGBwNNDviTE
bX7tnAscBFuaPUAu4uiTXWmY30gmqytspFcNBH49P9f0Rj5L3kr77Py4c7jOUp8N
3tpztYFLwXFl8h7LS1KOaJLMbKU3UF0t3Uz1FYUJ6TdA1Bx+owRmbsg7mgivlD+A
AOtWlKQBx8vAvVtzQQRFrFMlAxdBkpOaRJ2AsNFPu6NOe+lTvM+60ODtl30taZgb
7AVRZWSASRBueS+UFIRhx2aibGfGeOmCjou81JgviQPTGucqNkmSOP6j3Z2tohEG
XFl06dpuiYOulngbxk23TE40n5A50bGKl8ME6SOSxYsPxRbT8CaGZSV64OxBMKAf
Z6gWrKu2+4/eS/mp3rpBz0HjkRmPMp19fZHI17dwQJye+dLAFUT5gQ6rH66dPBsy
Ri/Z8Di8CWYC6lX7+jtaQf4z9Qk9xG9VMcDtHUz8nQR6ZFoU10F+Dv+5pikYyQRN
rM8WFq0GG7Xg0+YSjhFP+dISAAhikiLaV9BGSoFIpoh99EG+vgD7H2caGW+msyW7
U/agjw08aN2v5gYfuUQ/ue5aykmYtjiybMqKZSge8DipKO+o0zESwsn16tvD3+kT
Q56IWHRcDl9v8xeLtRGBD0lHQcGpKd48vMx0qWh/sWX29enaUeemQGr/M6TXj198
bBRd3AfflIkCDKR6+PIC88pjOD9HO0JcwOFF5rXPfL0UBobI1RRLvhkGthIgqgmw
ZX6uI0+/jZ2qH5YmKV6sKzh+09HcTCGNLT+D18DJ1k2hJCbrLIhoK//KrH1GsDSd
Kxn0W/6msRG46uZrkapBkS9b7t01karBo2WX457Rp8PchTvJYYaV9UIPVe084I43
UYKwenRVwX4Z2rHH42MNNEswfAIZ+YRR71ePSMrbG9/0NjL/xkMctinXtOC2Qt9n
Z/yYUhU02zCICbYkBM2KzBVvNNTGRGluMmAGYRqjxErncpuOyt/+mXWp0FvIO/d2
ZOFvOVqQSEUj3fkMc+vuJFvn9g16qBhLRG09GQ/QnN+PJZypd7wkrGIlc1syBo1r
4BAf8Y00lyfKrL2vXJW2EcwX2O32dy/mHzMHBS5MQighjXiM1tk9I5xSHiSJJ4M2
MH2UzbX1FSE2rf7jJyT5Kc7516/R9vAWcdAhspJ4fRyUIyP30uwXqjHvVK1JFeDC
z61SGWjPHsKC3gC9ujSrn/92o+uyhdNvJXcvFbQ0eZgYvHrbWD9/XvZsKQHetzYQ
iVhF0GFgW0cKePvA+7zJf8G6yZ4KhPRhF/IOxwKynFTdKyV7VrzDxdPCB8aWIpHW
GjiXZZR+ZulJviYidYZhZ5S54TTgNuyr1bA+SOTsHzgKafkrR3EX3Iy9EsLuz/f0
zjCZhCkJF/B4tF82G/Jl2EVKznZj3Z1MalO9YAm0EXUu9aVctwft3womRaqkPhh1
wRfbktvZOnvIwEdfcxTLVGLFclokPEFviXlQuWx5uEi5IwEH+5K5bh2KK1oPsIt/
Ke48Y0Vtuwxks3pf0C+0f3ZMf5spRK8yCcO3Atjff4lfFOREk6V5KsNB7tduMACo
/9Vo7VZV5egcbg4Y8moL2svfOktslzPwHKyMaa5JCV/pTGwPE/egSt7NldFUbxds
hUwsE+bwh7sdjDToRMopbgke0IbpHWm+58szvdEHGjEt5mkRVB9XwNXdU7lziHka
kEmQySA5aAURa2k3fVzLLsjYJ59Ir7yjvyoX5rs16E4mUeGiDYBzU1bS7Z/zkxyz
Ya6MrK3PU5wHnDCN6lgU5fAeKl5RePx1bZsrDDdMleDJb878jmtG/GGGIhv/EjcR
x5CKyn32mOWqNYI+4EU91ItmEPgnIKEdQMirDmMP0eE4YaiIcblXm11K5uBJL72V
qe2IHHpiWtTo7A27kcBuj/Prlfb2u7RVmajcqw5xUYP1c67k56zoKRTI/D2/txef
RDUt8P/CADUJiRDZ0k1rijfqjUFRqeioBRBAIJ2WqYifWBCCHbZC5UuzDb0Vil5d
o+n6DvzBb+cbukn+/piVLtXl7RDKUgy7fwsHw7EX81MZ5wYOWcsYj0HmjReG1m7e
LqhaOO+ZtvrZK7e1gU0A9sDB+iHRqZyiN/tqOH5fAfW+nb32FHXXL1IrLXFTqeIw
v2CixGH1wxWnM4p41DCS5BAioPmrnsPHF2/eyEsnlA44uUB8VikGLviRVYdhab+o
uLBcgCGmcz0t6JkuN1ch2lc3vENTsb4pRjxo0C1w826oIrhoe3ORlrNhR7HpnBHn
LX8RP43ENq+4KZBulwRqYhY44QQYqfKOcs+NTpRe7AUCjpJVp5FZPduYKEoHFZTg
VTospk7aESxxbBvfvZVKd2t2N1t8APJ2zy5WzbLffWsY/L8l0ZLqZ+syktWdUa+2
kP1Nu4z0SteWnCts3NfEAdRRuw25pTno2MEif+gA5v+ETBtAJQWNk7acMsm51kmb
TmY8MBaM5N656DQGe5jjey9Xvk/M18/6flN0cLDHln4qcHSUaHXRG98OC7d2Q1b6
DJ3EnU12w8oCuFbQpxnstzrBHQmBCF84qow3oN2g8s+42jZMT72BuqftIzV97qQs
+NIiZHGUEQujTBleu0ruqj7oyOZ4NLTiy4HW8qcZMpehqZE7h7dQI+ZoGaCYBd+m
FJYOWtseKKRiHNWjiCxvQygMYysO8A/3sUUJcctMe65lPuZIZ0bMUfqymOVXvsm7
jyPnywDwftMQ9iCGGfLGCAHWBQa6L18mzm1DBGPtjlKEB2Ipy/jSAH2oeNeTxjKC
abl9iXUfw2S167dsrU/cGVpeksI7btD8zpKJ1rsrl5nx8fEK8hQf3/mELTL+MBqo
RA3vPHKrQm9iJopcLWTuyIg0UBsuKJrGBMhnOspchaZbITwIJdrsGOvKl4u80YeH
Z9oTskijcnAm89/y4fpZRAFkxIiMoFvBZoSa+Evq6IaFfXvaeMwsf75UzMyg+bxl
s8p5hyf/4p5izhR6IwsL0GvL1+EP80P2eCgy5Q6hYRWbz5BTDu9HQJAG+65JqEnE
8xb4JPhkoWOyByoNqguXaPPp4ugWog24GVGuswjcp1KO65kTtqU47q//ziemDQco
rHUjVNHoLSabt04m2ATSRAehWJLD0F6TCDR6HcCsw2Kwfm2JoZN/5JQCJUxULYU7
3bGcZa3mbatgP+oGmrwoWD4sgKrHKXwiepHo/NfoxaFLX9diVfUPFSvFERoOBnZu
c+nx3WsMSwqmqfSPaHEK/cgeh8+w7JSkdO5W1M/OZb4864HRrQIbiuRD4BxIja3M
qlskeXE5TkTIDdu0Dhkw873wjDnp30ba7+HqT7nHUByLIiieq7aGonMINviXermG
AwCSTxoeY+CjsfZfI/8J+Jp4cjgglFy9lA19/HmG1jjnfqlSUSuUN8aUMxF/O8Eq
iJALlB9rlZ4XbTZguNT8l6xEMFsgq0QvdLafWcJmHYJOyJifS5Cn5u4MZoQpFtk8
5IAmsljGkWpax42Tl755QE68+0KrxZSeiyi5XEXc2ssWKY6m/kiq7d+tcOucXylp
uu0cskB87UNysxuq4VT+EKGbhF2FMIp1s1OC8pDXcP3oPQh+2NTc3ZRz35CnP4FY
BaMa32efZ/zx4GZxDg5VkJZESJJSS6CFQcp4J+ush/M9bYuEhaY6tKpxB3tQDjox
2if/ZQ70+b3SMvwz6ADPQKk4HnPFqz8dxa0VnuGmxP8jkVwkhMQsU64FfOcuTxMP
s4eYY329OQzN+OOTZAAubfhZPud0Su57cpMgRp8KNPsTvibzMXBQOUCgI8CuNkWx
drOK0plkRdgYElOvKWPbfTYOH5mKBl6sqcH1wOepliVpmPNX8KBETKxXsYvdzRgd
cJdRE+VCo5ltLYQCU2ET0ffUuFN6DUGGqz47IyJNlLXXAFic4kWSZNNkYX0REGEi
ALgBibwI+OwPdr6OLuJ5H/T6F4XMB7ffKx/swRPw+I/TN3b0UXvNKW6QYhJi5leh
maxe79ffeWrjg9Xulm9vrWQcUykKYGUHnXP6BHu33TJ1+pcQ9E8TXY3SEnkzMIMV
+Nr/i6vKFHiwv/oJ+oMj2keHcRt7bR+/RffmqIKDIvS6c66DqGsqKbnwOBI9v9D4
QYB7KzQfRID02z6VeWVtwNxQULsK5/n0y0sZ/xiamcWy+wPnNwjndEr36K9yt5d+
4qzE8beBmGsTMZLr9RCVyTHB3uta8bJ0bZVb8sBWrxzdH3qRD2qjT32kKVajy+YV
VIXtJhAmkO/qzNLYpEwVdokYxdv7Rj0AECJfVlJN/gxAvTdUIh67Jr7vJlIum5Ji
IWaxhT3wzvq+XCc14LIi+gm3M7BNlxBWMYdS1KwMC97Vk+/V+fX9Rc3vwgHnn7pJ
A3NGGgO2r8KKmtoqHiWlfaWQEeYUabeJjSmM9jgFiAQPpM8+DINS16Fw8G1hWltn
KK74GE52pt6r/4M1TaV34zR0oWkZI20RmL1ZF+1qB6Osb3W68p05pR0q52Jiy9kn
eEZ9K0NfQgld8FVcpxQYXkmDeIxruM1wc0Sy4jXwkGl91+hBxiHySrkrCInUafbT
S0ykLXwmty6GCSWhdFUMrhiwCQd0VVgKo95y1Xnn8ButjNUrLpvlZTcOpTxtl+Pc
wOaKPV83fQEtvKCpPuSgYDQwbaokAyC9+LAWAstaVhVRKNZJ4z+7NBUy8w+1h00v
nLFYq8m6yw8hf0CCc2XUZdxlvrGyf+OLGT0jboZAQ6n/YxJ27epRyTz4S/uw1Rno
D28EaMhrp8htmfAM+h4NkZTSAXisLsmFqa4JmM6CfPYUIloFNIth+HQdrt0cbKm5
cIrUMCuJ7U2P2Boopkns5RZmplHWX1ioBHB6sWU1pSmed6gJ021yon+somWVpMUa
r7nvMsoQ1YxTJXtjd3rp5XQsju4s/+DkMaliqXiAYQrzAfzpgIT6XU2bt1R6JWRk
Vu95xGvYt/7U7C2s4SfZ/8mRLgTrDlDuIJi2oVGJuysVngrjdVxYfg0FUiTfN2JM
q2yWepKU2nDfLypGIaXEnPBqXrBK9zBW8a/Nu8zM4wOLxBOw157OXU4BGPS0KRHD
5E+73W8oQll13IB4Ya4akYn62JAzOwuRZNKc0ep0QctYkQcNd3NvAmfkHac7IPtK
1iLDOQjPro7+TmNyZuyFUwnW2kT/EXUhhJsU0XvcgOkuKKO68fssbM0dHlc1xIiC
Z/WeEJZ1d6rhC7nTlma94mBmULPIqkaA9GwSJsYSnRtoI/CJW5brO/yEt0DEh+Fd
qGpX1JCxQfY94/AqooE0ibcyl5GP+8MiCHNeL2zexfPJ8ugOkMRBuGgFOceAqpKr
OUHssE+fZWIqo2hIJTXdrWFI68ge+RXMqLmSEKVz4AHCBzMOCSE30WllMJqe+EtV
yqchwXhcnbn+YHsf+OGegrCJZwedikbOMS6YSH6akXGXn0wbQ+Rz3g85qI6i0z37
N1JTllE15TfZ3udYTGmLVZcA+xX7su+HIU40hKuMKwEJF4GEWcQWcfClq8h5J65y
bpezoDw2esmoKIhtTNLaApEjC+dBO2LmrSfqgFZCrTkDUqjyoxZC7/45bge15cVV
h8RHhFFLSfGfU7CZNzVmwy0hr0nd8x0MOztitsmNnnz8c1h8nYNvnGv2NyDriuHT
makqZbLNOxhH8g8BkbmmehGhK3dbF62x2PGG3Pq+uas9dSnNMWMheQ7Lvl6970Bg
qsg8T0WB+y8ofulAqpyHMXLE/4TezNCx+AwAdKgtAZYB+G5GeDqX65I1IM++AO1l
mT/U5YJLqoF3XacRMjiou7M8m/RszOYYDW69LPTVmzupif4CNinTQ0mTHuOCVYOH
wJKOvLYdP5iK0r/QPUf9j9vCJp6E6s0acNu3ARRgbmZwgGbAQFQDTL68UvCCKXTf
GWXgscy2PEt4r7S0+i1fkBMnfN8EfoF8kf5Nqx9Mgu1nQZWGW+j992urVl506Me0
5zWZJ1EiQefILK2iUGDLk2BWL/X1WOaHp3kJscdJ1ECYGPqslgFjBmPVtbuXeoA6
QN7by7ingoOlgAiczVapfECYAFVtofRO9kCAVOmmcKfu3S95mJhzbxD2eE25kTEJ
FCKnwM2jqVb78arrS3LIPaeBrqRTKlsGgJj4n9APKmFn1O69sqIWwfuCzxCmPPjM
YrVl8qbrugxqKYKMJFJKIoVY6RH9BVZDF6Z+2Lul1dfL9HT6GL/OQcQjOeoAZG8Q
W1ZAzas5FBUXRlpRGoWlq1aF9vLcoXEuZ9ZYClmFjIxn73szcks2gnQmE7khuTI9
xmmyGDU7QvxL7fbpk//diiz4LSfXWVei6BFJfsH6BQm2p6hdwWDoLBggCH4De2Ee
Gc6CPX/EUnj1coQ9dhanJLKdxIpOrGPP2+CIhZVDwVSKRaX1VDGoch9Ny8pe7MCa
EzwNB0wG5GFlt+y1VNK8jCtzy9vNvoWf2rc6obRTxxMhHrQxsMoZDODjXjzFwqkW
44Gx9dHR0DUD6SvVlXp1IUoE83qoAj5qn6z0aYB5B6KiK7boIU4lLvoPGHsFTbEK
Fxwx+U1meHv7veOyvfloMmTE2mswG1OjFz5CurKaFTYhPmzyaxxSQRYaRq6FQuDp
NDUT3fnBlTCNd9EJAQdum+spEFagEtQPXARZfEVGgwDFX2GhYGmR1yxSGGCGsy0h
Pws6s7fjf44OlROzyf42KqP3nEVZLvBRiyl2SCKfGYnticxinsMXBK2uMCihXjHh
Cwj4TvwKOWGq40U9qMJWSJvK8aWTrfdjk5AcYGSrbmAEke6oBCKd6kxeYZBJ/xeW
7WZ0aKBzZIKQTmxifHTsJatbSDLhWgeA8damqbYETXfqlCs4p1jIfwBtX9RVMNaK
5dkEI68mWFQEwmFnrVkaCqlyG6tRhhcoLJjODOk/koCk9cDlndgn6HEbPOWMI2DK
HljNdbGUu9YyuBbB+lhCFafWMh869NC4Rj9k2kuK2eDAfmsmF3P8F31BczI0d8b8
9mciSYikPUA0bObivkkLmfd8P36qrgTB3Wv+o10c/UExQtmh0X9WNHmNF5lWt1nS
Ivt5IC9G7K9LysxtH8CUtqH0RhRV98gxoNkMluJmXjszkq2RLHABuuuZ8Sfd1xmx
ssa9A4Nz0XNwGis0U+SJ0QSiR12NxL8zcgRoyT1Mlmr7beV56Y0Jl2DrKggDDyj8
63sinBFFVFnbXHa7OF0/HDHo+uLir6c2oYRMgFK5t3k8Bjt3W+pNNWfXWu0JmCtL
Ui5NAh5rpdTCS12YRLTfAucdMCOYFcLxBpp9oZ9VFrhDm9I0JEYOmUW/pEG3RygA
kUHVPs4t/9wOLnPx28Tn3xMr4LSw7SiXCtjq3jzlOWQzuxVi96UCiyd1cgCkDa8q
CU2ml9n/pPqTF9PFNR3JQgbiR13Y8ICs5qnT59YtAlAWTxDLenh5osYHOEYQHaqF
Z+NLh5yH4KfA/HpAfyd7CHqc+v1rLRJh43ko2Y9vi9JciCHqFLkv9sOFhPiZ+u4O
0iTBk4K5d8GIZl5qNR3qh0rnU4IQrYVoJKKubXDslEKE9aTAM8Ty08yiu6GFXv51
davA6dKC760H7zeT3MyF3cU7esu/70XDt75N0Fljuf72G/UM/H50cbt0/r7xA6ZX
3CLelDlVxa2MtYSsz+Vj0FEcapVM8n113I9uQI07HmJNivGMGwI+91K1KYigiQaY
3m+LXbm8BCegF6lRebgLdQ9zLu0oagYFz0ARAB+KObbh0YmJTQExX3QgUGJDK048
zsmwakdu8Vsw66ILOqXaie8QjuvWswL4xuKZALKvniNC/7SPtGX1U9SRvxQmPWg7
arHJqJil9Py9Xq0rgfqVhQ/TnhElcuNivtU/S6/MKf59PYa+IRtDO2wsH72uDIQB
P7ENWI9DlM4kdbStx84e0PwwWFxpwE2A6YBor7KMbBkUbqX5+HxSUhyspEleJMPn
4YkoHMgFGa2vil3kEtdebjT9/RojlAZqfoHRisFxRVO0K/zOc8f+SfOuYSZMUHCL
CGFcSc/VRlv5v8ZQE+zphDXHJZIEXBZmsd65NqrmYTCWxt/gMbNVWvME1z7MaIf4
HdbL5yNgE5myhYz6NGwLeWr9Rwrs+z4DUsWLB1zGhjVWEn+0BVxGpKv03EWf37zR
6AHtIKO1F5gaG8Ts9cBoP6q2IfElcCQNOwlXHNsl5oWaUSj4cegzJAlUc4TBu600
/RzuulFcUvexNk2/xANVXEBUXMhcOmrm6PZyHaHS/LwJ/h0wAMpGzzwmWXbOjEK6
8678zP3gGQhkVfsH4AAUkukyyM6rYAAdqn122ZaTuM9veHN0AMeGGmfn5bmiqBuK
TvEJoDumy4fHUCQkOGPkPIYsaj9m9ie+5YF97oruqLEME6DfX6AQN1RpfGSlbZ/v
t/Xlt3jkfX6SaMbAiXFs1LLX2eYFzvqbAMsI60PACbzNo+/m2FZKsVNL9G1WPMTp
2rxCT1dXBkh0rgmoqxfLkYm2gnmeVZEV4R+tu0I0quXjlAm7Me7kIMNagKMiasV0
/U1BzhZiWdII8BtTpIk4odyKMBphUTK4ZjE43kyBPOQ51+Xx1NGO1FpQDM0IMej6
729kIZxZXubQ2JLcKq3VuIf/GoBf/QlYSnYkJs5KNugSTTjwXCyxMHndVg1Qx0yi
tszVcE2/tmk3P8wzbrm0IJdMrszsAe05/UMETXnVkBjxOu77UYCTg7yCSu0/D7V/
U76oj5ZpKjfljjzBQyL4E1ZJ0EAc/dDOersceLH7OPi4c4FSaxMORyqmkjJOGLfF
4x8CAxZO+0CtAX8yHp6dD83S3tbgMDjRACYWKZ5DZXebDfJ4ZJcpxGJPCA7SDfHv
nl4odt8ItTDbUHenTOvP01UPcyAEZkyhx/D7qqQnSwFeGwp2CkiKqv4oOzopwY9j
SMvuy2JjcJr1faTTCEQo0TfFZjzWuHcf6Ah4pPO2ONyfTBrBZ7fGbRD471aEbGQj
PjAWRoKfAXBlcefrS0FPb2a55yw9tN6kSiF4tn5hBf5AtPFgPGeYPRyLUjO68vfa
/pKFpUs+lIh3Su79/hOZmiY91+2DeoQm4byqGI/HMTM39hz6rm7a0fkX5lTky1Uj
D07zwP+//Hk5wWGC9mB1rObVHnb8gnbka5DSv971IPc6jtuZItKORVIGi1+6zgdn
D58VlrOCeTK/9FRcI2gaOsaBfeEWYjxclBu2guUgaoGzK6whHgEzEj7oB2LAXY06
AG/cgUJ4Coj99D9toxfNkE+hRGht19KFtFgAbkU1TrCuGBYxlJf7RuFu4bjdSnin
hqhVWzNl8dneuaQdVz3HcEsBxmy1bkEyI90dr6VgaCQBElzbziOrXkMw4O1dBoCu
A9hu4V24ExzI/Bq0bgkb+ofC71NzebRZJwMyEB7wenBrBfEiWfGpDOV7NytVpTnp
rO7WN9J+RXNoOuITaULsSeGCKWk78stf+/N3VeHaNLmYK19n45soZq33tp449g06
nWflmyt43fqEZiX+SZ/qGnYlqoRTxeskqc3lWZdMQrsp5Rid5FshXbh5zmh5zkC6
qrRjWmh9KPrmzL99vzAEdc79xki0RJIY2+RX7n31x+iEjgHYmndDReaVYPgoP8Y9
yWnLWxlsthKX4WTjZr/F725NC6HHySI1rQSUe0lyUkrUgloV2r3ovjOpC9joyVsw
CTOaxve1PSJIJ0LQ4qGSc3jaWa6JE7Y2wcGOPO0HONm/FZEUvwu5NTCCfr4wugKE
SJbU/XrIyKVctK1sH18EmjEGRi4WSatPTPpOF89DFiBKCh3cPe5jmQjw90Wkww4U
jlJrtfRmhevnmZc/YXwxFb2h+avDl1HeZ7+PkCWVPut/JAuiHnH+J+JC/L6gi6U1
Zxftgk0WKb1hudw1Vrl2UwBNfSOGPQd60lgQ56j9bPvLKSySVEFy5q95//0bZLwp
fMyMqJJ/s1nL4fEyAcOGjJ0jA0MJ9wppUZbJKt/wKeo8glItxPlgw7g0CbzkvQIy
t26nINDgycDuddcQgdeG1eIg/Apv5E8p0auh9IuTc+GGDGXLElWhj2pZURIBYLNF
tgVYo5ff96tklRBkMOt/W3GdUpEpTkpH+c7Y2SFtWTJZfQdLm2CK8bguUidbbQqT
8v70DkNVSZpZtiAE1bE9H7gIBeScTp8LaAdTUPulrqG02Drrg58PIyKjAX9r64x0
xoM4z3BDngYksM9Tg3x4jcV7l+O+BrcYH4EkKD+XSd6+UZD2qB0yQLIwK/rJCc1F
fvZLVE8qb5uYvnZ/W5htDPq0kCmifgaXuf+q/VkHyxFpUH3nKnwrm9fMXISSr+4O
NVbqKq69BaI6NyPQli80CrM/W6r72jjXhsRyy9oMNHFuITHspVQNML09dtxU8R7e
iK385SAjoPfzMDqVnOhn1p91HMft9BGNkHAspjEnQwNemas1ShrRCF8yWKBzvnz9
BirC8oBWkYykSQrBAp5Hc1wqHzCoupa+1se6wyt4ClSM4+rLoATErdAV3JVRd1XR
6bbEpr2BpZFVegdwXaFIvDEfAoFfTjd/6fi0nIWGzl0ONw8RHtKQzpkf7LFRaUyy
iQ0IYq5tx7bOnSJLoLKB6vL6W/CRawt3OiGPeTQ5HIQvVJqojjM+HrD81RHve7Wv
eij4a1xhtokpPETUGoyvQ9oHlwKYVnZ4Ia4gScUoMc2s/j/9a1qDJdJJQVozfPUT
gXhjn73wS9JBQKnCy/PgUtw+ZB2e+FUkQjyrK3Lbj7QrWRL8knVxmjgXcytlfIgg
wVAxsnum8ePRWiSsK+f9M7LkxuNaXCvzWfQYjqR5rE99CS/Ex3dA6dA7xyO+72+e
Z3Xa39EQxRAHwFrCZbffsKppgWBqwyGsCuyE2dbENiRuTZiDwdGFhEvcHup6DDxz
ogp0FBfqQtKqqiiiAMPOvp1s5URDj3J07t5fC6p7jt/53oLsx+R4RDWxRq1OuUby
wBu98UNi73OTygsfDkOPsI57m65swEyy1K9slkv+RiBxmUa+wsvcv4J1ic/Z55XI
zBxNmLPgm8o4O3ODFJ5XwKmrRPa3vepI524lZQIRITXska/VlIHnmZN3+DHk3BV8
z9uBbDMWw13RJiy8e+mvjkeV81ZkNxHVj5QgYZov+yDi0qoU77aoC5sTFnVq/5Pa
6IjJuZ+I4RU97KY2pwD84BztPtr3Dz8HzNwwho8s0I5uwR814RZ1DrkSypfxFsaK
RH5HvV8Ay+SAip0AZ6LY0Vspm/Zv8oh4DpRWn+o3DLWijnWllHxt470kC660avvR
BsQWQBYuhPxUsjWHhGrvDbtPERumInLi4VnmcgcOumEL+/BOQ3+qqi07PYBIaLqr
m2DKva/t2CuSLo4n3b6vCpyyYyn7KzmVGanV1gD0DgiYOrFBnYhCV0+603inal+w
s2/zkkLD5adfotNMXMy8rEhzD9v/K9O1vA1Xlb0FmjrLvI2/vyMMcjOKNv24ybxj
GAn+JUNiQmW3ddN+UnzRckC9Jef/1GJrb9G6MEmU+4rgauYkLihhF0vBKB1HaNN7
7i5XwxXRE/dzLahLvC+VOc1L08MmJHbxKl2T37ydqWHK9PylSS5OW2t2L9wzGMXP
z9qSY6RogJ4VpjxQWluSTZaG7H+SJELipc8dsV/DLTGvr/hjHXpeypYO7yDYH5bd
1F0Vw1BT/90uvu0jGGZOCb59S8/4E0IpSpIGuVkKwBfJGohPMaE8REwjPodRPrUH
AKK28H/KwedeAgUFgrhUs3w060R1DuLcSRGZ8PgEwsktn8i7iMF5Nm3WkhH5WpcZ
Cyqy8QvJPAfsMROha27lGgsA3HyVogeSSH+KD35/8C8ODoJEQsU8SY+PZWpzfyE1
MupkwNWmfD/vpGkAmQfIOFtACFhmhqxoqPsRaU35cqfCnFrBTc29aXr/qGbZqTsE
Y0SzIsz2vWBDZhYl/rjKnSYyVaAUmPXYznfwdpYsBC8O//FTT65z7HcOnFgbraYs
NnjND/Zt8B/gSm+it0sx4GmXeRCaaji3wk5k4OBtG/4+7uK0sxPJnrgYBNRjgujC
EfWvECX/9BvsVQ33jkP4XUMSZ/X2y6nr6wbnL13Ru6o5bYvVf08TZEk1rrymyxHK
ZToKVBiBHtT8SG35My2KacNgjacJSdb24SG2HYp4XtqhzQzcGasMFdKJnoZhdAaL
XYOwpNc5gJcGuERuz3A6WXsuGAhIiw4muMf882X2qbHNH5ZwkBEe2hNSNq+pRc0d
ORkgdqJXOsVTGxYLU7cKSGCIG3MLjWQ5e3lOoml6x/jqOg+UMDBwTw3kcyLgZjvV
oU1zBk2i/8oAEkdkrj75tR0ZoLqFtmMHnVyaIjOs/rFoNTGDNXqkCsPCf544bQr4
NpyuE16aaykn0jPE2BaRMKHBzvBygoNpz098h/a30rOfHOP6azqDA8+UA7YsIUL/
4dH7aMzady/DdBpBaYb3LG17SvLWS0tS2g21EZk+r62JXdXzb8Ggn63b6zJS0e0F
OOvkJhpNSAmyKj37o0FK7rFwhcsoihc8J9URMG6uV20wB5Xl5c1Qe57dOUWp/9q8
gmSiktPzUr/OadIfO+dlR06ig3K3/eWOAgWhyBTbuBSHSnZRVB3cnbQBIOpKVb9d
ko1o7fTXOtDVKp7RVFozGZDYxAQQsP7guWDBwn2vpIcpJ3RLc2l21FQZeUTakBf4
+hpTzvDtULRUWi4zsBDKukSdkV6QZy+FZk9AK3ICr6Iv36L/MBQNsUfE5LmpbW9S
M9hkZaiKq4QYhj8/d2tPuBkPm4qe1V9hC7bYagH8PAv5aoneNo6s2J9RvYXVJhCd
8wJHkYjNV0FbDCVFMgokJO9AyZR5Eu81QWPHNKLsdAjPMCnOpe2hGiUDKo55WAss
v7hzn6cekaudxjpnKTG3vdZvpGUXCmMliDssvcbTfOvJm/Dug0Iz8KEL+yE/nEMI
C0ZqRNO1XqYIKct4QGe+jIOmt0ojsE50CNBSGmVJIVyLUNkb4RqHE4GB5NjltJyX
lIWmglq3xwyQy5Zsiu4Lctdls83IPRew0SapsPls95sbHOToaHH7kLyX8x0JXS4t
nviQoJETSyknB7iLhwd21Hf1jmn7w/hRL2L9D+bWNFROK0DtvsF1nRlMTIjWTEBf
smLqwaP6zDVOlMdBWXYzO9PqzAwil7JoLTKcoMLsoKE65nyj6ISEChqtCsZ9XIKd
Q+rdZVKYnop5KKxQBEVXk48QaIJgNJHasVS/uf9rAOIgsilPqa/PqW+gsA+oRg+g
BSU3SBmktSIFLkFPk+9vxCaxVmqj3MEzSnsnrfdFP/7Aa/5wOsGUPeq1IpCd0Eup
lOTSga/YjghHld4S7dx3MFmeErfMjAp7X1Bhf8Q8POmikn/c1KqepsEx+mIyKcev
lWIgXBbbSEIxdmqRb24rbH8O08gRsJNyaMCc9zPZFk1rahuO4oYk1IG+RAtIlgnf
E5Iye3KDNFdSzzL48C+YK9290dLLnGANZZA8w6SI/b/gqYMJRgKxjtvho3CkQqta
7Y1fXHi0vRHZAylUSROT7ul4WffZCYXwiHG/mGuX/VAFjxI6zFrOzX7F41JcJn45
LvpS1dTLanJSL1CBwJsJImTkzYIf3+AWBlRg3EY61raNbYJryNtZFb9JI5JfqIgA
Q1WVdzbAGnxvVcTkur2fEgW+OsD0kaNjWUDPlHDxgaxLhQ/HeRai25CR3aTtMN4v
zDI9270DIMw0nejEAhrgOgTKSBibjIhCXHnWzQwfPoEY/ITnTd2AR8wn4EHrI75T
QE8EiLPjbAfpJHmOcChYYz3oADVs7AChNV8T9WWdc57lHEBhPf7SFqa0vQxKgeP9
s+9XcJAyz4j28nuwocVXq2VSmkyDLpEmhcqLGv8ara/XjVf4/IGLQ7W3oQ12y5er
K1tPeb2tPF4JWxv4x27fNUGokkJGqZ5X9Q3lACx8gtiCPJY1CQmEPy9qakcdzz1M
v8DPx/BCspueEK890Bjk8SUVNTLlkWDBvyJureXc0i5P7QeE7Fx84GhdTr2zNvL7
7S+4PGhuJpr0ay5r053bkucsp3xhMe3aVFT+9wdA2tOUPDgWTuvbnX7zQzYi8LTr
5FzZ6JODwaJLVhmr+Cp8is8Mv8nAEdP0MlQSkFimT3/vFg7ASdLAoHbFZGqv5/c2
Mpcqtxs5C1vzuw+XLP0sucZuy9UlKAr/+C75xbrUrdsI8hRLekqOD4K8/Cas6ZPT
7A868NE/Cs+LRXt5gMRQ2pZiPQMNlyys6dsmjAmyZ8ZPk/q40Br7aNnWdvI1BIyy
RtvRnMd9MxYaWP2xm7HLzYm4oWITaqTvvvKbCZikUUyH+xj+yEw+J+XtEnTSyTMz
rr4Zux0kmWO6KkHTfxytfFx9ssMJHoiOUFDj87VrXA6fbjAi9pxUuKgnbi/TCZxR
QCgW7wHcu46tXlPrgodGKFc+TmSzSOjuSOFVPO7ebK/tDtyaRJK8ZI9R+iUEs78v
E5YY2GzDq6j1zzbrq/K6/A==
`pragma protect end_protected
