`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
T/mD+NaY8n6p68cK1fWYYwYUCVqnc36h9kgOZUCUUTabDRw/0bSNUIaGdlhUeTkP
UAGBlYbEAOzVcWPZ7AxTx/hXUhkUcU+ImCyXzbgpL5zq8FCJGDmcXvDRoKQOfJcc
muVE+LsO59W6M7OGBddlxv4DS/D0oopw5qJ/eavIlIc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15872)
e8KIAfKpwbCsLgsGw0U++un06HkB7AU9TyvN/f7HSpcy0CCNY+YfF0WeTzCd03QR
E+SaMAuSw99TS+evA9qiMbZTld3G957WdV4Y2/ARHAbjrPQ4OiNqeTef5dnUFPiK
ZhFd4uiszPNDWNgN7GS4LDEfkpUOXQHkOxh+Wmy5osAO9DNT0eCrPNmcC/U2QEbx
njfrnUSbUeJKy2D8JZiWtX4KPpukbb4hJxLElKJox6RzO/g1/A38qeiXyN5voKC1
vS/FkWQcTB7lHsl+/TnAUYGcCyN4N974gNCRss68wi060bG1dXyzR2yNVGZsNsc8
tZS6SR16ZPzMIqLEOmKdNerSPJoiIzD1U/jkqhB2HPSZCuJBElTBPYj8Ycwi5p3g
ZXDYNAF+YA1PUWsNxOXEaIWpWv8zz34NUvd7GV9W7fjc+7WKUFuhK8eIjiMczi4x
xqjiW5vf6lWbD9VvRnCxYmQRCR/AZtvK4k0pM8BVWefYTxApLkFrovbdXyxN9iC0
rXLHt0NQPa3OheaffpGBiU/Kd7QACYeBq+XDgMKksGd4li6QFEBP8d7Sj03UCNwn
drVe7GJnH4Hvf2/kfXfDH3Tzzu2Z2dkUjxP2RfmZe996hr6q+kFvytON47y1lQ/l
qtiYjPDjUvoeGGFgKeUY7zIisMBnpyg0i0QYgyqM/mts+tgFwC7C1JKMJ1xymAoo
BTSezq13J8u39sWnMEB8Ps6Sp1kqH5oURrkQN0Mld8KnPDRdYnB5xEzVRfSmeWKx
wbt/wTby9H7dOZpLe6SiUnOh6yhT08URV9z/7qN+mEi3buFUtli2LaGDerWJXw8G
1jjjfGTqUmAYE8lkwTaDUZ4Jm9D6PPSBEe6up8paH251ArmdJnjrHUk6Q7iTcwEj
uW/inAodiDCtOGO++8IAgcXQEeVw/Aphrwe5orMiXXIX7WgEHhv1XHFpijgKR/F/
nDOOy5yDwRKvnpJkAgK9TWurTroRohZGeW8U63xs2XlADKhIB487S4ac1vfHm1GQ
Iw3/JJqjEEMuT4y50/deKmBcxrDNICdUno5rdQSlP4Y6dCm9h/2e/gN3l9IMeK7V
bwmJaVocnaSoWODuAEmpCmRv8tV54DJ1rAXaWrzurnOU2+1eInOyGM3lW4gi0GPv
LEGy5dI4AohluNooKUj7PoJW10/2cj14DwCSlW8jPWhzOlZ27CLkTfxMg0/8vPKV
l8HCJQXBfBEYb3K3tP/ycprwrflrbGhCKncfQrgKJPAKQi2S5Ku79HM7s9l1ALUM
BwRRjf4UgiWCSRamdXVJckwIkzc5MmK3iUe2EY3PHw7VutzsYwKzIbTnVBAhlqya
mgP+wIEHCrvzv+ApA9jm+MQCibGDz0tqmlgktGMJKa4PiTyJYkT3w9znV+3QP/i5
Xv9/oy23rhthpuFLsLY3ZJGhsnZtFJDxub6lTWnf54s8ucXNjy+1mYgPu1Djovmv
ey0yBehejjL6oV9vAP/b3VV5tp0pm0nQ2S95BiZpE4f6zcuya76fO4GHEB/R0aZc
toEBJSXyDylryNC8HKn7J1UMEoDjdxfCn14NvjQZpFQJ66PkPEhbWdbN/x/9Ulnp
0lelWEONT1MKrG4q3MNqLUQptx+yIyrGhJkuVk7nE0moA060Yx9CzQ8mDHzvl34X
hzmTok4LP5vwdpYhzDMWYEEVbnZ0CiwbObcIWR7UQYaGk4Dx3+tVIo8tzhIp37MQ
cQOUQ0L6RnG5aevaPQqpEmYGqHKudfHsTNZE3P3quHs4mC9U7rGv0AjRHvE05r3W
nZWx1y3IxIGbWl18zSGTwuck+qG2NyVxl7x1A+Hu0vvhqMQJsAjuNtiuGIRvyNU5
eKj23dcC4kMZWFute7SHqw00xRS3/lvo8iBcUJrcb2MHnbFL+p1MJdEdyM4mJFnR
FyL1nmbhkyl6+UKzEVoDsOSxsVam0JCZN/eR10/pDvTP3BsixntWyuwvYJ1CctQn
mFAO5B63Itkhchu0yWGw5poYsNvNsKdTbhl/bDh2tAnom6SVQqzCZ/Lyb9g1cWz+
Howd+vkRQiN54I5KD37bOHpW+hfSyal9eX3r6vkd25TVo0A9Wylan7yOGU/ipaVA
SDS1xIUdq7s4YdOaGOgVVeweAEsUzjw7Lb9bD0nCoOH5NmEa992lVm5u8MlHJlvi
ACzVtgGrmtzhWB7XbmQ1fzlCqyvGHCRyfbQdVB2AoyhnWNTei/Q9qaAoSsr6u6+4
/NEtwlGWFlpAQSY/GAeknGnv9GVWO0Zk+d/0mDINIWMoXlsyo1QHx1vY0u6EXxKy
NvYs6CkC5K10d2JmDX8ASZV5Yrxr/P3ef8qevFOBZME9WA8j+NGJoLbTvFlt3fag
AHqPnRgTBcctuWztePQtM/aTxSfsWbI/5WWRjTxiqxUKGzsRkLv9X07stAp+9FoH
WRKWlMJ4eGwv+QvZioPileRHWE2iccvUbbDKS1+DCI7ap8+oD0fQHQ64sFQpnomb
4rRDDXsrwIy5AXqY/E3npumUp5y3VJtREFXVBB2HMX19c3D5QNihb7/QzVAUEu4M
s4svH1uFF1wR6TMZUBCjlmeZDNEzAT5UwDfwdQxwguvZwPAHSid8vDBJr0nnorWa
bL8YpXMcyE4lTkvNEMgyxbjaUVM0oi1e7JU6nAGU1goodP5Tq4LZn3yVE+M7aLVC
zpEFrs66aCQjkzwahkBZTCG/wmavUFQ7uI9ONJXSydNb5aUtm/0Nuhb+vNM6k9D0
uL6nmoiVvKXxKRiyzK7PmMe8f24lM3EXlqJKVNcGACAcwXZXNhe6QWyAv7cGDlqz
dythxnlLbR72po5JaFjfArLU7vIi7Yu/bnVlJbofQ9uDHxanU66tjPvkDTcr5w7L
SDULAakdiOZ+iDcOmoa/9vWpKZDMtovwri4GGoKBdnaawGdxZzzizBqh5hgeXKnF
s6nJ7rl+CjmLtqi3XV/+AHstg66QWsBoMYyejcSkkXeZCrHr+vxjHBpOC84oL2uW
jVd3NfCoBzj2W7Ue/GNGOZtYIG+m5CqZJvJLXikj1sLIwNhxorX6RnQW7iwuXzLe
pFTlhgH31+r8iFge+xe1iXmAyeOmyIxJrpfznZDQL3XNctQX/8Ln98p9/FlCd9Vf
PHtxuDk/4kt/TvAW2eAfhfcieIZ+sjNz9ZP4QbkH9JvZOOF1Nh8fw0SdA2XvdI/S
fu1q5VANLKqh81CViRyKa2J7ky/GIA9OfoLhvuxH1rJDoJiq70ZKAm2sTtk6GF6A
DYs1qoC+f0tHRVRbCkhyqS2g9Yyk4q6OJX8/knylN7ubhroBlOwQqpS7SwV/b2ua
spRGYprUuk/Oh///7HGtOk5KOjLK2abtE8lYu3/d3w61syFw05nbwBa7yi0XwUiS
zOJ0wf6tiar7iuYud1P3XRQmyNyJpsd9o6WswUEb2TQwI7ogXnbGUjkfYpPuX1xp
Njzy1mGEXHa1S6hjvjdv10rMzit8lSXGBF+9GwXxEYBI4+H2HEzoxQovlUqD1AaT
6af7aPcbMZovTbwI+hYva0XiCxl/lwb9GXptW0WJ2iXeAvuRx4+DWNxjljlRJIzl
iitzmZ80A3cFVCA0ALAS+ZUfiegOCdq2iAMA04d0T1PUzop7uWebYwA44JBhHZMl
/Uj091yg5XJsSvWtGE6t35uh2XMHoQfKKa2lwxxa6zfL3nYD0XbWecqkXKtVS8F/
0CCej8U734aSG12QBolKSpqTPv665/nzRXyW6m3iVWtFEabhkltt+LH+xNFpXjF3
N5AqEpqGQKYUVI3gh++uqYNvL7LkO854qoMux7xFRZPvN395n68i7dq8RBJhOb2L
Ww/AsyjicsLNRjMyupAz0SD3OXPLpLqry5cHj5//EMjCeZwLTC4Xc4Y6pLbiRe8T
EOiGi48ZZQb7raLhTowpI4clNQXL2EbosvWxZR8MxoOiW85nofzlfkk29laYwKpz
o1NxwAukzjlYsK2u/ffT9R3rLgcj2dnjWI7F2Xw6h1mkIaUAhmtbMTLFl77Q1yHJ
7ZRM2Ig+FvNtDkQiWCV7BjzvspDqbcopGU3T6mYhsW1SKIA8TRJHZTfL41Hnr24a
8oPwAUGQuTSkQz/fEyNhw6pYUCWuoUSPUqx0vaMlTs9ZSdmlN/d7TFbKn8Znl5/i
DgOW0h95z3DGwQ1lTvf92dl+LLlhLiNoq4H/JEvnty7rQyDHki2ezPsEQLsI8ptE
aI0PUCFoRoh8c0eV4lYQ1j+WgWARp7dqaqQcglwZQ24GK2zeMpb9E8f7GdneRW4M
CTM3LFhokvnrG8Rt3wdNq2DONBymnVhJ7QKO7zXREPFtpRvcFWibNiGuLAmGoYDU
sf2tFxYr6Ufyej/XXtumjnjgidSa440cibIHgzfo0nMesS7IrUTma0y0kLgR8yga
OSHUB0IorgJDlXiAyjkxuELWTYWVQiDcXIfAyi7zm7jXTTmWc/aAgaXMtA9pYwes
cfTSS0NIpLZAZj5COxtD3HcfMFG5dwf9GVgGCzntLmaEfGIo4Nt+koQQZnhXuTQk
VZDW9gA+VdbJ44XJASEbDYFdLDEcy8HtEdN69jtT2RQec7UX8GRghfbgUQMTqCNR
f54PKCFSQxYo9PlJB1TWoI76bC5Pt/7qOfskWG+pxzpSWZ3bimxIxf+o9efnDgky
2VPdiqHwlZbFHyMHv6Yp4RX7lQ3Ze9VUuETSqBKe0hssfS1q14fakwpXoClSoSwf
mk622OkkA6QyP5vcwpCC5M5G6rQCurpGut/cQ4e3ajDPUpIsDMKPkeDYW0Gwrx7c
aag5kHRumXXEqRrm2MKkqWrnk5PeRODOUYk2hHG7BdY6eRJ5hgXBI5c0h0k4YXCd
tTqVDZRUqnexUURL2aguVRgApSm2E8XcTBy0r4uYDRtp1kjZjp9DPUN1E81bMZbv
JtkC34FFhARwdc7v0S+7J9JVXkDfGnIYaiK/9Ytx4aJoORNSmEIO7FNa403SwSIq
lewubz92baYSfxctY1+zneBeNmxRUBUHuJ+idYozcAEsDJjE5i0eA7RGTnNetEVc
UY7fijNCyfoOqk2ZMB94xf3sDKS5hCcVbwtPg6CM9FEfn1jy0LszJaU8HpwwW/RM
E26P6fbjc8p6dc7OnIFlcTkd4sTFBkp6PW5UhoSN3Dp7ckW1C1zO4OvWO7rQeVU7
U1vt3vTQsSjBiQv9TBG+vvDazKe0WvRyp8oV7F4EEWH747mYJty0U9kh7PvnN8sJ
sHuw4BnaZNeTCtjXCFEDLyG/SAQh1zvSLXsm1oJm7yaASm0lfmODb4aSTVC6VcPJ
5PkvR/v2/aoVoEy/c0Ty2K01DuA9S8f5rw9HaEMjAaAc1+3iNOmxm3+LuA10FHeO
gEGXAP6LFlBG2kSqEeRz2hPvritromL3PJgjk3Y9yJVvI6tC9atcZf+Ka2mY0FyN
Yovszq4JjoKe4LMO9r7XIdy14wIgCwraTLSoiVhvvLHX4JeLqThEHDd//5bkW5KO
e45xwa1v+obaGM2InMblz8/cEK8uFVO/94lpLGFQg6LjdgJBb9wexbXPiYUjA2rV
1kXiVdS0LdvMqmqE6XDLx5V7v8+y4ocg7ezetHXpm94L8vFRjJ0UKxSsjTOh3uy7
VoCOv5ozhM6fyNSjgEDH7dn6KJ5p24bLxPfOXWInrHmOjJ7LC7GlWE6NUCaav45p
8Wi2d0SYiSWn4cRDFBuV6yGVuZuakuK2T1c0/r90xwOtdW9Wybbj6Fu2eOOeMBPS
wLOOPxzvlH3NwLP0wPvE4jSR/UMufl6VH2tk4M6xMGaO3YiM1BJFaxVCcQimzX8C
0B3GqqZA1bfPUzFWOYvo/fYwi8Lk9YEMvDsMxQrRHVuASlaTeIXOAnUw3FLOGID8
PJvLKNMkCAwSlNIXUoRlmJ7KGLNNUfISlRJEcMFcm6/qiByI+3RDYkgbu1q/QYbh
ocFVChCAhWe4wFNwWXKPFd7u8SxHlUgj7hi+SDfWqAzZno7rQN8cbyr2HdwxSeWt
cT/xpvMRUNqV0Gg0J4w4I9xa/GVaxOzmvT2AV3iyzQiVg99q9cv++uO504wkl8rz
OVUIIxXWvMiM9lgj0f/4LUKiC55RilYWexup0EPzfq8q95HJflp/obT3rImTDAkU
UmG7zx7xz8K4V59ggsGeT3GSuOxRBHbRPosTxnEDWq28oz+iWjPBk+Yjx6fTycWh
0/xREhTPStuI6ry0cx8EUeHZZ7oAc2UYJBbrV8Pnde7vAxaDF1PE7sUcioUws+iJ
sVMtSRo54GAfTOBYFhhxE3GvFLcXqE1/4JNDKRPb/EgsVG6wEUhDpfmjIzA0LsCE
mUcjzFNm8/3/AN1jEgBjSt7+SFjyH+ajhckwXMtupAHW5Boym4lDQydbmctl4yff
Yctrji5kpXyXwAaXi3af/nyyAE0uopD8yLHj97g3FoxetYhiYq+CcNWJaWKiXw4c
6HtDI0/ll/gZTATEYUGDmY5HhzGebSvWwChsr3KvXqwsmYf8BIeEOw7ChZRVQMrJ
4AAioFLIfnq+wU6H4jQeIu+0KFBoEK1rzIe6De7FGtBxrrHAm5hiQP1rSH9omKAD
b5k4ilOM5ZQ36kP8luVdp4VCTPr3iwCeJMV3tnMt+SIXUTlwvZCWANYBJQGAXQXC
4O1JvdX4f6p25bYLVTq0xvov9H8b5KQt1GV+0hZFkY88J9AF1ALWTerjp0on5yqD
00K97UhTMwFXnpA+Mt+XGMjUPB+NnGYpPEEOWG38H/YFQV2/fJZJhbNM3wxmJ8ZG
8InQZP6UYPhebkvGU99cK4Qgy0M01mLjgf7hpPBJKUIAKf908R5068wgVDKPzBgu
kQ/DytUdruic4PGyf6i/WfWVWUIPYx35416/xPgeAzsuvmeFNsLW1J84rcCkgrn3
SSGelfpfMoB/elCK9iULNieNba3JIjmyRuM6e4OxMaHsON1rG/dJfR9De+HyLdsi
xHv3M53LfkKnF3SLAoDXuX/SG9WHYzYJLCx9LpMwafESzKRLsJC7LU/jLoRqLYDB
ZfPgNIpbR1Y7sY2VdBJhvTGj0nqTB8bQlyUEtqZAxTAbeTTGrrJB/SwLheyfToIa
WegbG63UqrjV0tT5MTHtli2ERBPxCznVsJZLk0rs96pprYSi61Chp88RYnasvsuA
UBxz3AZfLQPiwrgoymSvkveyqIUsIBcxZ0fH/ppvWjMDucxKDOqSphussvQU5QF5
9PR0gEr/zUJ01St+KFn+FHwAVfSg2TolWzNwfGBxUULinkT+9OqNqhHYUN5bDCk9
3JaV3KlgfSosOEvNNAWvSqjbO8/Z981PMDm5Bg97cW8cDldUlJhHTsMrNA2lGp//
Xb3MIIhWx4Yfm/s3AxkX7lByLIY3JTmLC3O1XOZE5W9RuWZGpH8fuq+6GXCZuct+
a5StfTVB9L1XdaTiLy4hWwqnSKVUzhlN2AbHmKSkVnw3Wc+UfBYvMZUomfuzQgR6
/XzJpV4S67PwyNDVyyc3ZjCUVTePIpjZU0lT/vFQPTZVxl0XPZZ7qAaBreAFkJ6g
nKZYoe0jrni7ib1FY1R/GQ+F24SpKcUvM0xlV0EUszXlPdeXHly24hHeJ7NSSBhY
5czrqddaSLGM2AeUZE2YQ1AVlcCFvC7qiJ37mtO31F/GUZq9Aq6EXns6v88+uaVK
RioVWCSFDNxXc7ncT2PnUo+1Ve3Q+/1hbN06+Xis8l8UyTBqrEF8X9eWpqR7W3HI
Dx0JPwoLDHuJ1VnZvxu6yx0KI6Qgx4kaeYItnZL3tN9mIFIQ7Fgpi6QlxEM714AU
1zgT6kQThLflMkXejCrSF8GgjTqJ4lbLD1xmlAw44MhvaY5d5bwoC9ag18AK0sPR
/fA8VR/34FCLsWysWAGMnS6Y1jFsCP/DgfdZA/fSZWQHhtcNotzrz6IH/+/CAK/x
ZFJNgiDtFPyGcLH0jWYYJ5rYYC5gUpi5MQniCdYTbJjUjEi1Gyr1BZjIHQRz7saH
vEDgm5lOt0w0XEar2WfRVfSRrDD0Yp7SQS0assVjEG5lPLKbgvIC1pmIuhmi7bdo
NjFJqG1kNzLTwE/qpsNaUlTgSIUWdj3M6DwJSPf95/txmLdUVJeoIF4VbOl82xM8
9eApu8skRVGeb6V80Mz1sLLmFVwj41+At13yujnfFXvFat9clL6BL7cww37aDGCc
qy9B0USGeGzcS9nzS6EB4xBkYrd7MyNQKVLrzq1LeCR3Yqr1Bueof9ng17Obp+9G
pitWC52SDylZdnkrLyeAfWvjasmz1qjJ42K0X4iMEY2JhRgfb252ERbarnyW3PNo
9akSBiIF/SP/riJefNxjUO0cYQFezFAcRw2FtKRS+bOoHU+Buv0oG7qSLmbtX9pN
thX9XE1CECYoHmYmwxCFodjNhx9i38ZdUv6E4fBwVAK4atfGMMnnX/RCXKDyBPsZ
3JKoPVGIMwjSbZJCy361rPUegImGXYubD9eShZIEjs6aGd3MU77URr7n1rp/5Vk/
7UMBei4Iplbb6S2QdkCN1/BFxfyggwt+no95WedAwlusBDFglCoAK6TWVP6ym35T
ZMMgS96BvQ4Lxm/4I/scsCu7ZKXhSCWa9FOdpvdrW3vFOE4TFRQQBfkTOFpz7wz3
51YgDftpHr/EM7G6ju0n4NYDAIfAoffXJuvNauWjNiin23dgujsPX3sHWEpIVcFu
qcDuHp9NPuKbMOaAwEYjJIGpF8VacuX1h4XA8pHVstggnH3k2fE32gV/7G8MH5RR
cawGMX71AYoeL6VSme7hzNyQSnJtcqlm4S3qjMORmjB1/Vdz0xkMVa++ZStKFY8R
dpWQcHxabr9HaAxBLHQQ0eczcBrzVOR2ve7TjQ9rPiRCoknJRPOEG53YuWr58hdW
Z9gQj2VZo+Hb0MkR0dP9Z80LNa5j89F1JY3aUxN/wl0T3l0gWFrxjRlKEKC5H6lx
8D32QzjeFaeuc7EQXOhqTjCk3kSF5zwac/CO0uPph3tmIxoIpjgAssUEKWw+kIZE
Hly4kRSFpELaDImbchL0P330OtVscdm2toxctSmWl5CcykwfoIMpsGFutkVDleZ+
wmq3fvu4KnH6+BpDfhPYqytdIx7AvH7mgveWUNYZUuSnHqdbM08NBi2Th7V6z6+h
s8I3dApPZjERXqW9QIFOdSA/pldmIG7Aws1a6aykxLwmZQEQArP5OTYm6Im4taNV
VQioOB3SpK1pqqENwtWFWIXqmN5gSqEQpmGUCgUQazqpQu0KSwBWNSH/PwyTLCIo
JyEuK9+xcGlv0mvBW7CUUtwXShc5k9DSMBE4wtA5IONHwiYILPUDIdGdfESaaqWd
o1teuZFGDZbfgZwZNyBAQJ3wxmipH8pJ7m5XCNtR7ZgxYpuQYxOc3mPGlv5NYFaY
pzuTM5VBBKyf5GH01KeWW2pAxhhGHer/yQ5k2QEtdCM9aSW4SseyTdfOJlix7TGH
77osC3ZDIyPxL5fuKwDoYAvdrkVxl6q+Kc3Z8b9ICaSgcABltJ0gQyiAJpVsR2+8
KMO3IcwzDC1Mf2CbgNdDTZU2Ee8gd8rnslL4Sqdo6UXvLwfPewE8GJL8XRTdRBIC
DQS0p69G6m8pAkRKMLWkJMDGrysHn6AQ17FMMHFUC0gHF6vck7kvSTYIFY0Lljwi
YBQjG4NfDobpv+ks5UYGYvAETUVAc1I3tsJyHGC1rdTlx2Lrqt9enAZ2vfbW2Yg2
cVvOPJim+zV4GzS4jhzYdcjA9Ekjta8YIKqOGY8OS6MuqsK+Ff1/XTK2TcPEfmBg
Hu/aoujpvjomP0PKDZaf0lCdCA8xQJw1SVU4c6LaupF8Q6/JewaqIYMOSL25VP89
PDHfXk6kc3Z+MBIvMWhEQHNMgJgDCduyJYDd2r4FYlW+PF4N+Z8wpmkgTKH84vwE
ltbtIR5BFvpn8+NNDe+sDQkavkkR1sZQQcYhMIM0F8lU1NyXRmiLfbw3WDMlcm16
8FZQtmQMS3yEbSDiUIGvcBFCHCwTBwt8eCt/x0fsZAhaG3JiUxsS/sFN+M8PVb0x
nfl0EQ4QvkXzdD2JbRFMCFaqDifYITX1SQa54uNrsQV8E6XEMntK7LXIjkm+Rvd5
lY44p2pljGB0nEcrWKlxWUmWXng5FxQ/REK5HhuYAaLK3aRzYV6Ym7H/BGqk395K
oPuQ2d01VMhwfmywilYxcCZmTYDY6C7qQASD1yiLFbOJmo+mMgkhCq5Hzgm2b1LQ
r49TUxF3U4ekheN5tYikEcK5pgMG7koRkQpXyY9GgjsT4MFaxMi4ejwLAii6IAov
fplBCoPP518r86nlFXlJ125Ur3YCrAA82SGWzC2O7dOTlxwfWvm7pdLhmUM4oIHS
bMwFtu26FQNLqfpSnztGq1xRRPUj83DsSv9CcKoL4QJ2gTUjv4rZDhtFEBIbbCV1
vjeA15wov2xi3/rcw706lD25XBUUjdv8UjGh0fOwa0VM1VGfIjR4lbQvvG0rtPJn
oxLvjddb81YqBNtFnfcDefOM1QahczBENeqQKe8MWt1fIFv+p+SH5S1HGy/VKPxD
+3hnerjRlMYHlx4tquma3vcHr+5MVpMr93jHpOEkrd2u4fZIZoKXFMka0RQ0sNlM
bwCFn0/Iy4lMPlle2tKQHfxYtwoH+NeOcFLH5ZnhE3lz0K7o/vPvjpVAoKqln2Ax
r7W69MV2jEmqcQMvLLk3hbqaZcAqE5Ax1vO16TIR6usizW1/IYNKkG6sAVtHeq2K
FOc2lyPpgXCJO8p0faEFik+FVujQ068X8Qq+mnrDFdUM3hmXgcTpavGubWycgaMn
TIXBSU2DrL/BZGwgCp+glb2KYHRhAE4LeDQgXxw2hb/sNChUbHcV081hQWiGVpEh
5GE2ZxWGVwXsAzGgYSK2UZP0TN/fPUpkHDjCqaagec1YbLoWyGRY9UpwWLKXUtjd
QrBp5k+s5idcJBsJIFCpQDLc96rTcIS0ZJ1jjI5QRMummOOPZ5l379Z7f3XBFGvu
tLzr1ceawyIWuazmP+KyHfBSiiFEXaGZPXI5bK9pQHWBfFhfV9x7j9uB77l/ChlA
oyADe0deBJQR22Z15FEphKPAhrYNys4y5QRdtRgtZzBE4/7Q5N++CqyU/V1WOOYO
ebMlClQylHh/mXLaMhBi5Q0jBmSYOoYphVoX2oWaDIVNSEKUJnHfMc5eKwqZPpFE
/QCRChnO8R6EUcpzAhkkc43n7Ueti0dEeBIQWjytOheCNSpe2P5ru3mSe2uhazMe
vCms1NB/IUNlnVWGOA6T4bJbGoxsshkmhnYl1SlgSVBTT4aeOxuJJl4LuD7kw1Sk
TmWCHXMuvmoEB1NQruhVqFsHRY1cyEdA02xCueXMyzu/7uWlrsG1Wc51eYKGy5E4
brMvOI7jooVRbwFGG6T44WQ8M64F4dFJTwNknLea0ILuUP8f/y6MRVvGLATxSVlf
r39bU5gGblHMZNEJ+KKM67dq6BWxNG/MYlRhdxsBA8Dv2O9omeaDDf/ZIgGVHVcB
tLbHo68gFQ+TFJjtGbI1YFK5VgR6dC8P1xXWjJj5crEjWTCK6Pgkg2FC4GDkixUr
0A123MANLEvPA0CKbowbb5SYrQiteiZQULyU6cEnyia+C/CGcpgCCQLrs/zIM5AN
LWyrd9WfsSMe8u65LAjD51ce0sRe5LSwRtKL4WldLH0M7ie7IjqWu7AQNxF9U9UQ
rt3ihmkcwPMFvQ3P3e9ucWVB10djXppXBWA3K+xenLaCEJKkFikziJFSak1llbx7
j39n2RlQ9PFj4tHkC7okXBjRlQV67rlPT74rt/34W3OZouMpPobAEWFcv083c8Nj
7nUgI6RSogekh0JdWQ1OdJDcuHF0lA95ffAWKEPP7IKWddL9yJR5XBcy+/4s1qhy
NpQAZcZptOCAzHkgoywYg52QxXM7UjzQ728o7O2tIieof4NTxTp3gCflLxgAoNJm
ULxTpZA+SZQuolBDl9/05SaMPO9TUXe9tJ9NLqTrbdsPUg3NbioYYnksW6T6Vcyt
t14jUS++r2XzJ+gricoDzAD+glRmdGk2tfvJsCc10DKfxlSLgi0LFpKqXopXBh0H
nfqnbbBNoF78GqUg+Woe1WlBivgsYNg2pSg1nhoQPehj3m7kkRlHwj/t0RggLx8I
6f/2mn5MEfxx3cpT20j3WL6wmz75Gkc6RNqQIuNvYtfdhwYkJgHViUHMNO0wUFrn
pv3zkRuSNRhxZs8hS7Lay2v9ZbXDQ0dZgaKrak4cghmFwXJv3npgrrSnNSrL+wta
RQk4GHrS/AwRS+WclgReqa7m6loE0qEj8aq7/IkUeLSCwNSIxAkUeLXEtw8cDDFh
y13Ty+7+IZX1AiWQv3a0/wS8yHi1Qu7WCGNvbM0q31hWEgeuewuikR4x7z1weF4y
lVxKjxgdpPvWQr3pe7tOohcsr/sQCpeXLvFjPhf2REya7OC1/M+JPeePfXPf4Xhg
o6rw9I76MsroHEhpK0S0eRLsMp1kBqgEcppOD80+2ey9uqJymwii5icSeS6I9QPi
aLn9ZJn2jgNeEfokKwlZ52Cr6Gy4C25nZ2cEsHq3Wf8sjJyZiQL705htCmbFgGhL
luef9n71Np07EFbnXj7g1Jn+v+oQVfBo5dfP+uTRrQ4LFAfgC5EEbLPOa6RMcwja
4xKrf0lumSSaBPBcTFqoUOGbwMByHWtyIWCAPeeJ77WjluRA7g+QKrj9nlWAvPa6
jZ4aWGpy7ovr8PRTzG6Sez/VZ07GFTwdqJm22Rcdse2Rte2GYexSglAPCnthUjXr
RYd9tN3gNtKUIaTzD9sDbN6NS2ycU1GFrDuLBUqy0mmg7igMLbFWDAi/IpNi6Hs2
WpELVga9mxw7deYWtExgQGb1bvSUXQ+FdsLXHBRxjqxlDjzJjmcm/Yl9FTlzFBV5
dWu5BadiHf0FM2weGJOlGWrdKfRznacvfv/W8s0VEA/eXMdOpSo/fgQh9+peYDy1
wdGjz2McIHXyFBHPpzmVhq+fCa5h4mZraghLB2klJwLCoOJo5YttojcuVa2rUyGJ
I6IDSXLZBtbbrDWvhNqin5dHh14dgXgSXh0l+CfdIriRJy7KJyx2+1TjwrABfVF9
5Q5kMwrvFPejy5R2AKWhSGX5tlHv0KNm7/Xpvmh3wDpyOgliauFtzErf11OUv4e3
oHDtSIWZuzEfypMzWx+tMPrrOD6jhYr/Z8Ad+T8pmq2fBVvqNFTgbRtFt99TekVS
PVe0GbYV3weFy89lWOywPGxOeLI1sP065lZ5R5n6BfGoZUmo1VbmibaxXyIjAUIb
nkBtS45A5Tkp9iEz1EA3QO3J47n7kRJ1cDM8+YoiiTCXaA33A7naFhetD8cKJ+e1
lWPLjWlAVN7UTqTjP1Lp5QVZF5xh1o2JDwmKWDjwspP7FP/GQRq9dN4tWQ2NqN5Y
7goIFC8W5A9lIxDkj7Jdq6EJvhorMD8xUnl6rM1I+PQtuFRVEbGP8IfdOWrkoELX
5/AMSaoeXGUkY8pidUzZVLn+hdLUQCO4cPBX3cfh+eVqWp8PzxXYCG6Z7htpm9AV
8vhnO3pN3PjRvzZVJIPGjg7K+gKqb7dx+LASlVilZ20BSodbKWSOQ3djOKabaH42
rooLxj1HiEw6aXaeK+Kmd8ImlY70281hs6sChVMcf0bDJgYUwxDsNr0Ex5DueRoz
S6SbLoPPQSpuGV97136vl+1aDrXy6BfuVvcwe/7cQcec3LRc7IPFftdSv5ECFkI2
wZphCCthCPbmjQIR9JLuoQzh+CrPNWtTeGCbawp6u+EAqJNnP+QuBhKT7/psgXnm
rjiy94OBOnSfZ8jlLMo3Z1e5m1Gq591RmFileqsCVIfnzGbtPkvKX87d/E5OiuK0
uED+lH0SCwqN2POyrUGiG794I1C0jDop6T0/n/a3oFVP0sjAgrDbgZfas1Q6ANyT
2ga5AMBKSyC8FnovQFMTQjU/FehBiVTZbq5YTcAJgg0pdJsDkRiuMohMghpzAODQ
DRmh+Uc1Qw+YK9lRhNr+ay08E2N8YQgobJGyZOot/sg7Xfz1762Y9lmfnvL/A19S
qq+w48nWiT82TDqkQ6Ffnrdx4MPj3jmh1fyjWu8fJrOwlbbiUJMtOSbs+rgduCV9
Pg31TSoVWkgQElXxaKFhM4eyrUqEInWr91ujzjJJ9jqVJE0KFXMl0ctE8f4ruz4L
F3gAwBx4F5HUYdZZTYQh+tbtEqb7eF1AYV1L4UlPbhIayKafawtRS987NbeGyr/d
o6hFjklAGr7I9Uf2YH+UFNV99d87THdMtLqWdTreBSYbKpUCodAh/ZsvEcRov3qI
ePex0MCJV5GB169z0+X4mxULOUzJ13uEghbRLo3xfIYQWcnLiVUXN3nxqhlqJhOW
2iWOMxRISp4OIQbiaicR/qkCNiN1eryiV2IFO3IJZbi2OdYZ2FtiWkRDcWjORz8Q
8Ck1B/iOp9aQKOlkvVqWF6OAOMYcOI+HJj3eZtSSd+wam9aZ18PJD5rPUizKynR/
0XrVjMb1tQyPaT0rSzHLZqipI6qSslZiD3xhL+WU6fuNpRD6zSGXOoMi5IBYS4GU
r3qPwYfJRU4ouk4B4QnjjX7NfJX6FWt8zUDcgznrbGj7Nj56xLgy/BLbN7WauMQI
zmrwZHTO4oJcTXiWJI0CKdn5IZ4su1YliocWM+IPnRBZNlhoppz9RzhCHxt0JO9L
txDlAggQsyfTgfDPl19JIJVm0MMwr8XXBMNZ4gJ3Nm9FEsjkQG1q6qDkxjIvImT4
r3wIZVlWIDASLh0h+DUqVy+mEaT9luKljaZvbfDYbf9//X6WK1tiv2Br9wQMgME4
Umrh4CI/cl6iitGvWEudTliRPJZ1jZDMK9fuvMvADWWsxioV21rOdDOcDZVGS0pi
b5xfEhcAhHzf1+sv+6mqCu5H/iqtBYkMtnb8UuWqGnU9i16yPRciwXKKiwZRLxfN
i/jAssTuZzUIk/iC2JDkjCLdvs3DdYGSaKuAeoRSfcVSggBPznIqesab0Onqyo9B
GaYLe4sJ8hw83T6A/ArDAzpUbYJlTMDKH3yh+m75Dr03ATJZeP0RGCVRhgn7ra9A
nFDSqLr1Zm+L1xiXevQGHyRZe2jH22raLW8/XFvczsysZx5UuDTk4jly0pm3WCLU
BTftt6FaL1i1s/3JMqQByIo3arUwZAScOU0/oZ1ZURh9oF3KkWDNjyoeBHdZVK70
5xaQi6Dm+hWhkLeCkg1BO4Wy2g2Ftjh1gDDXAWGRWjxfzET7D0/LpiYh2CFBJrYw
/mRs539gZTdsz///RfTEbCWfUe6sqwRUavXBRV03VXpetTu4FSKQAife6rB3Xj09
tcpLPbA3asAKodWylsQIQkY6fDq8kyDnc/RVtZTMir4KMZWZAUzMVbeWWJoFBqJE
SfZHzrwX2XbA93Me7xvDhjqWq/Zm8pn/DlB7aFLlwWX8VRfXy6sXgnTA4DN62ks2
IV6QTjFxWi2Jre+RMZOXFacuOWW+ioKVP/FL6Lz0vhQWXxxlF6UWjXCTnpQCWWUN
vSQqpdSRfgwVDfsq9kl9eRx029kIHSWpprGRVgvJpPOqdKuoTD4B4pzeCzUATtoH
r0N3vxGy54+LIwIjZR0RZNHDCZ8EsheziNr3SXNlvwymmkosqKYQoclTtqFO/ihR
sAyf4Fyo8XanXaK1ScVdE4mPGrSEPq/KQVNObIcAhl5Bw+jHTJnYCi9ncpMQl8M1
9e4k4rJe+WoihWIO3FDO7zB6QWH+QTFz+ZrmXaqT2Qaou4NBHT+veYo3xsghIrG4
grqq/IaZXs1LL75eqBk4kV2B321nkq5KOmIYqZMzQf/o6/AhooKpB80hD0D1GJ6T
R89w1h0DEA1kdJs3x1++to1b42DgErL5LDvjDxO1rMmYRZkbVEgl/k0EZIw6R5Zq
RB9L3+HER1BUaqQDvQ0xZ5xENZZZZ1XQ/JX91AF+xA60FZou50WjOMdF4D0xLxL/
rNylekoycsi7SGpsoHax5YsLvANyqCW6jJBGshGdwiEWN6PeWXu+5oEPHSnQH5mL
7Uixq0ALRxlUKx3MEyKS5eOR8RR1kSQ4Rgjkp6BOo4n48f4oJCf/tMYsV0DPI4n2
3LnLmnnAVoin8pd2YQp89TjlpM3bu7OvUKUKSynxlore9s5Y9KPOCn8WWp3C6G/i
2u1aMy8t0BbjMf2f3p6Q3GP8zVQ/4MZMMci3QR/SLbiVJlasy3l/NYc3+LwGle3N
XQwOTEvQ0UYb2ERP+EMh/ihepkG8oZNZ8aUMac0fqvSpkwbHYTxzHK4SjBglygxP
WL66YReClnTdhgBVcp34i1HtWICApz5lRbedreJLE84z3sV/raZ0gcAk7qWpzorb
YOR98ysINNOL1mZaDn4DO79nutaAgoogENI70dEojqj3g0UTJD8LomWjptjB2gjJ
Hh111LY/4j13bYHhCeTTzHkm6d6JqCxrq3jJwBzCAPcseqDx/N+wOHnAbHKXE1PP
IvaC5LLdG4c78sbaFe0jaNYtXc+sdq7vPkrk3F1iqd/bL3VKlJCbbxXjS7VhTEAr
EFlqCSVHkdQvIwEYLqyuF1Q29BtITgO8tvOYzJ/wYtfJmTMvee8lqXHlkTF+Va+g
+l1F1OUwTQbemE3VDncYAWfWLY8muVjKoXQbaic7iLQpeNAN7OKe+fHn5cKuxaPL
PabyBd26Tbr7yJPkiTkMGMJv0VoiE/xljOf5DYeBh0xV8ESlPe5mIg5b6aP9BXQO
TB7kZ3MdKr33gbA31tN1FLELbagJlIzSDm9HYzB3HjkGB7sdPaiVly0HXRwqfQDK
/kucguxAijLqptpCzVmFblzCVE9OZYJgESJUwojc4GG6deAY+YAmGiiTQiJGc/Rf
ETl3ElIyX9+zH7AItCCCIXVbRiwMFnGsQq2w939yQCunqkHt8PT1+aAkuYcbSzdI
/nnHEq7D6+ORqumhcsMkSnKxOvvRN35SfkrL7g6t1rEY4/qOopJ/KuL0uYIQdPTG
JWvZ+qvy72SHPRpoYHtCJaz+HxGf5SDzrgrKIDkFtF9h4esARDv6DmscuxrEXiF/
Xu2/gKJlJ9MQgWqybnpsuCzrYR84vbiYHYPJonhcLuPIujPXCYdbO/7s+F596yUx
geol8Lvt5Gdq0RZlNNjK+NgcjCTt9OdNv1N7LKquchIQU4WQqL36RoFC0chbKD4N
xbSCzDSx+58SA4PinV5XwyawTOH6gzQP7OdaWxcLkkBSl3awKrms8yzYAO6dlzXj
TRAKTGyyiLE71V+hhELAIQQEqIz2sgLtx+rcBnz8JpbUP9pGO662l6Lk4+sfBS9i
EdALpJRagQ54BeTP3QLd2TUX7gPcycGYEbncZkkqCzvCon5mvRMGvuMW2wez9Mih
734vfaMTiD6I3Zz9ylBShObcx5SipvQ7eMYB8mFPJv0m8QqqssrHqH0Bq2pBMq/z
rKBz3RLkYJ190MhF7HehaIvasMZB2DdonB1CgaWR/uRof6CG8anc4gEjKRsMsZi8
pgmfxyO509WY5Y/d2BQg95yQ8erAHnkOBe8BuF6JQVvfyfeZ8vf7lLWR9hlzIbNc
m6s8VNYbPtHjiJuZeFGLwTlEHNUnYw3EUCRSJdCGe5Q5PINlch1SMLGdkGg1y52M
jKPP7HddDgBla92frqnG0VMtn8JhFJO/qn74u8Jp1DnKmkRTDnGPm+AfDxPPqAen
iSF2z6kbYSv6QFM7rhKPAdYUrsjJOpqwZII8S1kADzPeZTLix0HFCw+RWY7oo5Pe
1PKzHnqYWUK5nLDN491oyLlGb4f5PUViidlQwTQirQlxhp7wV5UC0RiEWwnnQrBc
Z7B2N9F5K1joGe870abcwA585TVVpVVwN+m/p0MnNFn3OG44bQ45swIZxrxxTGtq
UaF7SvOioNQZdTFMQots+KXq7/E+AXJG6aJXtnXG1B1Sya41NlpIS7mRDqc2u68t
1fVUJXJjsxLsa9r9pXZa1cHNpGW+ZkrH4dZqJv7aa2PA6VhHJxZhEsWFCnagiwhz
Ls/vjkJm6Y8/HuTmBOWF8/z2KRT6pTUTyoj+eXukU4JiNHtYXVH8eQZ8pF3/uNEE
4N1GrEJ8Hq7cgu7mdM4tv6L66FxzVU5QiQmPhaFGaUJWJTMLa4HyQ1nOv2eJbT3H
tKOkH6NaHfDwCV0O5RUBnnOuvXzwcYJ2SqQd2u8LkAcl6Ob5lwupzrcmSBwxH+CQ
IZEekD+TZSGX/nJ2GEGU7vypaipFnfAKtjmo7IL08ntm56laTxi4FgAwmE6kkeQr
j2A6aTPCmAvpXxyPGwi7Bdcjkj9QZiXkdJB1RRP/SWc8B+NpQcnnU/cx8dQGfxrH
XOmr97GvcoelB6fF0Z8jF2njgKEEZC7odraY4P36jXwCo9volYX28Okm4/WNg/IV
7eOe4a6fe3XVG9dQ0uyV76FPuCouSmKKEt9lK1YpdrqhrZmPemn/e9HjeHcugSqJ
P3VdqOIl8pjimj873oVQy4mh2sG9Rcl47y4t78tJwzgpN2q/RriYCYY+bgCXlofT
Gw3RnYAx58K7FShqvrH0F5RnjB2wFJM5Oumycnkj5zKfFVncCJRWp/Q5dEPOFjHQ
ZkLZXi06tyCLzqCaEAYsBZSZbvBtBpXctOnbW3avycQcTM1gTKjbvraC/gALFTN0
yizXx3gAy6uKu11hGXg26DBG29d4KcAKK/ybk2cZwEICr4ntJpwHVyy3jlxLh8vT
dxS0f857inxh06VKt1skkvKNrp2RDrcdPowvhVfjeBXNDW3eIt75XMU1VMtjRNKT
WoWO+Ko7QEgmPvMVQFpvr9BWcUJX7jKiUxAun3ytutLLnSKMz+jMltoFrZ/JaxS5
ATVIEO6WCHFxRwbTLCye4RsSCkosZSjFefMewh/rfgWebSDWCI/2P/EEeHbUn4hp
cRkYd6k+D1/YKsIWEW4ruSjaIvLgqQSUZvwDCXSvZ6SIvdhcnBv78ZJjB7j3D///
HZDArkVHfq0TDXmpr7G3QSMU6zWarIL3832N8tqUAmfactmbZSoE3pFXOvM1+hSS
Ex4/uKOqKEwAvowwY/avSTSBA878VSvbN9+IoQbvgwk46+xMPe0sPrXHYJ0nKsVS
eF8ybfPFqLKf1CWUS8x0T6AQvtXWQUd29VPf0afTNgwNVlk13jzqwNuTA6mnaPAw
mOMAvjJuIDwh+GF2CCEshFlirbHgtNJPiUPKgXeR7SIH5+gmKqxWY921oJsRbpfu
CPvA3Bed6aoyTHTuA5VMkNs566QlfmDORBkFqIWJOZtD5wdAlYMAQ9uPzA+JZ1Q7
oTElSCS3no/tNP8HCOyVcYQGKos5K0yyzGnAxymuvafcVqoS+AxWp2IOQmiJe0ZZ
f2zAuhS8Ge2p8denqg66zzbcFrg4xvmmCMfy1qpQ9RqooQUfrsf80xZhQCHJN/Cl
+8iII4NK1XTNkoufhIIvWKpX2J9zZo7hHHhFpUn5a2tMj7awARe1SImJJVaPsdVM
oB34UXKPy/TMaMU67iFgyiWXTSMOrazjVObSzKZuFHfHpr4KzVY2lLxBW7dLRG2a
saaW7jSLs4i0X8d2rd3a2kkzvpxEEJ5NeBr044m2hP3ZrAxRrHJTl6vFsy07U8YW
oHFBrk7rbZPGJD9Iy39/IoPnux68u4W62uxGiL3x/l0rfiMTSZJ6wjs7Y/QVa0wk
7GgRWGGobLMtTQUrVoeTLcUQCZOUAHfw5LcWsOAJKGGPvZrfuDhA5BznGTzYlxIl
J1+TxOjgqy/qBONQay5X3/peZFxOCoa/qZdKSTTBcXy26qkbh1u5/70pY6qAOyQX
qszECWKUCPWvhDKEZOqjVk7xB4o1jSQdMEyqVPgoaJ3G+ND1jpXrK/2kFzfz8ojb
kbnXkk3FiK1GhlThyKrf9iFBjqqlLMc4eQPkOUoIXm6wxk7YIKjq0c31ghm8KJSp
iLKB4UAZQ4PMzNs+rE4Drcl4Q+sLMQaVhhDdJdFSM/Zr6cWg/s25bF8tQBI5qFlf
s04VHWiPUp7qFmE2scb/9lzDGdqV/AdxEueZkth5LMGloBaQkq6IKY5EZeUuzJYB
53suprxIxG5cK18ZHvZL401GTWXcbhDnywK+aZ69z8s+bGoCr3TolzR1TgQRITvC
7vgxHoV9v64M4YqfJB+ECf5sdHBUyZwBIswgDQdH7Cy5LFzFfg8ez37m+No5LTip
Opg61Uoupn9NtGRoESGMF+V1k214jc11RQgnKkGIqfuuuE8yjtZbak2MNNkhqNJc
92wzuwb4MOw5meclOcxC/N/IyzkYuah9Gjltb3QeE3AQ9s//c4SQ9rC7huzwXhqr
9hDkApALApTMWzje6fPZ7xo+8XbmCRLlBMggjJ1POLgzH/NBVkkMdI9z7Io2+4qj
pOCsmbPrdpzb7m3o6Iulg+XUVaUj79NUtTO30XGOVZifZ6B1o7UKRtntK4eql7Aq
vETPCcug9hrjRvGPrmONRAgqlpA7YxAdvTMjXiEqo5QKVcJa7pYpAUme8rMK0vDw
P9FCCrglZ2+QNPYudVc7mCkyh5nPPLhAp/8t9lczRVoUll/2xCQhJJOcUw2ycDv8
iJX2jubihjXQGWg+yR1RryyMhGfL8DoB3DkA/nv1W7QPeVKXrQFggPF1+1zc/qC3
4SOkVFnEPL58arD+5cgXYIyRi4UjLO7jtYBb4uSLIjVwU0ivSHHz+4Zu8zUrkbBZ
A8eNx4QRiALAPL4PzXr2yfxgNI2eziQmL2om3fVY+y5iJ8Qn9WS8FLaD5iJIVIRH
VSC2M0gEPgK/wStOdM69WyKA9bzfw6k4J9gMRdSGSOBVh5NqUnAFbbCN74w405D1
4CZsH868SrQFUcfNcd9joM9p8Q2xavJt2n1UvLZ7gK+qw1Vqa8NUiBku0ZNtuKqH
G+mSeeQoSG0lVUIKxu2y6+qNhkU9izs/mWK1/wzP2se3O1uJZ4L4KhBhBPAAoaV9
ZeeWulXpFvNeHO0A+62fx7L7KejJsIu2vnWgDg56evwpoYHyiV/1/siHhc/qvMJK
mc7ikjm0ixQmZVENz/R63wTG4YSuzVw1wkm4ciN9WYHb1A6Q7dDxXGjO0SZRM+GC
hO0KPTta71GN5n4xbWL3agIhb0zfdfVhjbigDLoG4gU=
`pragma protect end_protected
