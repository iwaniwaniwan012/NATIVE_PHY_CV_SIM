`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Aa0RnJ4p+m7b0qdC/KRYoJvP1gnvnVJEIkSVhjx6EJL2EKSkDLwcLG2U66jRXXIo
d3ASggIR5NIhM6oJzTZ6/l/Qv1MMlv27R1+sia+r8C70QYjSYj7oD+AryJbv8W/D
++kyT+fLRrDCyd1exscD5bY2bZSegKgyRdyYeFhGKlM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2224)
+6skg1PmpFEisp6q3S+zdCRy/bhyPXdf7ciuoeu9e/E+5Lr0Wy7FiLkP/rUa6uxd
6369q00RHWK9mxA5ht9Rfg/nCl12VoI0Xrfq4R1fEXX5pbDQe9B+yQUUiFPhEyLT
sL0HFCt8Gy5K4sPC2o/B/u8BxCo5VdAbQk7vzDoXQu2bl71vKAdq4DxtlNg140PE
LW411Y2KNvk7zxCIrRZDb43f/r7DhbdfpTIhdHKAJ5aMBUjKYhK84LVTMcWqPtrb
6XZzD8Ifpr44fZf4Ox+vfLGlDLAB1Xjw2TBlDUv1jBMu2M5JT5Wk/07rFZGNz2kj
bAKLRPcNhFjKRKQRR3eXC5adppqq2iahvX75u+0UwbZIVpQWWBpinuEoBZwnv+ON
3g3repQ6yB9zaw/5NCjosaJ0Y2cDQxH1ZUBTm7YLIBlRSRpo/wKsqZ9YQHuZKiv3
SX4ORwyyvpnTKj5TN96NteGIUPg3eYL8DHgNHgZxVLegHwOkuSVeImlQRqENgflC
FERriOodL/5s4vwSythN6fZn28oWLLquYqgKFKrzJDHFUAHp3az2ye1eOOeQ9hYm
6Z3eFX6bLus5+pzMsfTR4BBqZTBBjpqN9yoP6Q2oZIPpeDQOmNzZXfVciEZinYcA
SKdvNXJItx+uTsglVwW7FDBvg0tZXMEpt91LpH9hW8gFiDcZn+TK1inQ3cSrSiW2
kGoVCzzFmrHBHWCd5H1nmQXEjVlhyTdSdon1h9tOuYjPLSJ52GLOmLUxX0nRk2aB
Rg7FiTv8lBmPMkOusnQAyFH0fHtWTt6jifUlVCTd3Bt+5JmNdak5UrmgLZyk64t/
JG/vTXbWAR4MPNeSokKgWGoBNrOb4n+kq5wA8NSIz8wuMycZDMSNpXz51Hlbxiwv
+OUPbf+a0jsiOZzqxiLp4pYDJ6l9pOisKV1L6C/hVEL58pvOk99zOHFQSCSu7Ak5
+xn2BSHJlx/hY53Ku/JsIbM0uyGaV/4HNcEA/pKoai72tB65ARJlOSprspK+iXJe
UzHskVXaYpmx/W4hxODSSgioF/KGrvp6SEY+WBrYKLWs6v1H+TXCkoHTZvbrdt7n
/rW5mLWfIrEbaSQTBHDA3uG7I8V/3tkIl2VgqAE9VbqFaGtKEmWQ7yHjJhXJ6LQ5
X5H1TlUx2ps0Qahoj6la9z2qP7mn3+pakKxZgMXfrB2yQreU3S2l0JLSmLPzsqPe
63xej3Hh+pRFcUwy1wlfAjokxGHcGKACWmb2GBlKGKC/i/u0d0kIGQl5TJzo5q2m
phbfGNkY+eQWHP3gv5j4oPyrd1tdxmAu2duWksedymaoZuwBvAVwiOZNTE0KxtXJ
r90UALKE4ui8hEMlhhhaYKu11wJeLnepAlNhjYCKCENkSwNFxh0ct+2Z266KW9Ix
sYC+JF1FIRUeVPHNgpQ2IszAqMuT8TW1dl/0nrJ2w27PgLX2SNjWH/aoUKxPW33c
juHssD6iQmqlmXdtj7oTFQYX5+MqEKsaXxBycHMr/gZyg1L1Eav4Fx1AQuz2Gf/B
vtwfxBgX9XdR3oMAioUzlrC6xWDfN+ruf8Luu+vXj7uXgQ+YrDNsmaWfn0+nI3yZ
ZlhSnLor7bPcXrWjbr99aEgxuFR2toiSDqGuMW/Y/hRSJxG97Nbao6NmreGdTm04
FpM/BN0wu+FZ1lj+hkn9GKJBm37cTjn2s49CzQDsuAxI3uc8ZnuQiLoZ2DucRzR+
09f19O/Ucas+mPVGIgNgOVO5iQw2Ss9A+jwTj8RCJIWDQAatDFtJzMOCLN4RwJWF
pyK6CC+5nQlBAxB09BcGp+cO/8Ix/TOajko6+QaFQWlGZ0nMop/GzmeQ+XDQupGy
ixLxUUgbYIXa7S7TRAQQEYB2jwPn21aGYuEkTevbuY+dmTJSCda0pFIonQKcvsax
WUYOEEhYtFRhkWxCRKPB1uZaZA9By8wKT6l4vw7tiBnwtecZjzY62dh2MySL403T
9EewdSzXl2Jj+1AN5Prb/pFThENi2ZEMcyGb3qV+XdgkSSwKkF+FFyl9XVZexjai
AIIzvdFordOD5zvHQNQhg8SyxteE4IuFX6NQoRGDvhgi+dHcABCcIUjAQLFt8TPx
xrP5DhSZUjMp2x/ZgpPjx8WplIQA+RoRicynBPN+fVQZDaChwXabFwB2CR7NJUv7
c+0lbOSpMU0Shm9XL8NDYC6ypzuzoF6ND7nQl1/uFWmxpcxZ/YNf1yA97OmOFjdO
Bxdz859IxBL0B1Hd6hHIk4E78aiptl+/ixF6dfmD2sOwijmNxS1bYT6iufjYmvtY
w96dNFw+RSf2Jk9wO2o7emNjM6SVg6Tv4lJK5bP5SH1dK0gXTthGnIPJXZ9Ye5UQ
wbvBhNVGc1zP+Od6y3ucHrQWdhgBubVsw4p/LllcGyC/8qeUGS5kq/gRv2//mVse
dUhyaW/9qmOE5P34mjKF9EGhCxYERWh0FkmhcC6xFvcheb/ThMdX7Tm2oGIZN2g8
uT44Z6j2DpWotqX6mnyOAM3dFv5U1ndJ+7JRaZ1UwfDSZOyizGOKSpJ5U8gBdPY2
UFg7aDTmQZDOibkYlivTBfiqozlVS3jXTIUB5711wJLebn0qkQwGxpT69pK7PGbD
WtXk/td3/SXJnwL6fblXsWUhYMN1vX+h8qQnwab6aEHXJaMm7twM8JkQTYslCni6
640o67Z6xefwFxDqiOsEa/HnGdVBF0VBgeLFc/sj9yjuVMN0BYq3CjPbGEg8XcE3
/R0ybfpqit+lEZUXUkBgIRRqOu4cUjGceU61OoI97T7Zy6yi4VvQ20paRwz+qQ42
Aey18ngiSQMjXI00bv4rKHt1tngMMpyYuJTgP/mK2xftz6CRTytuUsckjlehB0Wa
8lzkrYt/b9wVVKB9Cm/GRrhQA9qKA+4bg2++ubvB4W7IYJ7bpgyj/tZEDnGLnKFg
+9pyWIwKLdYSYWEwlyuvqw==
`pragma protect end_protected
