`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KrpIDYs2Je1DAb063F4pSP8vpgDWxNXdSBAinQuFALFO+H3C4BhqcbwpXpz2fdX4
g2X3ZQM9e/3AUjALWhgXkDHieCJcJCqYRSKqPwXAY6BsSuI4htd3zkDr9/MjBPmq
C2VNqimp6tmKFLyEGiKR24ughEEkcOknAQgNXbFz5UI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6224)
WexAmw5rIDPAHHrTJTOsaXTpYr8iZlKO5dXA4rjU7U8ZwgbyYYh11mutb5VE34x5
AIyNMVlXz0HU63vrLDyI9/6UkWTcF7roPsjo8DgEYT7U3mok1af3RBrZr4RxKjF/
BAY9YCRZzR0Wia6Lo7zeuwuDCMmE37BTp+4bacCysL85A96f5FSGhgUrzeve1HwD
esbn6f4Mtka/NfOkAJDdHoLqvilBg/3E9t14/kmMEb2WgeUyKOViLe3pvX9HtPy5
WagvQR47sxN7IXqRhBotJ3jdaOKjUE/jF35VNMUPCeYLionCT5ZrhWJqclPlpFwg
rrDjUQcedG/qfzLzJ9gonALUjIvEDud7RXUYBaw7D7gme4BkkSPpsxIbdOTC1rsk
nX8STIB9XddiVW5J4MEcmdXtN23YQ5xtUPpiCCotOnnUBostf0hrT0zqHKMJRhM7
uty9ICfLv0sZiwBNgPH+93MFmeSZAmLDmzhPHmL7q21HrIXWYZWDgOvIS6iGsRdt
0CApOdDv4sam+pdut0EAQt9+0IfF1Vz+h09WxV9mO73AWnpG3teHogg5DGVt7z9q
2eEeBhTmnj5ajFBIkKK1TedQhK/b9Cb09s1p1Apks6VbwodNQS2Ea6AWG+lAk7EI
yJ9DysTOWCEOzw7AcpSFolMvh9t8cKPxskjWfGXsodxMAem+mFDfxjyRzk5yQ+EV
bnotyG4p/wLjjgK+ieI7km39myzD2ytKXyoIYTead76qR0anQcoftMVnomUkkmNm
aG2Cnw6PzHxzBcD1cLYy5y2WWgezJYaBwsWGTNZiG2ooWR90dRUWsxTdiyqd9eF8
9AcMEdMltHV+TPwvPyWGv/MhJUPmXPchL/hD2jGBPcD6L3cN61w/Se2XMEBbm35A
BZ0CP0bv/XWOnGgPF3OxGvFcZXYiQIytSboKmuquM2oe5KFWPvVs1+NCAvf7mQoA
uGVgYSRWv/eJaEe6cRRtRNmIxB77a4xtHI8aozmLHzAPkeKsgCjLJ+XEIdzIoLmo
mnxuhU7o/CTQYBU6zStyg52PljQBoq1WO/FD3eLRWR/qrKMPNJfY9jFp5AOKmVzR
A62S/u4/7zHjd/dxo/J2iNofshKP7KRVCyee5SD7deJi3nRWzeCFkgzPvVI+k6QQ
lKVQgk3PIC462yT+p+tX7EvZN0Vn9CcjPRTfqLIzsskdHS9zagsCWcPnIe8ppv0d
gDD1NE1BGcb43kNKw6Su60WE5kUP/m/bV7LqXX73+ltyODZlEXrqhIgDRDVeJ5uV
opdQ1LLF9YOghAazpKTPILDM/vnE4MuThH+kDUSzXy1P2smDo89V0C7poHf5RXij
BvDj/gjWpUbCtcywFyoEROhuePV1jyZM0jmCvVZKN5Fkb2so7yil4e/NAkrf7yjk
DCrm23Xjg+X5+wG0L7V4OxUpGbO+T/ALzfoctOq/0LIOeUKIuL/inP5Ri6y36KwY
pQYfYqwLtiBn0OD0KmnjeRJqA/e3DO19XCvph5fSGCGsf/DQO81Oc+URgVshEyhT
vSjjCg4A2rGj/ykGLhaX0V2BY+UyEzTYs+W+1YXoALUYb2z1nkb4Xh8StKFjQjEC
4ZN8VikZdnegaDZTKmzLcA+mGSGxugn4KXmaWG6ninGaeISx7fEpLPQNqjNBqCIh
sYSDkgAkmvnxNeYi5/ctc+2rRck4U28EDuQdv22l9xiwYFk5wgenN79fxx9H3dyq
WOJP4DaQBjzhiLtT6rAWceRrfUxJFYhbB7GTvw1U3/QhhlQCkybkJJsq/AoIgDyn
RsQgNIq2pG0BNbcsYBUmEpeGnr5u+JF83GKdSL0ww1ukqU5yAzreWzbEMKwcpbmY
hugaVMxSlbOTVT05pWf4F2i2QrSSPsbcLNfVPpBQih7dM2ltEXZ4i6gtAYsyZku7
IjVBrVzoq8yg5/2/fc7mNKgooOa6FEZepjjGjK5zwxnWH0/OkKVRhSyWUxKhOVxi
kvk9xMzxIsSWikrE5Vgof8OIuSbG2CTIOwhyECF0+TPGu09m5FP5sgKSrMirqv2a
j+2pPwyL8LD5FCXyllxBXnWlKZ0MV5KAiaxRf85MqwePEHNuftsvMyAwYK2uwzYJ
H9JBvJ0YHq8QyR1noYdj+oKnralPeDUxF601l+HMOWVG09Amhyx787HWXiblgut2
xmskOmO5Xo6wBlNV6UhxL0nR4YQn60u1oGRd+JTR4IIQSlKZ2BcjiUw0YVPaqJ1B
RjmhsuDGevmJ7eFJrnhPp4zdDQGiC2mcgwFvxsMFYaDIGFn/TFERliHDDSFixL0m
faLhAbsuYTlqSMCinH7+Tb+OBgFp6SJtjgyXjvfLQFhP0jzOOS3BGx+vBE9FLgJQ
hyd71Mh9YA8h8qoQ2nQZTRboHf/iKEAP8tD+EPKuNqiNlJefT2rLPMxHWfCvkLV0
X9bTLviKI/mnEb5qSpKuKTGadV5hdtWnuBi81NJBdgRqpajcy8jXU0CJ2aoTxDx/
LzzNt6B9/TIkXAX5+tk6vEzsfzFtrVmttQ0+gNylYVq/ZLNEnws+It24L80SfvQJ
1NpqmSVyBHLqfX2zdc4bMyzP04DxsFyXAl8c+pHNAhmLGSR4hFo2A0UWfRS9wv47
T5pRhV9IJHGqMsq80SxoFa8Z8/eFF/lTk7hMUj+iSWZdzdK/RWs+3wY1Sr0gPCc2
fQ7N7ewhbygpZEL4lY4sGgqFBubUT9p1/BvV+4ykFK4gtGWIrjeRZIy9IsGYUG3o
yMCn2OuMELbxAcl5wDQxtU3WLDJ5sAx0/7BHc+nT1KmJiV2mpSE79B/crRsUv+n7
6njNgHf6PHdzt5iRuRrLzvg2aMagLynCT/7nmm8s2XJeqLGIgvYpTkFPKZhc29O5
sJ72M4FZFBBKHlJrmU2DP09txzjxRD8B2xD6/voVG6lJ9qRfut5vcWXA4iBcZRpI
cneQ84eQEkG+3+Us3KSlRDCdg8/ZBoa3QjA+z1aY6VQ9ai6xup4DophvAaSiXYKy
jlR/SZncVyztuTWSyNmTfEhSclRu3rvwL5pqTetzxWE9fw8EQ3L7j7Dm0Ef+VKXH
ocPbZkeD/3vZKUt4rCCQCwZ9BJn//IdZ4IqXOsdTEx75bveHv7Te8DPAlh6MRBm8
ZrWy4Acm4u/JX2QGNb3tRPi4OYdNYqKucBTzuX0OqfjHWVvjx64evLrBkKQ5nY78
A2x2gAKg3iCcO1m+qnG2M268QkjIW0qCk8V4h9B1+o+F/rhaPjW3+ODHu0Fpw+WT
V7e6vR/kmxx/b0cfPvY34aJwYTxEk9XqdwtU0J+eSn2xK0BcgMqIJQ6O3aLtjXRo
82DM1knTZhpsTkeGfnphZ0P8uUDnOTyRwzJbU8650eA7ccW0gPBYuomym9Rourhd
pguTjp4XhIXoBIjHTtG5cKXpEBteN/26VjZ3jjQBWvt7eLDL9kxRVzSDA0HbSsh+
AxwMxfECi1+zdHY9LbbFHKYpAaXfn3V+zTVPgZU2+miMljAyYx4eLz+MgP9BGJcj
DyW2wQqhZAGyk2i5sUO68gYfMvQW4gGP9lvLZMaRPjMT/oJkEGkzaz41g8BOtMlq
fBub31wJLw1dq9gj/v89RjgRT9p/SwCeR95U72BmkPHoKm3IMF9siDO1mWNeZ/dR
U4GERTLi6I16sX41sNIMezQeU+8yQ59CwgCSdABvHLCKBrnKuV5LMkJ8lJtrNU8X
v0QoyjrHFJQ7MB7ANqF60ZGtObk35FKwmz3T/DuJIYGyNVzqGRQgLNAJLqWqkavb
xikEA6RAzQfZuTdJzmqyJZ9aXTYD+8OrtJ9F7csrK+RnE804KS9K4iGt8y9miJZX
pi3ywczTruoLd0Hyp6rEsNw8lUzI0hyvfmgnSgqRKchw2oXfVvmavcOnZ4yQ7CBc
R3g07ipENQD/Nv2Y5CFsZrf9DYhMh2NxwgWMdkBYrGptgBh+WVDAkaM7ZSqHsuMw
R5foRW+POqKD8+AIyulYkpmez57/8+jJu1vqrBAGwENJ8cT+K0yj1Fz5ZglcroFC
+7M5UKp87Sj82Zzzq+JXWXzDX2v0I5uYLG4ASS1pt8pMoHQ1lGS0H+MNocY4YHyY
yPcUcJCcgIlah6aenV/gWUT8Qy2K2TE4NJDFlz61UeJc/QYngL28aKkCjuveR0Ph
og8a7NNg6q54AySnqmP8n5yBFaPlrBsUvrSS4fHKRQryEwHsFgfUqFq5fcOEsSkl
XZujV7rJAl2NGqTY1XGTWdPdMJqR3eWjZgLB3NknWFtiz09UXXjCrLxSObmVqA9p
ltut3DquCSvy2aP7NAD4/DXQ+VEfPwO8oAEqqDNBpCgeI9ps9Eu0bxS634Bns3qG
Vm/PJS93UMdRQI1osnyvqCaR66zu5pVNTi+RlfCywlaqdfMgnhOEbbscMLA7062W
UdZrNr7ReU2mOYtlNQ/tUZwnfOXqq+g5FpgCS3VVv34JBZek7wdD/r6H8BmAeGl/
8alowv4aH5AHb3UMc03lGtdiw934Lve1i7PdMFUOzQXPI5ZraBBM51McaCvk1+YU
dvaMMcDjEvgfPVQ55tW+Ie3E6on3/mt9xTCrob+QOUFDtRG0An48kYcuI9JAoMyi
h6PHlPcylUDg5i7n5v61E4E93bIUswp+fmql6idU81n6yncuRY6oVy6nd8yaGCd/
raFbKyFSX3olsmdyLmP0oqO/wB2VqnkkeTkZk1CR6dcF7T/B4dJXwEZzfap1Z2z3
Tt+oNplbT8n/UdbqyrX2kMllZhwOvAX8tex+DqZUkMcENmnMkadg0P46w0sYoAiC
1DWcQFZdiKhc2jknUETEmFmG46HgB1+GARSVQH8pB5xq79xl4VjOhdhgng31pFrp
aru5WBf3jAuKyggMKGJgaw8grV106Lawwxs4SAAzf7c2nE5ljyaudmH0s4FaEQ6g
B0dMnSCRoTRWQ86EmWMHnDXVhe0GQvxojVkcWGjOxKPRSyyCwJjeVvMQJCOigUhA
3ZeBdmeL9dL/1rv4VbT12En/4l+vn7xae/xSvWMEDaIWXpGZnoec9ZUfLVs/he5y
QJY7M6FOUW45AvTO6hsERFh1FsubP8pV/moevGV5dh7Ahd1wtYBq/RNpZKA0Cv0N
TMeX4AyAUNyGP3EXqSRdKwPtGd0cHsi5frDdWoKZ+0T2xgagSRnzT6MpMRDVTIog
zV8DzW/5ViyqvmrEdO7pn7Df0BsCp17mbFuTSsURXEhYgKRkI7BDNLZNowSRDC9d
dbbLp0ygS+EqeL746L8HXXM+cUTUEhHP0I9Jwf8OSBEFT7cmXhdKEUgOWtl9X/zE
V3Iv3kUcDZ9wvxvp3f/Bc6jcGy4+pQxxwbUVyOGm01s1tiBm39jqoHupFhqXz1/U
QPCRJ4gJNcxiZLwdpWHSIpDRc6+F9uU3xuEEHAL5o3RQd9l5cK2EA202ZCKK1njJ
QNlC1D+FeYxI4xHeYexT53YMJWjAow3tv+YDbQ49aiN/lzRr6J5xxddp24WxaxKF
fD/NcUAfF7sfbkk9gpXOhfNp8JSt0nefjbNTtF//EEyEK22th6vQSUU2NTkbOO7M
frIcqz5Ck6CzQYVpJKi6KMBoZpT4JywnF1VNEFVfFSBzW5WPThFUQUeMvbDyCSI6
PWQSoexjxcTqEvi1NUCMXv48FSFMDPQNHMwE8B6ljmDjXJKJAcYhR/iaxSfrNoz7
IDDsffxHVPxVUjjlSz7/eKx8e/zG5dOS6pSAdfi596dZaaht2ZNDEiBhqgR0P7O4
Q6Ez4ISDTJRVJ3EiWfBQ4rwQkamVzHhfp/50JzWCQEuhYQOpEYp92PHtBcj3xKHF
FH9TX0EVucNBGrixiQUzrLVZP1Fm0ny2BAzkNf+U2BAa9fQSmQLE9C7omUSLWlO5
pB+pQYgV0FhvQMg58vN9Dwo2S7Zd1vMBG524p6kSGN6UDOvZu2E2JBKgtStpG6nx
dc0FMiTgYGbXDElUIq892IHk7ilnNCtUEt5g16lZRrDoO8w75FbEz6YhGEAQjAvY
illWdRE5XKiAOKuzHyiCFzb+RDWv5n7p7D6oI0qpAMuAvufUSgQLnSLVWq6b2LhQ
uHJ8zcgz1DATT4QDH7dIe2+fedxZAXYmCyUYejJ/feYbNdp49vBh2R4V99dhF1O6
OCuc5lwjRbsY51Ugb1TGoMGFZLVYXTHEoIVyNGTSl7XqW58QFFALmrpn+jeMp9Ks
7wk05NmEe+cgRElDWnOqcKI4fXkcPmguUQ2lJa6pkOU6owyrGyrkjWsAtCFAeGey
8wUMEmurY1pBUS1SLwYxSiHNdikY2xfu2Sq2qyLb0IhLNTwUQCzkHzFB5WZz7xaw
cNUNeW1BdUxOGWbJJGFnFsiKWXct53/+PqljSxjP1VhzWGlYmba7N6NiWcvBHRg0
9tli8va4N5D8NX2/H2E9Vl+ZqNLAt1yJVSHb5QSC3KAUYsHIA+7rHcrmBDjsUugB
emCYV5X/jA5ECi7THHRbWOds42TxCfdTA6thQL4ZspoUj+Ayv8Capws0AUKhvVHb
RkOIj76jzGhGmt5pdL48kJTRWIPrWaAvqAPpHmFM6nAkNWaLdN9iEAz1/OROLtc3
KaApeYM9CryXEqPw1CPr9nRajHmKHEMuOvsay/3gs43RyMWeE4ala+hZDwKlZFo0
7b2fc+7Y9ZuVMtcSHBDWbV9x5b2OHvj5eB2ZTsAIto6EszN4WToTwEGQ+TrFi22K
pip3J8t6j8roFTUv5hsxI5/yMzbUKrRKUEyF78Uf+LDh0ClOBy82oWn/UjFma/3U
pXe2YNdFvSfzTNppPfJj8Ue9ekd5BBgXToDKfuAHaOqlSIUuasjBGrVw4bSKymtr
sYTOo/0d0LT4veNbhAPnDDY76yPLHLqlrrQleRsavhwmqNM4CbpKhHTHDDCYjx/p
9TFMJXxF1p7BBiEUJbK9yJB+XoItm4y8Pp+oJVMdPsW5z4xOkun8vXdJJw0QeADa
O21JCUvzeP+t8Lbsb/KAsuWECWNqnQWaFWk3gAXWKtd0zMSBaSfY6mDWVD8tcpnS
gw1HbtKE56boXzpq1FZZBAIeR4ZUNtdvRndf01I2oCEP1tvhMT+HBvEDWApGiJ1W
ej6Le4Rqx977dRGQ8CK6l55l9MoAi5vDWyMPlfOE2ykGmuG5QvP8ZY+Z3o/yr9Ib
tLnsanPgteK369fdtuvmt5XadCtYLBZw2qlh+DlAhcfwjWLq1y24t8hdwZ+XZjp8
M/jmVunC0JXHhWhO6dqgBGh2YJKQzbck6ZW3Kj0Cfj/OwHHUXmuZra4F4G7DUYoH
k932osLZoJBTfYf1u/ECLW/v/DqSB05kz3qVZJEzBsJpllMII2iOTJbAv9Vppsyw
Ye3BIwifcJ6QkqbgGL6mHwkd+Uc8WusLPezukNXamBT9HmfLvUEae2GTPKdwnFIO
hEGnUj/x7ZAqyGSIJeOEjCAdo3ppmVSipuAxutUTZMYjxMsimQo+vO5Uq4P9I/Cm
w8S0+JG1VAQrvwdwoHwtymf40X5KfuJxLbHJ0FD4kt2ZkSglMjhnCpU2CCKtHLpa
dmBGMQBfn0S9LCts01A9U3x/t5z8zb1yoPSl/x+OTp6rF1mqgBc8ZNTblfg+EIfg
aDfjKTQGYZ8vBndDxDtkO4e3flnC0FBWp/zJw0Py/kR+ZTO33U6v3t1yHuMklAqz
+ImkObb48G6gTnRwjJPIaljU3WQ3Xe7DtvrrmSuk+cE9kt7IiwBEfkErI2A/XlcW
9ZxYmxe/LIe4RU4oL76Zu034iUIiykxc6fGR+D9Eo4LuKMOESoUPmcs8Q6sEjpRj
ploNN3VDlYe4uW2aa2JB8AsMUIMpNEqigBv/J7xjfDCYc5pBM8MDVeXRS60cDf1j
Av96/jMWeGVKYnNXkufo6fpq+x9kOeixNuihed0PPv3CSyoGF071zc5uy9E+Ml39
dKZzcaZZCtFWR0S+QlUwOweiQ3J7bmNWJHe5pbKFPAS/kjKqiozOvi74SCdV3gp1
2kvy540BYkcw0qQcnHHSXVwN1hscYrZU3aApeGvd1+4swKdLaHHarZ/dwa43b294
SATXCuSBQdw2vuN5qX8Hn27KHwr93sM7WJ0LTY9KmSkTcxgJGhA8eht1HzuZaV0x
iUsDJUf8G5blccD6LZV5V/quxtX6j3nqNcl+Ql4zeiH9aZ7OIbfQw8R26lGjk8TJ
33kx3YYwm1MuPCUhlGYwN7RiLcakAAA4IlAJITL9bK0IsrKnPgCXY80NWzmZVQJe
vob4NT3o6aMTC9WoPE3s0ZmjSPy6kxAsSX4KVhN0UPY=
`pragma protect end_protected
