`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
teHMqYzFyOvxVirUdu3wupnRGMpHU5bf62DCMYZRjCkbH8NB3N1Y5DZ/hPkYl/U3
cKuDLtMFKcLFnlFd7KOb42Kkj6XQljUWQJcBrwPARSJnadyNf13DsHGZ87YOasFU
7agpGxagsFUWQSdkA03QYQu9mqiLTPkQZyo3rS577Bc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5488)
2s59vgpue77xcodiOKVyhIrj0rSkfy4qG9bFuQE3UzWeywzOrEtbsRDcOidB85xM
hvnhz+2C1Jo4SIMeiVRpOqod/bWBFigiWa7H3i/4ll+AHrrzhiw3+LUyLdPDR8Hx
WJye0eA24nL5Tp/kIych96hlEI9HeEh6JXto0XeBvMrtY8AY/PLHwJo6mB9D9KMO
q1Fj0CI0Wj71mEGioYm4OWp02X5bKLgoOVvfe6FemPMXEJZ2s0tr8g5Mos0otM9U
4RjCkwi3+d9EVCunI2fDpWxVvGu0P7+TUHqmpNweYZNSWOJpHDa7AuEdvzh05HqY
Drv7CVKP6hW5WyW8EnclkoFi5JHQZTx6p+qzKbc3g++0bC9IRGXMMsx0Mo9ezIq+
lJv0zrwil6+lP1qWydb19buR51gFAcrORqQ1bn/qIzIRw0k5DvyFYvpOau0RHkmt
rh6JC+TXz/3J+gyXmMwgncShUX2UFGW2EzuPRaEoMQLkZc3AizbhWiroE1Uz4vVO
ryfEQUf8UeMKQ0MB4WvL71onGsPvutg/YzfS9y2KTk155mtcJ7BGf3Rtu81Qd3UR
Fiwuhz9j0rTtHM3L+7okhgGqxy0HmJiHWlYBRERNr7CauLfpCUBanf43ohzDk8KX
3FqyTg0ZBnvv4qnBpFnwAQizCZBT6pA3PLMcw3W0F+X9CUaoPqPSp+LMWCGktOCO
oL886UngrITkdeFc38V8uKuwbzBtJ5IwE1Nx1CvgDsbLJEv8kTZBiBex/A1HEKsf
OCJv5wGLZ5fK4rDBwKSbGRdiTqdPtTQiHj4E8wzvEFLGW5cqclpOBwu99fr9Sv8M
+tcg3yKbP/ssvymDsgT0MEvIJ/PfD1SNpGRLJkniGUiTm4b5MYX4Sqt58n/fxxP0
GED4CpLjiD+prbIWpekbixdVDjGmOf6i9ZUUtx9LSwaY3BOGZVUSYTU6mDAoAgb6
BgQp0gahzHk1v8h00arYXmimZ5phNg8i9Rdq/5+jI81xAyZjd/zTMELWwTdEPGP1
aotLLf4X3cpdxDvKo64tyy8lW2SyWU1LyNsv5N16X4/Xhh3ktgmcYppJsZmXFeQB
6fUYQ3QzoLf3Ln5RwGqrAuVvxTR2CGSWY6OoPEVs04agKH81urTGbLqTXkQPtzCy
HX/iaxXKn14hakIC/S0UkGgbdLQ/wG1MscRo+z41p4sR/n6mnvINy9HKUX41d6QJ
ULEdcZfD3wpYhGP0dAvKway9QrXUfQEI85HWRo0RwrZOLlI6/fn+2HnERXasTWe+
b576oV3iGrijfoeQG+BPKl1n7/WEuy1WHnwnA+SHtGVKHxM9iDCr2y56HYnxn4Ao
2t2Lz5lH2g/zmVEPobYGHXw0fQk6ebLNFuFlCLf2PE1Y51MY78Czn25ZzHi2VbkP
rLtI4jPrtCbIndMK+CzG0uA90DBH0otwdZCdGOt1/cpOAnf0pAeeeAfA8ptrhZLR
SSaiM8b9ukkiEIvO+3d9zVDiZ1TdBjU5WIHpWTL/dR3LUCKAv7ElbZ5TQijj3wSb
W2Ivd85KEPG0m8qEicyWLikOeGuuH56g+VnjRcUN8jAXd5uQc/hxiNK2hheO0CMt
XOvFWxJb8SughzAzYpJ/DKconp3bo2bFjSThefuIxmcqLT9Nui5P0HrWDppT24Zx
K532IVRDZRwtEApPOHJYn9Cn68CjEUbreLqAFu4ondDw94m9o4GFtv8zs0zDocLt
p1QOVlFFTLwABjZ9nWAVxhp9ibRuA4l2DImYt5GN0P4Ril0/h2y2GZ+1U22qA0Jx
4F3trVWIdViiHMMG9IXRe9Aw9l3E3gqLI1M62lBe9XRDQkuzhvFvcWYf+j+Pjscc
+7IKYF5ARixS4M9wKPvG03hQ1CaFcuayM6i8kr+3VTeaXexpfLi1iZUK6DrleI3U
E5/l17NX3W9agikbmZi3vEOgQcRV6xNzSvmUVmV3mMkogcKJHYQ2mw+XB1QEmUk+
670rwoqVNM00r2uQu5H4rb2dXlcnNVERv1LVM7lEdycRMAGRETyQAP/4SJs3e8Qn
G9VzUkgEIbXey1ambPlIym81fo85lBdPd1c2hZZ1DcNlbIfPR8M6ID2ilsczpvEi
W9OHIuq4uX4Ymv/xa+4BzGal+6rqgWfQl4WeV6DSda9dAlBwED+C6AkwSFGAy3WU
q/2poKxpCgGm/wmwgQyiIavhJrZ7PQODlO/ZKlOOQJ0LjVIIowKlbRClC+Airz+g
IfetsNtdZIoZ8XY2+/ZJwmTh1tEmyDtBHud232yENaPrYPFgOVITB64R9W60K0Al
4bdpXU3RAgsUhcllMFfiD7MN3a83g66Wt8JBTVjXOMjikLYPZYFLFI1YAg8eI2jU
Fpviz5+ivT0vIhl3QImJ0N31kvNulJ0RvHIPAMHefxjs7jOK1a3gX1iczi4BYeXy
rOdnUHqQ03CJyzMRtEuuXq7DWGQxJ4RKSuGR+9G7VYU755a/i/JdnhttdgMRGd4G
vHcfmhhB8nvrCYYfmOzW7TJ3S+D7+u251CXNGfGuBOZSA7lqYVITVsTF8tCruos3
hu+KqOZuFWEnncW5m6OoRSVlqakKfadM1kAqedfNY8CX0n9oS6EXrtwwBphyZNQV
fak1LGEZTFD/6VLRqpeTEqZUB+KxdSDBpqBgHcLBXu/W1Og5ZsPu0PAD/rlwr3Cw
U2f5IzHCcg5VHpCh4fX8FA3Kac9mRy40lPESkWpdvtqNbb6g/Ak9uLQMGaK5j06t
YlpvEPnlsjXKkmO93nDH/xlsSn8bsS7gYA91GcI10TWxeFjUgTywWs9fUjoC1TkV
jDhkh/aFicgwwtUbW5tq6xw3UG87hppSVNgun6QO0zsLKHSgcKOA5PbyVLz9XKCx
RpWBLt2yhUV2pU4YTB5U5+UfHpoz+bKwg6WBFU6xYXN+Yf9xpo8CVmdEG2Lam7v7
rxO8tiqS1nA5FGm6WSq8b4Fw8BvFVsf/Ueftvm3i+hjbAnDnAum9yAWcn4yHPNqT
K+PqSNHbpzDXIAsmajOW3WWR6ZbBBSClX1fnRyDKxKeSecR7QaPFSUOK8VFmPIcs
AHRHB/TmidN3aHLPEE724yd6PYo6zxUCpaydKhASOs5dzorVEREmFxZNP2AVXpyF
mJprVdVVks5C3YZcGiAwz7SNHXX9DHFP8vrDz5nofBQUXkMTJ0j0vqCR3jhSW0RQ
UvD1uE7/yP2zLz8P5H++7JzrMuOwp0ACMrLJrd8+f++blbvIPOwI2Knmav+qC/JU
QUDJyIXhZgdFlJjEaVNhIH7oih4p0rOa8SZ4ZPVlJZd9qfHkqevf4mnQULNU2t1a
qzAVeILc131gGVl+1GYgfllL1gZQBOCeizz6w62oa403LSVvhiua1q9Rou3MGiWN
Tz3YNvFELaqzITfeLzq2dxz9mGovvMTccmdiNVFqtbpnx0PXYGQdkDUILGRP1+WC
BVbjUkogWul9bBk26OPxEWNA7gfsABg6uXR8CKELI18J7ptOJEI9ZaIGRuMjhiWL
SQc4YVVBIYZ2jfE+22Qe7BwidF41Mcn4AqqMeTRYI4+V9GFi8ja0rwhS97ZxjgIb
bi0nP+TCKnSo2CM7GZOikWNt3HoaLR/jlUJf8iZ2dCKKMRkSx5oK36wt1YlMehbZ
qlR56VNsy94s26MLTNAJ33NxcBN7NNIMGL5YFKGTEPaSkKBrYHzb/jlnqGc/c+Bw
sIibxR0wHAn1Nfk1uBYGJMBI79xuEM8gCBXW1IPw10kjx7VpIJ9dVyDmP76q9tp/
lK0UagRbcwE77Kld0FewhRzBem7qqis2Gom1Kv3k4KMVrFfII/XTOKjaARfPd5NC
Uulxr2I/1zd9pPiaW9lFTGF/PHaN7bQ8p7Z173+3MBjp1hxkosnCQHUUzduQTjHL
43O8Me87D5jzIK/w7GKLL9Xkid2Mo+d7KAGDspC39ostKoFzvBEU3MzoB7vTwnTf
U/uigLE/Xs62WrYyzNLQH/IfMN1qouD4K3ni+3aGOpAatXgABQLGXN/JTJOGL0wR
wengKIxw9su4P+JMoM99S6zenHbtlF8MJ8Q2pRENEoeLAjyjgj5qNu61YQmeCJP+
676nqdPjC/OvoSZ1ShlYjvH6wxv4MzpTeADPfPBwh4prRc++Uc78L35A970veMO+
oVbIWscSq1kDncCReKgvnVU/7j1ejZMPw7OIYBuDgh/07EHm/xXjq5ttBSxKYANu
3uB/EYqOScwpmpYp2q/PjUwZQFrRsYAmd6fN87+PZmYonmRXE2zKeuyxU6DV2hNz
rxreWQfy0euMp8h4lJKcB5IBjjt5dvgxVrin81fuX0TKoHTJZhXNqi/LLwL1yyLy
oFWe6qG3z3osmVcBTVt0TapkkOTju3558dubLzpOnYUWNGOfovc0Q6eyugr2ktNe
ePeCUT9rVLHwyYhq02s6rh4OhjZFLfp/zycq/aRbOHOBlsQ04cY+ZE89BR/DVS5R
Gc5j6WZrKBj4o+Lejn3AfFT+HfagSFXWtccibvCM7WchGVKvo2NbCQZ6+8suC6i8
+IAf8WOTqHRn14DSvg2eEFovYqUpmIZpHEWFBbgceC4qsWTfELd64WgsbTpZ4owO
GDVOCaKRa2/tsqdZp2zDsWjTNUt33J6lhPq1v2dbAnr7WQ/eq6mpME9MnE81P8zs
KgsCfIeWXqa8CrjkKHkWaCEkjUWJDaJ0x01WfD33ZO6tWRrIt68jgsSBERMxhz2S
X/dYBz4XqwtySqtHMuyHxTj6pMnv4oZivK1fE7DRnBZJ7cR7KR6UtUJKd/qL61uQ
bFSptBl5pp2w8oZj8bXdIdHhLwLeRH0biM05hirnLuHxTvmjsDkqmbAJAkJYPcMl
m4bWi597wfjbyU+FW45lBpTfdv1yBxuGJkgps5tIsnQu6ckeUjpsLioiUvy0prko
gw+mvUfZPFnS28sEbyrGSvHjwoB4N4RLLIbD1Mp/boP3x4tZdV1NtQZ+l4YqafKe
Rbq6x78N6GcZ+7yB56jQ/gTZyvg0LUJLkOh6eEZhojbdlvpGs/qAJewiknbJzQxV
+REumkUfKVJcbUEPE5bOEA7MBHu9RG0zaH0WG7toQI3hHVki/C1wUkX67lk8Dfjw
3AID2HRmNbnzBUoiU2zeUWtXJ43CMkoxbFnaAFbfDMkIO+4zcEot/GBVtQ5ekstp
z5ov3kNbRCSev4Uzl//3CfwxX9adGts3QhAkBhGdbS1BlrzJUOL4cB4OysrJbNYe
dgtAvDm9CaHRr5FEJyXEopMFJCDw3xAe9VNwz46oCuszGP/tMp1FsXyCICMEdJIX
daTot13rJlou72ocOD3zCf80pnSvvuNwDds7xCSE05b8VaaQTy9b18eBA6AHHMbA
v4DUcz/0KKDi4D/tfrcMnXG2wKazbTjSZBQXRIIyZA/ah4A0pzZnPfpTXEPek5q8
04122N2vNVT8hCQc/rucjImF7t4m5wgIaMVX8C2kW+0H7wOwt4Plhn4hJD2aHOaE
OxGn8oKkOhwT9l0YLTvBgJPBtIXsWuCJr/btZUF84oeK9KemgErrp1/Qioedl2Ze
krPMJrgl7lnzxl9l3f0iPPXBF2Nkl6FjhZsquH75yG0CH4VV1cPysl7K8zvCNhmI
Pig8vHTMFRI5SadmBWhadU0XmctjJ4XHID1pbczEYqOH9Kuok6ppmhQ9pEdz3sSA
QbNsJU8zgxXXjfvzHfaADXu6eQeYm7ruXLPyy450/Y4x8udGJfYBPd2Ve8FYo66s
eZmFZDOzHf8KLQHbj0aVQ2QB6xmQssIxB4vPV26pxHz6hLm1XBvf2jvrRDzl9Bim
F4aB8akMcmwgqBShZTBaDDiw73vVwIMvLfzqQG7XmKcg4njs4k967B4AR5O9Fu13
ic2eKx4fVa+D+mmGZUxkc+JNRFnIK+9Egu7ci1AeP1f1VVBWb/24BpDoisxzdljJ
S96tyURreCEa5t3Xr+ZqFGbrC/g64tFHkyrhbPq+3oLmHb5jqQXLYgrfAqJztaUq
k1dH2uaNhDyqK8xG9YeRFj+OrsdDfni99HQp3LG3ClLOzrP68pnaLGZ7T/aylGkd
TG1Vb7onG1hVBPnibZUoQ5UFmDmhN0k/VtMalyJB4MKNOI4xS6ifGu3A53aJ7DSp
cefEkkQXZw6ubcd3MEvOSiGVlzxiLIUKrpLKZecgG2vMhOzWDI/VE3sfr0n8W+r6
B2M9SfBT1f82AgxVbRpMP/JAmTzLOleWie94Omy432J+kH+UjHRaboWuEc2aH9FJ
0jWlGtp8wCKN2iDPGtEOIApo5uXBmoZe+kQLzbQK9jDKKRHox+sdzeKbmOvwD9dv
t+KPJHGUWPv5s9iXMFAyhgPTVEEQFepk6jFKwWktiZ5NMYMd5dOEPGFnxUIHYSq7
ObG9WjN6I4IW62wv3Dy9ukDdpIxd/hzikTMQarn6s9eMy5WwaaRf5MW/z2T2nxrU
uXnafI+LwmeM4a35cGKi6AlHvCs3VLcRGFqCv5pOXX1S298TL6d6WGGaZUQFYLmS
GihoP7lJe6HS6TPGZ+Z82PuCn8izTNphuZ5nTaE3YYihGufQONr2EnjIKct+VgKl
wl1gZfrIvpfIaV3fSOklV/QHky7ktJCyfzP3V11qGJIT68dVa6iGFIdNc/TPNc6p
1HmBTuoyKjtk2XsZONx8548HY8ZbN99PfQvNkOBiwdXfTJXd+f+C3MMP2H/k6Seh
fdKsbALWgTkY+IERmiXpZkx6xsVVVZvRSv7t+kHXMrvnfLP8o6zZquGQEJ5Ox1al
CPygD3GgN+ppixFoxMFZz5f/6Icw/5oMV1C85L4zNuNNAGNratZxehAK4jRxS54l
Ot8aejbhHy11Og9hYRritH0bkqVGmOAcahVyrLs8Marz4Twkr49DhYFexuO7l9AM
Qr10Eu3J+JmmcF1KART/ELjCgr+N5+u3q0Omjo87gxDVVTEK/Q+ANN6GaXIDBM1I
bH3m0ztweGt9I/jngbcUQuZJRzElthurdcAbTH+lm/eLL44SqyhcyCzS7scgwrML
Qu8UPMw78g2xECs/9zVp4tDJPvC7nEkpBgT8kur00P7qWX3y6cbDATJsQsRjiErh
6QyxcmNHWcGLVkvCq39NIyzatbrWnhyE3hmnZgxT3CY9w+zv6HNVFsEIhOuwdG2U
tLTwpcum1FISbxenRd1QUMbygbCiotq0gNTVsUkJpMOQyu424VRfGfyQxEXCggmd
pHNZcrnRbKF76Dl8dDMgvE9eTwcbRW2YcjzhuRNnqmYq/eH9BRMOQ1OTDih6jDvZ
NV003cC2DTB035pQOdsyyg==
`pragma protect end_protected
