`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
i4ER9jw9M4xNyznXk+ZqMuwbp+fYcVYsCwIFWoJ4l8xwPP9VyWcKXy/nk8teBhZI
6rMD8RliAQDmbXUuJI6WHG8gnW389IZ+WhuhbWbZrlqTe3jMefWQq+tJonXOIMO0
hXtiEEVh+PuCKFwZcIyeQOpnMlhw/EwGq7JnmkxILUE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32048)
69VlOmPql/TxbueoIyRcDcwjbl6o7hsFyveDdiADTUfrn1pe5j3CupfYROCm4iG5
rwDQbWphdkLQszvWbBrkVivLPmUinq9haIORhK1aSd8e9iKQRU2Ll5DcehodKgCy
CCKfUoNy43IvAiW2njNNYmLTHgTbzKzCBWvTfb8BckqghuvmE4QMYMv+72l91g92
yYxSK+9QgyZoTS3wQrzdKCZdpk/2rcEq9LyyJLUKM5ej0s3vdUMhWNtZ4YXu/j6x
MJlDmHNvVjPCyHPDOmacpt0E1XA6ts35B643EWKGo0zmiuGTHFX99o/hTA57VyH5
4zb70IjcZlTycrJczXqmn6rOwKyzqPXOuHk1oztrd8jvazeIZSsTcZbs23HDg/t4
VFjOHLzWC3FxqsU1X+7DFiZ9xXBfveItUGLjinUz4jG+Uu4YxHRHzQleck7zA9sO
NvWMbvMdf2rscELNHkRV0q6XedULTaWtd/h10XOuvZjYQllmIp7cdYNCyMtEBz+H
tjIxfWQokeDl7WtbKfUseX207MiO+ULm/pXnHnSYCCW/D7hsYywoHRStOx5YBEsj
tTsWbyFs1KFzjzOanbje84JibVvzLrWgxmKFnRoQXensNlBXanKl3n3T6afpYyLv
Zw5FeJE/fvim/t9DZD9AmGV23cP+iOvDwxKDexm9hlvgLW20PZpNHTZcpPTyNy7W
GhWfvfsZPkLK8rAGMa76djqtgr/9zsybzjc1Zt2lqUYAMHqevHFCe9iLqoZdfMl8
g8EqDxfsmW/UsrOv0Rx40FHkmoGpJ7aLW2SZQqeqfwHyU41IoljWT78EJFUHJaYu
/7I4lzR1IGQ0fqldRX5zsx5gzl5r5XgDKT6/6ENt+NqfNVP7XgTZvNMLpW/OauOb
a1ffYhlk0UgRLrF1bxPfWGw5OGHXX9aAYavWlbUKnNzq54VrKukA6pl531KdExxk
U0oPTAxKNcIwGx8TLvfUxcC0ntCg6R0SAI68p23ASAN/iMH10qm+PytWD6d0mlP9
14V5+kT2KSTGfWqZ0/vGpllzsb41iMcdPDOxFhh2nKMSJ173QmPjgQtvINiDMPPv
LKDzts7HpgmPkJPXL3Qc8f/MWKlgT/J6D6uC8u5eSc5qTeg+D06aIR85SzrZCm+T
E8KzjTqYTFsuVUnLeP0pYkUtVAYjDUyx+IOkv3wDhGn/NkOG5shMDQCMvXHNMYyn
I1m1FNcPtO9ubkxzL6sXI0ZXi2FjmErrr1NncluBdYym1PTmGoiq5XbmZBxX5zm0
1abj1fdH/UHzLaq/lGgJJgGA1tNAucViXZ+RpZOD5gfmqSo4v0SK/IVX5ikkWMFw
OdzagcC0CalHPmPLHYfSztEQdGKrsc8MSHPhDIu+YeQrDAmSdIRCTs0x2d+yqRmo
SZTW0u6mUM+h1ZE+/LyTwKG++8HLwkKJdhpuYCG/+BKqyT92sRmb3ahIoxXjqYi3
4ec9WdouazrUEkyEibL4QzugySa83vdmBTfF9FIxkAEBrzxx9l2jocQ3hlf9qOjS
5WmlXJMhHwz1L5HhdPW9zMHUjsDp2UEeaePn/v8S040fwM4jdLOG44pHCkEtFpQe
eTLrUccoRNO9YYZ+s4PrEVX9NSeGynBS7/zQkSeNIvRv76bentEK4WdIENsKjeKa
urxj6adGcNe+OeeSFbXfxyfBO8fcgY34w3RFeGKW+JaeeC67DjPlvM4JRgsI33AX
rXZjri8tracIzVchDTO4CseNjHwCeQa8IdsTbgcd+lrJ8zjJRWAtebLd+DUMlMI8
eo4Sc3dVzLR4A0LGJ/V/eDLy5rZ0rZVePQ97A4zRzJGiz4biEp+pxVztsdVJVS3r
nSYtUKs8lJSvGWJNBnkrUHauu6Fl2iKXMU0fZMhH44cdmNq8qnAqBtpZL71t+pjr
ar3RcpYLIQojp3hpVC+7KzKHyVBnMjpTSABjOQcSlPi9SON0ODa/zbPcKQhVgqyv
H4qyBeLAtJI1R6emb+1RBZZW3fas2LBWzb4iqyrp6d1SfDjL0p3IQ8hmbrmInBJ5
CuZrtSd+CP/cE01oQeC2eqYD7kXR2XOSOdxna17eaaoFbJCieE0p0oZn3IvjUK86
E5o4oVbXG5crxqMlRWbHYOyIBlUm/ON1EbGjav9CM1eWGvAX2M7r8iNWQcRRbkmA
KtVUKU5PuXgbWp1GMei3IbpPnvYlmMg0Uyxicxz06hr5stB5TnYxNSMsaDWRIxaT
lvKPKCqB4cNWdtMBzUljKLGLNcE4Bq60mwPPIC2e3EDDtU3mfiDx1sAis7eaeu3x
WofFNLwoRtmShlRSwNQNE2/+cn/lJqLzsBE/g1GbqxAswxsKi1GpiuXCozK9eHaY
8er7g/mZ3YbjxRBDBy5xl513pp7PBmNV+WO+sSrhLtlEBDTh0DDa5rRFwM+FjUdE
tjR2Zz8fOiX2metP30m2QLNFcBEUkbZxkmlMbF0So9kP2fsFjMpppsYBDVtRaYn7
NvxTUa0N6BzYsA9rhIKdGnX55u9KDmn1U8TRo2obtgdSoHviQmkK8d5EyhWUU3C3
C43VO2hO5Q8cWtbVdw84injGljOqLf2P081crgD1WNF7WOQN+pxKkTj8MZqr7xKf
fbJmjkTnb8+qeioF+JfCTYMqowE7weciW1bHww0HZHi6w37WpUGAkUcMqY8dcOnK
1BoRd95X/CeKJyKserMbuByw1fd/BfViWeiBa4fH5JbWCiQl5ZlfKUVjRpU3uXMu
sD41DuB8sBwdAvwfYPSOdAtjsyJTpT2tvZjomv/ODTDWDfTHO4kK15BIKVKvyqeD
HbXzWLDWG+8ctfK51n3xiZ+pwywoax8QutdEv1jmfTOhJ/QWB2PUJmGsCcJt1g+N
9ptNG6LgYPH8v6pSLLYXCWtfQzvW3P4jaqMWpWfToKS3ays9YkjsLOHGL+LrZhFX
x2p81qw3fuMVBxYZi29c3WgMdNBI/9WSW9iHwTwexvs4m3jQBhTDtccm/bRJgcZo
cUEKtJy1m0p0yTpzLRBEOfQN9wkD0/iof+kV5edN9cwyyG43hrw4pRZoW19RprwE
ziqaEUGyqPFTT9z4lau829TgtJdYq2PdsgvTlan3ODf0fFbvNiUhfncFbp2okyi7
6+5fQItvA6k3GH6SuYJL2dnG3PoZqdtkyPPIp56fxq6QUMMJdC/yc+CIIJUhIxGE
twvqavLqU2u5mtv1fftwIYLGc82O8sUN9259FU7lYh/adN+oDCDjFetSLi4JA1Co
0UweauQXU6/PCjep4ypwdr7fOzzSO27IpzAF3ieGogWlaoXUbl/RbVlD96PSi2fz
7CMAcztWRLpmEj+4MhMV1MvVCUOR6Ap6AN8JKlH58dk8FZ4XNrKSOBsHfyokAOww
k3yAB50Aa0SZ5cimJpQDG8mM+EGYxG4GRQFovrXc92DAsHOjS2LeYullentcIdof
ynofi4ymvweTi1OEUW2Tbs0CwndctR9yKTE6DRdmVEaRhuJsx10L89zoDJntZgro
dsvpEJrxcBucz/KcV8DYCL6TcvuPncA00yQZ0vDkI5G6jWrieOVu/52/MbPW+48U
ygu0Le5WZ6GoUU4J2SLn0nwCbqzLe+yDH2URWNETeAth17SWRHiNXXO/mJHxaN/3
oZPzUxQDC/YWLzNCPZDkJa1B9kW1gV/ugg5vIkjynhAOJF6s3kIu2GhCmizUsK5s
E7e9fFADjM/leFydxPFM3Qh8+tsoFltr38Chvk/lryhIVV0xues14+kFnntjbWtt
of8JXASM/G+eoFaUMrznAPyKHGaU8KfyIZmEFZetdv44Jz6jW48osu25D/ERZs6K
AVFxz2yNe4ZnZ//smEn8f56qnNnSEXQtfjFXL9yXbM49sKDxeYajm+94ziPPoPZb
4oPjb/yugpDs64lWMjgsVw8bL54KixISMVMrKTS5WdZQle1BGgpkFHf2lPCsRBhu
DR21ljDfIItQ5qn6uiT3YuCE1rj1QJGVdSSTkwP0sJ5OGepg9ygo4Dqt8Jg1IS11
URDn7cbvn3UPlr6eAE/roJFkTn4NfmDLrZ2jRsgNeJErb9QHFS2IClC50Hqrfi2U
QfSRocRl1fM3PydU+vfC/rbhWEFirAHZm1N+N3zDAo+hbFXy1kziPIKuSXUCIaaq
zZPiTGh6vd8XDNso5nwe3Dhy+4o9jWTzkTFYYldHcLdVVaVdCovmZ07oMA/9zfJk
B0p/1bA3NGvTu1MzRWLXf3uExRnUNf53j+zx5KL4gPCUbZtWMSygo/BTTM8Iu+gO
f/21ZgcAOhQ5iOHx7iw/23jRh5klQiKN+7rgbh/WSWX/xnU0FI9HYgWBbyghzo8m
JSln6erD5ZyyoGIKk6mv8ohPhTA7SU5RRGZJoO5t9eVueuSMpQH3UC2b4lXUH8P6
AcpW9pJtcZ5Np+ZX5t2N87cVMNKLesvJuwdFL4cK+GW7+TlAMM6D9BWTntdUsL2p
dyum4abCnsclO0xe9GNR7YsTAh0d2/Ih8ucjU7zU+gRASDsS9Cl530gwaqo4h+fX
nSwznTuaMk5ceBWGR4sjJ67/3VJ37XiX8BEUK38g74DmEw2n/QXjGghcx+xgt127
EnXtI+R24qMU3UwkZLMmJP6fkLOq0JIUFgbLnTolhYcFdaYAct3tlmHPW0EBiize
4b4uUnlDC235JbTX60Mx+9x5wsbn+bTboO/uZWAuVukaR+CPPLK0Fn9+vgjL73cA
eMhvGvdR8Hsmi8cAJaS6Ispyn2ompxbUppKlGGjMC3AHGaudhVqpfdpr7vkZo/RO
P4t7Cr6c4UXbVKHVd7yzg2vxuV0z6lHWqDVvPtKJtjC1A71fBgmYO6MO0C21aUvi
5Tkmd4e1AIsD7hnz/DSBQluu7Iof2/hKGlX/rBw0tb29FasACcujZPLFuZ1BZhI6
wdWRYn1HVQE4Ee7dg7cU0z7IxZzTldZyxkU+rC4Wr62y2RaTnCXIVJH2E4tL4CGr
ItTEjuB0y9GIXEdrNds1PR8dT4s6Zp7P18F3HPY+0yLduF59UA4U/nWQHFO7itnD
DzUNlsTOh15uj7KJRdNTifrj8gfaaifUgxuXpieODKEFA40iklUlE8ctIav60GS2
72s0pAqV8AB+rqnJP/a/OdHxKif+0qVaZccPNeambyIyH9CjCvICAmD+MiF2Z3CJ
nFzSXrCh7yUbPiwXWq0XtEY3N0ZZRYPhYjY8i5n6bfcBXg/9NI0nWyi7uT+Dj6xb
4UNEsuPGoc0yTwR6ednnbZa4BhVtAJcmXaxG1WXMO8Nni2yv62QUtlhWX0rZ/VHT
/eIJ0BiryIuxvh5bJiMsZmkCfnCrv/AWtmHNQnlOEcZy187+jjobEf2S7Jaccf93
kF5BuWCZHeb7Vh6ZevrGhR76jiRyX445pYNsZ3cO8JCuo9vNMvSj8mcBULOHWRdF
mLnJ3koHV9vb2RN5fM3KmOcprmEdzvDJRu6WykA46fMK5OE34YHOx8s6FNMtCk2/
AaLsTwxcAk2Mgo5cX7ZGg1izzfc5rAIzS32NZ98b3vxKt9OoC5k2No+porlHNvKS
lTlp8g6cq+Tddm4eUr/QRI+joTyz2KoktguFzuu0d4xNF+tZ7jEdrLGUMZTZd8+l
rZCXaSX4YLSRm2yNfblSEjBLzjqkvK555Qy8lFrvZZ7FMrj9SapvwYHxkdMh66Jg
pIKt74hCvO7cvqC594UPrYLTNderUxGudiJiE7WtAdNMzgmQnJKnwu9EvEXMIW1w
d4jS6y6m9XkXQ7nM69T6BRwNQPMUsa9rUc4sN0TS1D16CIyRXOH3lMl5RasqTzY0
kkUTiS2epEXzhEEa1GlRrAJ2nLqYdzqiDtx6uS2ywTiFZhGt2mZWew3no7h3D+Ho
dc1+RZkbumt3pSnP9A9wDIVD0fe/+xJTFxIKaOimAVihwW5r6PJ4zQ7FsQh1kRMb
bQL4KGDFqce4rZ/mI/XQT/3c96sA/R7YOtDRCc8w1QAFk2qrkJSjjYMmVCWr9Bj3
SaX8Hp+xL5YfhiI/ey3nafJu/fIV0DeC8QolJib9YP+yDi73d1UA6QTl814Jsz/3
LAEJuCH/xbxvDQJDccAHuuCCGQUJWa4U4V5nsl4lZjnXoOpqd45z6bDcIGUTo5xO
fv39uOtykwztMcMb7Hpu1hXNfBJ64AQEBEF7iEYbXfb9nXDZZpmfqFdS50ABKrVH
VIoUAv1FkOyHH37NWiBimdDcqLJRZZBFilzaow3xyYIf1ZcFl+R0iMZQbuUlibOO
6Q5IdtdOSFf95akwrV2M1LSoif2095IKJOwQEnnnwQJVm5CCy9ZMLzrAy58jTRkz
/dt6susUgu7yi+p1BQvLE9lY+AopwNU94gGRgvOwEuNxsLunJmums/lR5umOU22v
4C/f/nidwicCz6zfQ6G8zRMyz7rtUFXTEK6I12pWdC2PUZ3YKx0QMp6tx3Vaxmja
+meTF+LRZfvyaIlmWfXReqL4g1EwQBK0ROFxBb4krapvxbXxxGpTzHdaZuwDjX0l
uk+wZt+gUc85iVMzrQzjJNRqRTWO48AL/6IKJU6Jnh4qTqnCO5cY22SxoqL9OKk9
AGIy3Jyh/vkuIiWtQ7w++sd+EaGoI+s4LnD8UvtWTqvBu0bYMbtYM/bhxXcCKjbg
F2lTvPxD/vOk+s2OyOhdYDFx7tpVGHRIfnlVMN3UVutVBvgVbnlVB1Sk1Pn6kK4v
ufGHCIl9e3waXiiBznGEw6+9hkjvPR0qK+Cca5tGOyIs+3Xfo0f4GxdaW92lbQyK
nmcSPJh5J0no2Mzh7GXl3gWtZtBaJ3xCtpyaFr4U6+9fKuKbfIfdN1y9O5vrVqjU
nH65wDq3A/GEffyIFqwKZ7xtNrsqs6NK/IjUZWCuR+Cggfhd6Wv1rK8OBSZLTwOD
t/axADHXLm1BMB9S6QdR+1fKzxIHogpwvvzJ5PUlkGDFk0ALDnB/MDwsOVHZADT7
F/F9JusZS83nKyJJW9sTJ8MV2E5h1Or10DsFVbS5XjtcgTS5S4LXmC/RtunRIU0q
ZTNyCtlLXqBObCgE33wK1Rq0mAJHny6bZ8++2oUalFhbPyyn6NXGicR7uEw5l9a+
0n7pZyWpq0ur5lVvR/HzU5/FX1tY8aEr9R40qRiRXG33Fz2KvCwTvqdQJ6mooD7i
h7lgvrB71FcD8CEE+XSkjor2kZvr+qNt/LwfFTICDupVO95Xayvi635sVxLRpkkB
kTsEb2zVGy/m+7+rg8ghvvMJ1EYEk8gITGh3fJXxegh1jd1DizVU6UxbXz6p5Wuh
y8Ce4qVWEabSchKnVf4srH+GyZ3VsoubdfoYp/ndtEcN7RTPq3TGzUuIfF8xkS9J
pd2uZchkTZ7UUBvHLm8xepyOzruHSrPMBv79f+jlQ4HmJCDuFUUeqmj8brBu8b4n
2yRG6p9yx84T4aLzcRgeQW0Zu63CP2/A/GGCqs2hI7rggP8jMvVcLo045lmJVA9j
I+PPEAXyPvgkSZBcsOQtQ7+DNiTdasc5609ChqD4iziyf4p/PWj4HSQua1ID/A9/
g8kL5PydgTGAivjlS/40sIo/3OL/BCyDG0NJcyWvWQOvOXscfSreD+6iffidbQWK
G7urckPzcEhkq9x939RZMmK0qAyEIWFBC6ka+DaIrORXke/D3bd4V0+qZiH1/EU8
DLdVTvDnR00QR2wn3q8SecBfU2iLK3m5VQFbxxR4xNsovxJFJwka3XPjt/3iC8HH
65FoyWQRv3sc6Y6v6Hr4D046xjcSXeJtfAiyG1i3/TVNkVhvQHSloRD0eQIe2cqW
IolW6+8HA4lkQTxn2fdkpG3XVGsnBncIEA4CJroFcMxIiJhM/94z10tAsAk05xOr
kM6Wr/bQz/8Xh2KoWRnz83MqDSlDiYPH4TkmlA1xt8yVTff8q8yIl22QxvYOWErz
5GCaJAETqz/Q87BFATBVLm4A+zsBvwuyn7+dBGwjhcbY4Wx08iSHkc5rA9juTzRT
ITEwPLmVWlcqo5ipA/x9HJb7WWnTTCTiQ7/cogutSRgIlyWDT0knus6gLqR10wtM
VZXgUWK3G1/7l8CTFa8r5aqSr0VBcSmLvCCVXM2GNG/sk2VU+yvWQM0hGiR851s2
t+GOqN8xvam/AgVKgMh5+SIdlV6yWKCFhejFsIIP2rD3CWJ1uDl0zapu4nBSeHZ1
BThbtYi9Qex63Tx8oUPw/Hn+Rxan9elVvUIzHe8ufZVXmzXNjDY0eqUFqD+6GINz
QHT6/1iuzby/ALdQdx4NZ4Wyh9dGi1CDtnMPLDwJnOsSY2UHo8A0uLBYYiPYthWj
JWjLPXWe3iUW4CHmFNp27kHknW5Vup0WNp9wZqQOKHzzviNO21jGD7JgPgxmfAHd
Vqxtb1sAih3W/aLQttoYP2Vyf67tyzeDjpTCqMwQIFfTKTYTacfJMg+TtCxaOqG2
Sy0wMB9SYHFPUdYDss+y4o6LlFG0R5zU9cMsxnS61zRDfCsQ0RKf/QI2lYrO1h/O
Ea8NjYArSo0H9j2O6MeoyVhMNiXhxtytZY19pGyW27g3CNv1CpfG/RiOaZ7Aj/u7
wjJR08jcagcbhb5FO7jlwm33AuPhj/XeKem3LK7cAkv7tLDWEv2qpIMDAUD8DXyd
bPW5MDxLL8ftBsM+rq7NcoW4ScjtS5dA6zP2Py2l07Yht4zwQbkF72Cd648tn7bg
uFEtsEF5DkyNROnbG0K9xcpTMq3yLirn7pQjuMEAtEjwA3pRzucqV5uiZty64d0E
C0x80kWUUmNsZk6WRrDn53l9wBds/jDHgRF1H+yo5hx9muAOM3YFrWfWz/TMkKCq
psvtlXnoH4yj3oZxhpMujxCU8OrD1D4t+YufoMBPgUHRTIp7UffLz65jDLZ/DkkI
v/TUtVbav51oQ+LqLVv8+PL7ThA/MDx9J9hjpGA3vb/7EG4XmhJXzudpofNsdOnO
ydMwZYoc7y1g2SyiJ7KPAwNfQcXinBX3dgTdNOeEdNIgWSnzafGk0ZqMUoA/GTaa
uQdS1QoEvTMKAAebdoYyHeuMcn7ucu0luBxuKyf5XjYohlbCS+pYvXUdPK4iwQct
gDzE2Qzx33lgK6UP0VLIyuAlxEQu4jHGo2COFhQ7T6LicBidLCAxFjMNi+2FgAFy
aUEEW4Vs6qSe9hHhmESjVckpepbzwYzyKvBpj/L2Ebn7wvH+6X8ec0u6Mthw3JTt
rqL3tp+mMdwN9c79UDWpQv6P0n8kViPcqdjKjNLq21jgg9XOgNdM/AcO/64ItKNq
7oNrRet9xdhR5tFkickNu0UPvLjco+pgx/UDjFm9DvLRtNXBB/rSsRcX7DLXCqs2
4gDpgKgAUzpL/xPaa0w2mnaQq3qlh4fcIFrSzP9easHnT8CAQpbqZIyiUaXYIQUC
HkSMnpGBTNaH0y5DrRpnph09oeWjiYU2q1HGGvnPxAF14+ESQQjXExeR0KvYqAQs
e6pfv4Em/OhOb3nDRJiNFrc6B+02f8HakDjfN2iZEJnt8L8uYnnLVjv87whjJXLn
Z81ETABgGUjUd+YRrkB77BzjCQV34tkE2X8LDegGsyg60GFxYyzj3FlIoyTgF5Zr
vzpLDojewlx4iIwd9gp3JFnbZI0fRCN+nFPRhuyizl83AFSDIRoaaWXrFS2GQgJx
ASuvBZzETMovjEl8Iu8XeL0JrQGIGaV+r0nrwtLBDHd7fLEvrZ5+FjEQIgscZNF/
HK5LoWxaHgwjHQ296wpnbNKwXYdVCHhkrkwvNvfO9o12g16HwJgRY83ySCUef6QU
ifyK2Hk3eCaBJScV3hzvi97hxdL0ie1LMUdChm0gJgEgK8BUR9LkKmTWtkOZfmwM
e++8hCs/DpP7R981VCwlBeInosCbK3C/idrVXYYKAX0mdxZlC01AH6XDGP1Sw3mx
gO/2GyBRdMeBPq31E3lworFxW4vGqXuLbGfI3nEvhG7LtDmNDLdCEcjLZlRvf++i
TXrndkVI+ifUUSul4QjXWGC4iRU3d7UX4egcBgnjoCaWgFJQ5nTUp4+bk5WjazxW
nZomR0IqJL60bXFMh+vb9hOP3MkQIzeAa6XCaE8Wf9Mg8S18RHddIWfYWHMu1z3I
T4xuMXtpIu2mZnKgRSvfLp8hxqNq5qafHzCYSzuVFgQjeHs7HZMRnBFE++OE5qHL
MchRkkkNAWbViyhPk16o5DLMf3mkEEP4bdGgrzUuZGKJkVcOmCubiFTp2VeT3W4m
MGMfW9ePgw9oRqvGb5n/Xzn4TtI8Xpi0lEi0U2mBy+dTXk4tBF66fAirV/4/HiGo
LEhXHV+MgYJLqvupCkeazlo8v9eR89XfSigcsjXtRNhdOKay8ND/cPzx2aSJaA/7
y37WzosuH0i7zzus9fY1zoGGCfo2FQZPWFPhuQT6Dvsfz+X+/Iuz+hcbWDmwHKqo
69xw7p+SQTGOA/vOMSn3+RTe1QJYtiO/ID0KUEkN8/M4pFdqGxp+IlJ8yP0vx1IT
ulFeqvyZN7tc+k9fg1zEY+a0LrHZZGLwP36oQJ+0uud+uRmlZXTIlQzg+k0Bw7g3
HkohKLrFXDlAf8inol//jiqFIbNxidsF8FqTdqnPShKxM0N4XGEilafC8iddNERq
FUzR4X9O3pEmNAp5fR3V1GakI6We6tTHQHsu6b7Lw8t/JENvHDrcSqOf6qI8dtxb
8dN5k4Nn0ISa1NqTQKTieHKPGUSzBKXhNo3QfM/VPO9A7A5K78dBDXNt1xqMDqPI
DBfV1ENa8zX7gajL358DkYKhSB5fG8Dws8aWDeNYjrTjieZqZFZHO/ROmeGb9QsM
O20dNMtyMc8DleyZffHITczhMKjFzWaMtMeGLxIczfQHRJim+rFhCx3uwjUopHhP
R9UOeyeT2jxr+f9zXzV/M3CAetN1qV1rLXf3AEvODFM0AOkrmosSseC/0+o9xolH
NfcThQFcyfCbIwHVqqjRYtfCLZklXV2TfxEp9D83nFJkH1+y0XagvaoylUixFxCq
+zlEsK8r/w5w2DSCj7LTCNeCnwiEQLx/R9chMHl4+PHqLDOqszT8HxiOss9PnTyS
lHxlo3RWanmgO0djXduyufn1DumuibxzfrDw1XWwNdSuJ7V/XMokjWGdHiDl2M64
FLRoQ1MiPWz1QWigzrbAVwWwClIN+nmiCnFXmxysUL3OUlI2yrd/MiwACPcE1cUk
sIyBm6OJkyzwwu/UqNXohDM5aq6gDB6RG/oCsREhRFjXVXm5RFY03n2Yv0037QOk
dLQSWTSdJfYuLHTK9kQHMl9p6bMyFjlHyRuhpjerF6HJD+uEmjEuOy1FMiUhljSx
7Z0ibgsSvmLofpdcM84iUvA8jwgbZ5z2Fe3Wz6UPTM/Zjbpz+oelJqxI+3YSt/pv
lcgR4axRgjyjxP3RX4Nel1FfVkaclUAiRQOmi3+vUZZJgysWT6YutMdPJr9A4G+u
LuiUbGmDm/SaUKffB6Me3/sHJNUryVKsf3kDoxqgBHke1tEM5Kg8FR+UVonQ2txL
SRgI46adwINcK20cg0AvK+5e7RG2qQH+kZbRRLjhl/uSHClInpbmlUyax95MVQD/
eDt0m2abKailRzreUCAvbXIz++0qXDajNjc9CiAV3qHW7Upf1Y43hEx/gHseojjl
rAnFAP1DuMVOe/OVX8oY0COv2nJp4ECHdq+Gi6DiYHuEwWxXxoerrv3pRr3fHiR2
zQqaZG2lG0X7zPrCvBP/mGTzKsUICF/l7mH9bu8ECFrOmmfZL5dTqdXMLOi+wKE0
+P4xzqUAvH5XRWpYTl3xWDOF74f5qx+crkqoMyg0I/uqNPnRfeG/JrGExJXiPuyO
Y66xMRTnJBsIzWqmzKYADDKoCtveptLYxBzvEseQT1v9Z8hzyX7iA3DVIGKGA4nz
f1CtE895uvE5lNRtoOWbrBeL/akfhjRqwNsuv2rLm1VGRIkX/HT/ckPUi0bfwy6h
Hz7sXZ/I1bQfKcSzRv5MyKwFh0AX37wVdsD7xd8AdczlbHBW/kYpURAde/X1WKC3
jA4yKFYPJ/4A96GKGo98y1aHLCIgVKx3RiYhffIb0Oa4xWQr4LG5Lfib2DPbDZWl
h7CDt3NKAiNsFMVaakNRvRpR1c+YmL2F6MwXLMKGoUa41RZ/wOD2aYncYo21yqCD
Wp89DvJxVa0NAeI9apeDdnEDSqKE6gL8Pi5MWXE5/GumKcvx1IHoSnlMoQJy4BSI
Zpq8fc9vFSXTEvNKDmRXlP0gkshWCjVojcgKq53tAThkfmRUQK5v1RHNhEXc6ELK
NTQGG35C8xuh2CY7Qe8tX7Gi2BphB49MhSubJGFIuEPlZj1O+yaqD9XMOnkg+0as
BW6r7E+arKq1dUA6LpvKM/9zFbAFYLxHTqZrKcRTTfc8+vs3jG34FC5jcFSvBZrR
IUKeMP4L4CojT3FPQTnTwWjHNfGxKa46YaagVaIJ73/3GN4ZF4TXadeRn76vJBov
4k2JxmDFs55/uKmDCj/PHK9eLfzpSKx96ANVt7eyioO6if0DUtEOqnJCStiiPFPY
guY48L8GIDrqpUQfXfeswI2PxeOODuBzqiDUwbJYWUeUl0hGN/qg0Wkhm22MmUUB
JPqwC0d9o1m0F8w2TYWGJUY+vNgwY9Y30GEL72WExfgxDaaOAXyRHeC97Nx+hC1+
w7ub5KUFxYouLWHatKgrQKG5yrbw8hLxTIiGX4+t1wzKXh2c3PGXH9jFpkVIebek
jnHLV6D6JOHvKhVaKVp+96pwrZ6zBLZ4yfozD0fN/QSCzbtEH2sSlSrq4SCW4RlB
VOLpk4UNJWZFS6dTwv5IOVC7YfpftMU2ZVt1GFaNRVvF5D9wj4+TFTiZiIlIhEJq
6lBxtJHMCBSTNN4Cws/RI2pRi5SYNVekkHxdJdjRTKnAnGIFYfoefvbduYAO7RyT
I0euBykXHckIl+dq3HYMZ4d30aZZ4kAd1YAHt7WIoprXzKFRayuI6fQgJ7C2v8Qd
do+YuAXA6KqHPvl1vmknaQ8SWT8eyEcgjayjlLbWwdgg4d3rpaEkggNMNsrDVTZN
t/sxwFpa3BfQogNM8DqbtYaNNmw/alT9fFtEaHBhzOf8yXRNqUyJlHYJWwkjxnh9
W5zzspzFxUOKW3KWxne0EZ4lk0fCEGcc5hip5APrpEvVsFrlTuqvkYaqKc66SgH5
WMwCHHueaBacinKF49w5nOrAhUuOLNweo8DZp4PuQNHk8V5D5Qm7ZaGJ75xreb/H
f5+xHKEA4KXPhjn1QqppaZLDuPNdVYZOEbpZplTIwJ928S8gSwet6Z+p/FamY655
Q3phvDEuHGbiYUkF6+6aBmouK49sMHzo0mclg1ByG4nbHjv9pCQqIS0TIBj2igi5
ScVqpSg7iqvkhxdhB8ZACShL6E9ljwzYMctfNOcQUzQrYW56vEeJVw6myHc1Makc
+ZO+K6ZCwSGr3YSIMnHlZa9WkplLxZbJxKz/kHAsF8ueDydKRwccTndpwxpViw7g
P3OpFr3HyV9BuYEBxwwaJN/IiBlKjg07MoVbQMAVH3RxhugB8EFQj6QN5LAl0K4a
YW+E+66GlEN/6bbzI5+1pfnisCBeWRJ6YDAcS0tUc5wTikpY1ZMm4fNcQ2GBFU7I
yAQl2if0BZsZZ3LUjrJC2RgDYYV3f+qlJW3Z8eP/lKrZJJKcaGZ1ZA5uxrhvwH49
lizTK7yAA0shIyUUcLvlAga+s5YCsyB8mRlVppoIGYwGiM1NzkNEZE5HcOq5DI0a
5fivDOLQrX9lNDyVo1hwJCNUEUEkc4s7ICj9JUoZQbXbJxxm9SQMQ1FL/1cLxWVq
s2u0ceJxfWk82n3jqp0X/PIolQ4Fwp67iJf6J7ENtxH1+nrq/rymWVeY1pSV+1pJ
sAtguo/hZAX0+o4m/Vic2SR4zWQD02MyubiSou6F7L0nZA3MRCNUzEJRi34Z7YlX
ziK08TfL2U1Y4fCKckDW1ktuUQ4h6kkRgLBL0qcn+39frlMpMs7Bmctnv0liHKvG
NSfZ7hbrPgXH6rCERUkiJFJeIHx4m8IqzHeOWBz+BNd2ezsFvqBMfw7+1x59aNut
sednjaOVNROcnzckkRa0SdE7ugUBW290UsvgWaKY2tBXKYihVtZAtB8udKZ6KCHk
LhvpsAZPS73og2A73bqxmJXeSaUY8jltgnQIHfFvhTF+bIcNLlCXJSrWtfu9K+K7
9MyLILwUo9CXKf7R5i+Bo/XdXPAYAEQgJUHw/HU/kjky1H6KlipwqXEimyc8PFPW
6TGTIXvFfZ0nXd946bDKlD04hFMJFIXm2JkR0H2uChjoB1iOsHMv9Jv1xaxumg+T
I4jaRBcGJ4G3hFwR//7LTwvlJESKdQkQIn3UxlVM4KA2bL+nzuikhdg/Ha3fkaOQ
D0HvF+FLctO2f93GSaNqpcg/6zUBcYuFL/CIv26WWq94MiGNQUsZDuoe8GXJFJ+o
9NlJjSKOzADceRMOLCvZK59ZpWFqzgzlju0fg2xWsLE7T/VtWyubOr2Rcf95FlLT
Ndt0Za0ohrie8m5Mteox+iP2xjMaLXCWJGOuJ1yS3AvF82pDmFVyjWOtVA5bSRVM
D/XeIyWeLDniG7rjrYG7McB645+uzerjaBVrx6OoMX5eYYl4abvArheoqilEJSvB
KD7lgTAcAQgzhInFlbMRjkRskXBQqFCExf94V2UlgTdm4FJj8RP+I4QyXi7hk+86
RXRBYll9yeHBuzgS5A9JEYFVZoi/KNnfwKwE+Db226+7073v60DDFKqlrszgM4Qw
N6hL2L+BCAaVGNK9c0MrloPY4BNG4QrT1PBsXHGSYOdiLgQfku+DPtELfx6Fpys9
mgNDLMwhREqtYlqxS6Vyxe3JrZvkZzZPBZjEk6pjee3bOgWglhnt+JMPt/df/yPE
O1np4f1KUsYCKrVCvCMK7/aAd5zw34MUQ6efibmNQ17+5wHgb5XreRfg0ByS+snK
D0UaLZX3G7XBs92myRw4Sue0wB0USvGiHftaHRN6BQcJQ80/q6AeD496Z3RMDH1v
Kx/EOdm6x08xuia8z6wTyYeStg2vSCXguVHs4PFHZyoO6mDjinjDpSzywnFAThNW
SChESTTti18xmhIQpnZRLsg3wsMKg73ZOaDoszkECW/NSHmNcAmaAsI5aK6KckRr
+d7xjnOtOQZzHeLm9zNHFqLBlvwkEeQlUE1iA+3FXWyAbVx6qmThr01KoVMqckbt
X5b6FbWpnmqNA8HEwGaRC2zrLsI6N9WefWul/An2fa0BCibiUzuoXTlGAOqOlgjs
LqEDb6U+9y5WV29AUisaIhin1M3zxwBYWyN23vTiLbtXOS9y+ZbsNtla5g8woOPH
kPAVNHnww675JOz/AUie3fmtoWSwmtAbdQKKVoYRm5gtIZ6w1Pqw/37Lu8B+EQzB
DY2Wm55UoQm+ZQuzGCNDOwBtGM3Zi3BAjq5F9GcYfGn3wHw7+9kTmZhXalKbHiBm
F1989QyRUu68uWE4urMlLJ4unDowo1jiosuNCK4GmQ+fG6vXknCtu8dAmfP7qQ1i
upX9JKTGbtm59eU9qA2s1cFR025s6SsBUcUP/mO+rz0f/FKGEum7PtnmzquQYemf
BNKIkZRsBt6zpKW2bj4g+ePSd06sWEa12TOIVTA+Y0xTmwkGuvbOzYe6esbkmcET
d1a+TYsI1IbWDgHH9XqgUBG652c5ae9TPUddQHHPofqnEuKR48Xj3oUkQilQr9s/
l07+RfMZk1RN2zDsiPM/AuCNzbMUXjqXJpFLdF8IPV6z7R82Z47jTrNYrLuKJg1Y
6nciAdoB0DBMEwznGAkf9Q6uJGfmrh97dqBW2vYIIPSvxC4wMXkE2F5ztx5J/xsF
DhyaCxpcJdSWChs6yeanMJUa+MLGRSCmn7OxMB452gGUIIFdJLj/oMDMUwnpX5+F
Kv6HKj/6jo+71B4n/T3r8jBzf6aUZCsEDq+mqtzpL5ifZ/TpbYQfFpBaOg4G4nmh
+YngpZ49CtlRkW+ANfE5c/Nzmqhgc/EiaVJlEZArrYeH1NNJdwiK1b25qtRXy5OK
sktVdbBCEgttflXMrE81IYtkX7SCUVw60HZNHb5C8OmD+nUFwkcviHLTnyLgxkaJ
rOUQ6Dk2AzijNyUeHOSJhTmjj+e6Q/ELZi7txh/Gz0j3IaDTwPIbwt2XCpjf5T3o
bVw4V2jmmHz8tUckB0ahVneWZ3/OqfNOooOPqdJlIINcCbclYa1A7dbA4QmYasiR
cKkfHz7d1y6ur92Rz21ivQdf14ygawd6lwAYscMNXEG57D/XZukWQ+0VkE3dmstk
/lSexk/IWNd0kyYeyyUBuuRLaa31NBmsnsrXS+aKEVPg5b5PeIfVPf4b4TP1pub2
20EMEJwi1+TyZXg9EZwqduxmQYfzOv454ItUQ7NmIkfuid14EFaTy85Z7I/cNDKP
aQhyQVyAnjdTCAaKamQPz6vY4IsK/8L9l6DQJ/+nUWArRPqgOJzuW0DaroGGC5qE
l5Qs76mM24VOGC4Ht5neAjsXtaYUuy1v53se/zKZQ+nVy+rASi4dKKZk1y13Nrhj
lBwMvN4u5SyXISLtU/lo3lCewXapHGZO8jFCE7LgQumyvJfiDQlHZEdJXR5Dm4zy
kilcUv/51W88mKTKKM/1X5Of5svQD0uzf/cfd20e74uNY+s5rlv7m2RMHRmmoF23
PtSjc6I8F3gTRphc+IHZYxImX3RREGN8qGmFP189XZaUhwADUrhD3rKYCoY5hnK9
ZJXKot4cMl9JkYuPQxU9zS4fA+A/3oT5fhbAZ0XJLQvjTjGJ8ZG2IjQ6BY0+U0BC
JEI3Db8oUeaoQj0mctkR0M5Vp4jsaTv672AumJiAVH/fjaFukwLmMOckdC0mdlb4
/62BQ3fZkR9ZUsl/Yg2hPrl7kHm3IciPmNT7ItxIljtDpTgNAfM6D3m65mIuBCiU
oBtB6W1ZT040/o5bn4a6MRNCPJKKQXPqtbFeaKALLFnuOYKWO1NTTs/NowxanZrM
vpxyKzk4sipy7Q6Ax/sYwiW7/NMrPAPBo4Fq/fCTgLVWCsmK/m0d9mWlSQvx3sFQ
1qTZ57uHm2MYZKJR8DPtmSOQqm64sjjNcTlbgYQ/xwJg46zkr7WiAFW0ys9lOuwf
NZbw7Zj9E2ujPpQVucodYOYu6p7UYVHkWq6YKkzhR2i/JZ//ayeOk+CfaPVDPwoq
WwiaVtFHoMMRpYSeecIGJgt+6ktWDbk1ZBqSO/PhJxGm3YVH+hcqyeU+pvfoI7tt
puxufgTjAhhDU5hG7iMyDzSHGKdwCjMmaQKZXZGwTtC83dYLTFV9NH1MRiv4xuXE
XCSnYln/L/w8OKRs+97TsuY5J/xxV7DaCf8dk+XaiPY80kNLvxS23j1s89AvP3vK
nCvsIU3/8FsJ1OL9k4HNDwq38ASMJNE4vcrF17KthLyMkW9zmFNtzGy0xrajdmnN
PYs1bxKBV6MDPN9cRS3oYpnsq3/hhHOXN3WullKaSfLOhE7krYK7SL4bZgycdxMQ
eiP0+BXZRi8c3P2rj6hENCdOfLrgU0zYwxmu8VayRzPncb3aKP3n85J67DHohQPN
twGbLMtF1CMke9a7A9t3PrslOAS7X1pR0w1sDAtvT/pcqfpVk/jpYRtMCO/wHQEz
qn6UsjMejriE7qY3HWzUVxSp5zsYVMi6Q9xUTmkvC2PUXr+W8ikkPDZr5I42wJnv
iCHUy4XK7kKRfhsUmViQatbT00kFGi3KkUcy4t5n+FrO6sxHAFNHvfDGbbv/uhzd
6dZTUG7z4nIbaZZKcc7yhOb8nhr/h97rGy+fPVkaBdRxHiEY/9/WNah3Jk9ZsIFR
zBdcQJHpo5ethVOlFkp4fyHXZnu4AJbLjCr6P0TrUFjAqubdm0BWhnkDcUf96yrt
p/DKgW/oHZZWXk8U4QD7iTV4PJrUXOnm96RryJKNd5MtetJRWbQeRjHR/aQb18wZ
9RolMpo/i0l25XUF3pMrvKCBNhcwAlXbKZIM7ZTltFoQXWFNM4gDDdFE4L9eCQfz
97WsV1MT9b4gma+G3Y5n+UtOZ6ZKGAzt2+20qq4227W9OVxFmbdiUAMSMHL8d3I3
pVSng/0yMGa6LpYGC9ceKvEkYG0w8Vl9E4YLpv6R+6W0QkoGaRYOvKbSsaySepL1
Aiq9NgrJfy5BSfqAgA3QqsswTcz5v4onFtWvefoIFWR9CiEUwd3SSk0PVGKctFps
noXbuED/EbnsoqZhqvogIIpYe9LSQOKvlpG1kaqW0XsTry8fxq2WDFMEe75AwALC
7uwiT/6BqS0p7SxUC+SvIIJZ3ZhUcLM/lJp6dSjX7QCERYVRh0LPQs2DTxQ/wptq
711+PnouEvYKIynb3fbqvt8FFdXJ0B74IWq1Tjrtoyw3Irt6wPHOvfMWtykfNzi1
HNF4P0pQIzOF3l1eU8G68Y9o+GP6aopeuf2QBDnrRGWwWB5UKtQxIkIZULHY0HyU
AIMZf4G4fKHmfIPj5tU/BFkxDuSbmt49/C01DhepMGISsyWQa9HC/Zyzr/RzjiL5
/ZaQoGkZfIqCUwRjUA/iqered9s7MlJkzAPByB9lSvT4ur2Z93skp5W+hraNnx/Q
0d6cYRTcy1EgOnxwvBUxFYKof8fsHWWtHn4svEuiYeEI1LRPjNM2nLNynOCy+8uQ
DCPewyAM/Bc8ho9gmBXH1CFDfWlQGwFFUJ547dmkLyyAMwABxBY9olcBsv4fR+9z
HBwRZO/RAYqrl/EEdhp2q+n9/9NgWmAGJ5FaLTNYj5ebVs7WwwLk9wvFFH1R5oeX
tMD29F9fzctt2s3/JyckAFe5Ix1tcIXhIWk843baEmOv1XPEnJcplKTqAFgOybvM
2Pm4e8BM8yBlUB7ahorOhd77WfwwTa1k1Fj34EKboVqoAd8DU3rOdwT2zVB7lJ4x
W+mOlJYarH4fhI3PIsq63d4Z3CkAiQy5GRvFjxn9GuL5bduxa3pKGYIXjXuRVrS6
zr9fxWd7NRUKeGhNiIPmKxMyyMRzwYtzJoI1rwiSAGEfUoq/pGOK4HbOIokXDp/L
Y+zEIU21oDTX1aGJ8URR5j8BttKBmXQglHYRWbc/knI8ub3ZJPgcDK02Zml/Y/Eu
a9zdnDNyWfw3maNLfNUzdNqvFITKoA6EdmaIY/tB9yaPGBB0bPMOFQKOkI+mnQRB
zgSvPONjs1TBkS/R7HBTGwURbVDYePYxOufiDvupJAcjDdULH5lYa9MmbsOY+WL3
ua5PkKNWhokLnnT8Nx6TAGn+ww66Ak9sCVi6RFpwl0F/qaIQsRHNX2V3ziO1dDPj
EnBBuBtxv8n56Xc8bJxJxVdxDAHhaDAgCRhrRDQhF/r8ZeZVRz3Dr6Jzl262AXF7
UpnfRiLZD4cmv2CFeWCwX924hR8i8xdiv8PH86pOq5sb1SatKrkvYaOBfrgAIuVk
9ucCBaI6QXAgIFxmoaiuGnX6DkZd8QKB87k9SoGkxEM77R6HyoDceMBu35uHiHm6
oznkkoL5aFXxh68IZMknYtnAVoiygEuBUeOPd5Rf47mixJ1WY175+/rRnExj+c1J
EP/BpM3kqee1l4Jdb1MC4lE8bvekrQ4XOa1mF2nTYbyV6XYVuefjJjwWypBQQ7P7
Le0beeh9gNDrScfSqqNQ8dLu2j3dEuLzqWVcH5TeX8bY6PXmVbqGr0AK+6nxA4Mj
+4WflPNDcRqu1Q1v8m6QGhRIeG9HDAhetMXfSJEZeCOnXeaxtIsPlOPGGSLQVgDM
eb07h0Pj/LneKNPOtgUGl4k7MU225tZXZAdeIPdWbGuoe6ZN53kkn2o8LGlwNE3K
fNBjg9fS9SAxsdRr8aFvj1soL3pr/iy5ZL+K92V3L3vjxGKUmYTL3iKvAKF97hoK
7lKbEpsBTfrSgwR4p0sm1FwO6Mq7ngMQzqhBQPdlChDdM/JIbpWZBo+dxYI9QyAZ
52kfkWuwmeb+ugq9Ngfa8euLK+tXyqPdcaShUXGA5P2Rpo6WYF3Gf/GKmXoakx6K
VZdsZ9pTKEejRff4dkiqugaas2lGajBSnrm53zoi+3VbHw6TGKz3JittKowcLF8T
CXswE3Pzvro35OVUoDq4v9WYsVQdR63OtTf0igbvtofLPRZwUA5su6RiXkzSPfhd
6u2+sgCS6jwRggCZkGgeS93cPmhzegoBjjzcoS20skIFK+TnvV3D5tmqwbpjy2bH
geUBNDF1RtmkupO0/41b8PI0bMWLkusa77dSdFWFsde75DKPzjOgJwm/3RzKPbJ2
2wXIh341QIChqw2mtG4e0zmPJ5DebioLZcy6iJ83+1L/eXTbYMC8CrWCIDrKx5kJ
SPdEzYq4UR5swTMyqC94gMhmLlkhT+2JX3CizYqKSUuIeiU2LIyTbY0tYg/G/L6S
9qGnzfiQttvd4SXfYEarRs7U7ObQwg/lW98dkvA3r+nEBQGMfvg+RmQ2W7JPpdz7
59FTnQBdzKCLId/Ab1/osZ6YB8tqeQg7fKNioFpWMHL1uDT9g1iwowqMJsN3eQcE
Uv1hvwRxZikjIXJLE+8QspH4fnJgbW1q4st/NLMBYCb3VRZ1MXThT2FceySddVw2
4Bmju7kIYIXUy3ii3BJtj+uduHYveQ1OqVG7qzIBVAlTDQ1UoSlQAxke4rMciLD1
FYXBechTc8uEOESzNVGBhumotr1DhEfRj3D7fNmgFIadfiULao61NCjaA7fPzwx8
uCQKd5XcjgFmnmrutNCwE63x9e+ALjvhf845oNJOI7sOSSil3Hsb5pPTXD6TVeqK
el9BpLbodEvxQsu31kmY3WBT6cS+WPus9/bWrK4a/7HHvHVALHlKBhhv/tJdL7fB
Xf5hiepvqO7rHaQeaavvchm6f4GZIUzRyOXGgxSCyGnAdx7GYYK8gNCSTomObIsS
kwuUIEC+i9OkCLahkPCEUXYe7l0mkY2LS5W7QkTjN95WBe9JTzjRMH6cmW0x+i0P
SwQ9fA/QIdeCyXevHJbV99yD6hw9d5GuxK585vgc+C659YGOSZBmqED7fyOR6VC3
kkQxyoQUpxbXkSGweeT+7x5Un3eO0bnESRTYysjlCCNNNvfaN1sAOSYQq+DdHKbc
1A5phbLZVZIZvLF41SoAbvoBdGnpxz3/Egz4nPcgxFZCN/RsFjsxB9n82we5fqcw
ua7vuigKvjIT5209lwonkmOrCDVcs9Otn0WgJ54nVunoXtORO+lAIuEKVnqrwDRl
I8QaXiQ1UIJIhV3HOcSuHQ1vyIQI1/TEyh6zH7ggLORRz+FCydgc9EUx1oUcDBEd
yk9zKNmOLfpa3B1lDrBYoAnifSs+C9RUwyXuLOYfnrQcYhJuXRs7XZeg6tSrgvZ9
ZMxjcPE7XCsMnDSInEpGwoFSmx+VbeWM0DOLOuCFMcWCTLMTqpAGODKDAsFOKamD
UZfcT4yvVTr9SCZWZCR1dx7w6sRBAYa4zJ7XnovukV7MZT/IhnLh9N6hKFKv/vXL
Fl33fyIIKMmH2NdI8pCNnAm74TKE/bbldzAen83zYfwJ79x8pKA53njHwzr6mtod
TaBHHAQZ2GUWxdjJ8d+bxmUQYLRLprHQAhaHvJSJQi0sRPWpUy8CgDro9XK3hncY
3GrSk7KhgO63aIgPErpW4eBsW2NoiJlSXPDI/pBsvz5V34+lT1FqrRt+sO5lJG2I
IUqDUaE5LMlgQasQXpkyaJ42fbe5/Mc9d3jmZsLR6z1Zbuf1wxyl+vKwzgh+n8qT
6Dq/vQ4gFeFdNJMEZnSuGz2iEBYN5em7dvK2SQDxpjWL+qy3xrI/06RZ5+qtj4yj
uDXWfmwNcZ9GdKzYn9caIDBC2/uVaIAgKrzscbbSFbv5WdwEDzGkYMsgD17ZiHmn
8z7xME1JWrWAH9kt/+SrLUIipKDy6MxsGiJfTKvVLGXB19vdPqXGGrCRS4L4X/yf
VmU2Mt4fAcGnwbSI8I375LQPj+s5GOqG7zaA8Dqs8BwTWPt1QuzBMIjEApJzo/Ms
obdgAAfpQbOfzJ+M2qK3hZx3gXt4IA1gqDILUir4J3Y0zp2vgkH8+u7jVhATBMVa
uKt5kJvJBaLDp6ysMNsqoyC0DGB92ZntxBzreKBTrKc2mYmDbq5on5yu9YjcY05l
sF4zYvzGPY1UwEOuryzf691MxpUB7liyDU6UhSdYJPn/+WmQ9S7CVNBJfGJQZHp/
i3U8qIYGbaS3dKHoHl/H0TklwOCcbSQ7V+z4tN8NNtnIxvEGN6WHiNm3jOW9IX1I
g8helF/4/Ct/ig63z7u501W695VROVWu2M0iatt5G319n0JzJbfnnkVGbp5OS3jD
wwPHFaDVDjIFDLQ/LQtrg06pS4obyGWwOE7zIWCcX5r6QBUfOrzMojtnwb0dGqoh
zHaIpq6E7cDz5mibGOuVVo1rdCcJl/RPN9rpKl0FPtGgbSb2o0k77vk5FzHT1Y3G
6a47iW70UGe6IucD93pWCkvTVC/GLxwEm2tTPjMFHOEdTkRYCAtEK6A+TR3brXTG
6XGNXSC0hGV9bbExy9/JEy4JhMCWNh9UHa4eddKSCiWLhzqxC59gScY/75vmHgDs
Vk3OYcESqjrZF0iy+HyNy6mLsZsC64Cb25Em32y3jAnhpB8upZJH/OMJ8XFWS3xW
7MT7eszi5U+iAKSVahyJ8QkWqoQfrnrCinAqDouNISXig+iCvMnyvhuUVdi6l9lv
FWtzkvcXVoASKDYIEf9e7GkzcwR9m19uYs6cJITxOyQkZv9lP4SYKaoZHJoPcBQW
VjW4AtMzjZLpZvdkElPNiBV4vwKMmB0e0nz1ffyo8pDxGWnP8FElUEzRYbo3iR1J
gRzUVzYFqvpmPdUf+9jBw2F3AikqQDIAU25p3PwgTuV+FMCNLFF4QoOfURVLYQHf
+jyaB0nZjMh14Q8vReWKXjB+LZdxNcFnxBrrDA1gFa8a+p+citf1nNQYXSgC78AS
HUDpnWZJGRlQFg9/qEHIgYdTe6HGM+a5N/h7GTFkOdoRn6vNIAG2g5Ju7Ti2j3UC
f56L++DWqNnvSeNq5A2+kuTDcoW1u+aBPdIyNabrzp8uR/cKTnSZoo8nqYPH8wFH
ojlVG+gMZyRyNrJQ/co9ILbL3B5D4cRJ2Jtd9WYmDBg/EcxTIXYtO0CySgv5i9ST
4dZK+RimPccepwl4Y1JxK08415M9RevRVVrTjQYpfvsR6g1Pg0iznx3kzkza0yhX
MUcGvbl/J9yveA5xtnPYakf0OrpXBdmklRUaT+Y09zH/8e/iIdfdNBmI2GoRNF2L
xDDWmZ0JHb1FaRXQ5asX5CYqd0geNPEo8grTYoJHUnJLq186brxG4emkL8ldhVrw
RcN21kFhjldMitrTORqCa3kS4hpHP+Cqc/Ni9FylrcNMJG8CCq7mUzaAF9KLV6NA
voP2aQpEtPDge/m4UaLqmGFiA8KIqlRLOiQunsscc0Mkx2U/1xyk1LV1q/+Leqf9
BZn7Zro/DoSrmoO0rv+G1AeZMGVeOD2zDgfQrMGryvrQEn/19aa/7zxoO/sp1Xxe
uC4/CLEYF0fv+Kg7JCdGgQIOPOAaUhgwTDlBhkufUhx9PCaqbKm0b1DoRKZbxkMC
7xppbi2ymMrxl+JIYm2auPUwcMyZPQa3r2eEe/nNoA+iIVARRW/7x4GLmRO6aWxi
0yWRZ7gzqzevRM23sOPk/lOv5mFLXsBw+FbA3L05wZS3dmbXLRLdZHSjsNdVqtsa
twUeDdSstbYSRt2uXdxmBKgYOe/zyttls5ONgnJhihFdeANSuxBmCO8OC0xlBvOK
+EVEdVpmIE5/dRANQ1sZoUKN4P+fQRf0G/6RW0N7z/5UE8UkdNmVK7zgNmVzQ+nv
b1dDM/cfc1RBcAGNYb+7/Z1PzlHLZcnt6krNWPH0mbTnbGKWEdxKMzzqM7MWOmkc
9MIOnZG374/SU3k3tVknZhvyk/tNfUHFm4fMHGZn56ejqTE5aQnGpqoIhKu5ylfm
YWsYmj11shiuShZFWJqtrtowBMUcj6WhM1HH9da7N3D0Lvlkw275F7StDj/ZIjoE
SgEW7J7IVlQupwgftEqObd1OyggPp9FkeP0ekOT6RMkq5u7Lu57plgUeRYjX4BfC
SWOzo4w95nqf9JsWbxJryplCtxEZDZVWmC6Fhcr6JknLuoYjvLK+5GCpPh4bhMFq
LjNcMna5ZFDCYdQMEI7H1JbtQTPb4HOFR6KnvhI+BZocqJspc/V4RE0ZrS1la245
md6IRrwiG8z2Az2xpaUmURt22UfZ9NgM0HhQEFJ5KdjvAUiaqnwv9F0DuOOtvxYO
6wa1IXsgPTzcSJKrFikPu21idgv1/BW967oMN3i1mBesh0cO9Y0k8x9GpsbuKmzJ
4BF4nNiokEWPWJiD4Df9Rck6Qu9MkwguB6tOYaF/ptmapUHC25B1znIfpHb/P7pK
U4kycdHIJIyh54KLi0cQ1QCvi11VyKA1L1QFIUd+rmCEwIjCAfKZ7br3fQRUxeMR
fnOWXrOdl15sDPn9zHxBoFOlbwx6zrd/b9SBh8AymHsfMa9YhVUQ6uhwx24jmtxa
GWFkAiITJOobWmyBlJnwoaUXvsuE+jwqrsYeO4mHjy6RYosVxLDDZbQl1WGnlfVI
mRakmbJLx34BSqkBwo4Yga+ZIxVeiYXNYrUa3UdMlpFSiDSPgjs5G/ngcZWerNE+
Vrgyd65YjYyWulxudNw89bMj0gl2AnrFs29evU4xwOc76YtOrnP9WTkLqcBfQGqI
fQXrEIIEWQKXfb8aejTXW5m/ikCd8Q9TMFrL2ziZmBB/JzIFZgLzrVLeu69zZvCj
49U28RH5irfLQhoFzmqoEAC/OXb2rSoDuhWfRCOtmD1yMMmQVe3yqv0597jLoWG4
QUvhr0qijbfbNm50ke6tlFPcPpBl3jwajruezE3UG/gbYGjeQ0cgsBcp/BGHuSt7
DXrJUpAHq9UqGaryxsJXx6iVc68depon+TQigvTdgMbLI2Hmu+8FlFfI0qkcjMmK
VIk8vmzKt7QHhGzYZ8P/j4jexUHTbHsDKFfHwhhKN5u9IM4immwhCWX4RKLrBt7n
Ht4BBqepCkoCF432zsazYAIS0k53WH5DNRxqK/w5VqnP0/CDl2rlVU333cHfY+RY
bWF6hkONj5dkXYVGLAKGliTl0taq8kqGD2+rz96gJI3CFq2/Z8LHuCaBRt1PEdRZ
C5p7w8I2iHZNY7Rv+hhRQKfKOOatxDv5S2K7mnIC0xPMIh6ZCVViRqvHqSAdIujQ
hmC7+J/uDIUgtErFGm4bSZlYglqzLTX6NzmEIG24rUXFbV93w9Mk0fKR8XaL+F9+
nQZoaRP2wXhX2qPxBum4mfd0PEUm7TPt+hutdeC99ceG/6tlXa72KfQvYMxyZCh1
thvNxNS+vLK3AFqrQB4oRX0edIOvql3lwbwAKQOLOlhDcbpdAOQQNLGou78qZc8T
iJPlKAi95VFOVhll41H9npwBdCBJQGjUJyv6S0jzkv4CK4FJHRNe9yzPHRG1t/yx
3bvjlu4xdwXoHg4SGAEVr1N94dbLIZfD2wkyuQC50O69bTft/3+9g2WQIkiJNhAj
lS2RvNATDH29jdByPmTMz+bwUjggE711fwHxbTTyqKo+phM3oIHyOvBoWD7fcL6e
KZg4iu56tWQe13U6hnRvD+vdlAu6QJ8tPQwLHvHtDZ5QWCiNoZwLeYsWl/+oxwRO
7aaeatPqLXA8M76DEGC+lyM31DiKoy4P6iZGtlpCRl0rju7NA0O6BrvHpxzLWYxW
1miJi9++F/P0m3ZUQdbBA9QIn9KMGdEUvI923ThWwd5FUT0O31nohpdGFZZqkOXz
wgiMMRoAVfUXeLGnNP6mYoYds6ix8tds2i99cEAVZUMqSSx9eP9CEABQu1jXs+pP
j7/krUtMT3IkeDNj5XBxhi44HkNpmsJ3fDVkCeXFnf/CakcxPljUvTI6zZ310hbI
S9dLoW+QmV7e20NcVCrP5P3ivJmz6sIXGNuDmQ1EvmVfYDDB58A1+w0lQ7TTThBf
Zbs7D3kWq7w96+po1wAL4/8Di/x/1U5sPeZHQuma9TtRF7PNglcuVEoTFKwA6Nfg
48ZE2/fdX8T/DlpBBvIY2L+kYSofaFQvbS+9Ed8HWRlximL1Mj+3U8Flq3P6SxTB
gnwxqPmmbsgNqB8J0INMZXMtqx7wDILBYmDsrqApDvsCkJOnF11zCvieWoDOZe4a
+w6hk/13k1SlHenJgg99uuoMqxX59NE/5YSiLb/aTIRzJjnZIHAFF6M/qXz3363N
2rcdcHWcNNdvN9P4gsPZEec3We6tBvQWCCHfzATgXZraFX3RP+FsCx0PnaMwQegr
YVL5NS44vGAnbyfiCUNCSHucz1+OyflpKOT0Ov1f1jaNmrrJ+9p7fECJBJlQyuoM
eo+MwafsRiJCtMPutsglIV6190Uma1R1ilIaBqmgHj/cCdPchJzEotj8yA1WATCz
CjEuKEmDaTkb+tiKBlm8o5CPVSrsWfKMdr6oQs5aMD8doFESBYY8Bp34/PvwXTxZ
uWBkTyj0MTC2D/iTkTVvDhAzA/N6SY/kCv8MzNYy+tmwYVLinVwciHYJIaAmaaBY
vhOL43lNSs6Tg8ky7gesqSV912lA7i5D1hdr7HJ0pLm6Fls0dFamD7sddq0P8CY/
m1X8R+HZNkjT86l9Hf8g4OJ2kIjh21XRh25nfL2Xst/h7pR9ECBAPtsRsfAlzN3M
jogwHsS9B1kAtjxTP5/TWFgrjlL67lHfAMX0QRMXUAdV1bJjtCofpHcb0Fqmf8aC
N3ppsW6AdwvrJOUQexhZOqgbHY/YXkkJTu24YQinZCmynooNg9zPDRm1vhNxpzhb
bQ50py1EzvwfIs5UhbKH4TfIf63VCSWfC+LyPszWfXEPd1K9rGdJg+8Fc3W6iw3z
3JQORZriR/Fb2jflzbB3wwmyqWv7BAwyiSjL848fUbVMOF3jyj/YWNbgIkrx1iIj
xlZnwfYa2s9A4PIlJhAakJY+eUUob8wupTyTDjF9NJEZjJneb2F2OAHxC1AWzaST
e3+IchuWceCWWNE1j15PQW2gprfRjzTcu7APEFs0ro6VYUumydQxnQYO27bR7d6S
3wT1PfKBw6GlMh3TcAiwB8BJo4398HSFFMietsv8ZwSk5t6IIqDrlCnA9VdNEnUq
j7aUGdEy53duB8J0bIw3KjUhRVMSKm8pKYI8bjpE6ZwRHzz/JfEcyRBM7FU+C82i
QjBYSix3P7yjmBb16IeBU2G24n44K9Md2xlGKja8cQHE8WwdI87nsxeotcJCN+FR
Tp8ZAf6GclIwQaAJHkNCsPeh9vaEPt+wtQT46oG8bAmi68xxIKYXv76c7aO1FN3c
2cZK6pTpJunucOATiN762uQftu3Neru18/uAQG2JdItFzDRB8xWMjVSo1Yif2u5Q
PhQ02fA6t0H/iDlTqGvkZqO6GaDvhpLrRb4p0iWwdsKY3odRbr0w25lfyJmq8rY/
bo0vM9cjTwrOU0bKOQTlpqA1nxki8cnxptzQdOk5bA7d2SAhlhr7BifsBYV0ZbOI
QvzVARJUhQ3czvF3u3ZcQvdGrr2XJWEvwsq2wQ/x0tbaKvVot73hz6FFOLNH6ETo
hl4WksYBsxmwovFlZleVinQCxBr3Sj1l+ar1XWhrWJQBMIZpu4xc0CR6p3Be9EmC
OCz7J79EOxX9QNhEIdI3giAiuAUCR5q10SEtooKSg2KS8/3CDOPCt+R2WcKHc8or
dpmsmV2p2o1w0A/LfkoCIt+nYQJgle3vrykESWUmCSpPvOV4s88ExMANcO0+1LpX
VC+vj+ouuu0Fgh6zOaMopSrHZ4KUosRuA8BKb7CUFTIAfW6SaK9Mxm/U3sD763xN
IVk1IlJ1XRX1JqIK9uvTCjR/xBbDdsX9OD5FmBYXRbnljVnQBLKrSrnSsRUNiEOr
Pi4rS3iSlOGV4zQA/KkdF09k+upb+WMtkJnDMjeauwBp1a+eaDZ5SHZKP5vSKX/M
aVnqdWBSVstV+WdWhJCUF2VEjpOniYqijIl9p6+uf2MsGHnL4dlyxrzxnJO/3meQ
JjSvL4mzVFGi07KCUnBCGn0qHWi9ttQzDfLrX1EJ1KQ4rrnCKdLHNEtRgghUdhAa
eb+O61dJ4uEv/Bd9XIPQUHTjm3yvjxgCnXinuoLLwzYRe1lTBt3lhUKTuGZ5rpXv
MrYNY6YjHdt/Br33AIgTKR7q/A2WaHRgE6qXozp1xDgXN7avYsltF1ceVko3V8mV
EDtmN14GQHQqPfoo/37TS7kcXbQzj85oRRAhx+lJ05JTZzxJQLkLhLC7zD4ejt4o
StJPG9ZRNpbozOGvGyyC01ouPrSqybCTyPKolIUPITPrr2vA8Y8vNssTbMWXdaZw
GuibjV5f8miZ2LyX/nq2iszzTlUQikmFcY0D7miLLMfhldjcKTcwD276Lc0P70Sv
AANz61fkw7FHF3C1GwSG57UsWFw5KVQFtcYUwAI5kAByxD1ZY3GUpCgMCnkMg5pl
ksf0IoCwHezIcye0uxTPel8POwKYeybekV8InHoZxYXEe7Z55KGX9uY4hxn5ULRq
nnf3Y0bEkR+wA4d6X41Hc9ITlqixh48UMLwI7UvWmxyB7sfVyOMa0SQcYlIAWkDf
kLgv82IR3WGHF0G8n94wXHVoXu+i3sUuv8rBAqqLzObmpsGjsaptE/Hyyj1m+h8o
2zgEUNRBJS031+rN9baIZeMNDF5VbK3uTAfTL+izh854cedB7ybb5mKWBP8fEO2F
Jhku9v9XAMQYO1bQee1CKeGS6BGysQgtGcxxciZyk1gc1PcZ1Zww2EGO4RrdGUBd
LFuNK4OMqo34Nd8ySO5s2AZ352O4giAljTzaks/3h6DLhbKwbPgsUqqEbyzW+20x
q6VF4oi/4CZHg41WqmCA6wmGkvUbdMifdPXEPafFMd0Kbk+XKiW8WLW6Mri/in6n
S1Npimlnskr1jgkw0SCLo7IyxMOjfypOKfjEabpm7VkeZPzSttkwVizbaqE/4po7
ZGaMMOD8xLDHk4uCGfMcoVhx1gwiFMITMQa15i6ObzCIfNamt15/7+pY7ZUCG565
C2V4jXWxFd/NDY3jctG0rrznHDP9tn/+mOra6ekwKFuqymy39FRcxa58UcsCoG3e
Fz+m2hqc3EZBqsvOwf3JTxP907dKbAuzQE+LnhXLi/iGhFWe4aNJMPdcY4I9jerZ
HdCuT26LOVQ7jscl2OwIOHL2XheR9AdM/5Ctqvqnj+XkH6hE2pMll97f43zH+nEb
U5t7hcjxZG9mGU5hhDfhDqkHPOGrKkhTsoPuCcBnU7ni58owpiuwURom8Mz+zHAJ
5PNy0fo4LkYpnFTbC7rqzpzPq8wf72o0Mq7FQtSSqylyg2NpoKvsPlJbgWoFEKBe
KGon3VhErDQu2URQLDER8nf7rqLZlQMKPOrggkEbbfMncluhYETWft0dJ1rgDvQm
6LP0qJVYf+g/goZqKmyryDdiKv1QSjvoMZClKCOg0V3k0H7WMpBbYUZ9kqls0D0E
VTJgtIen04wVnjaonPe5mUAcTzq3MCaZTqB1pELZdapiszmWsVl0xbQUHTY0UYDc
VJvZZcK92CMb7kmFltNN7TDnE8GKRpM9rYg/rD4e2pW3lT9yWDqlYK40zl7zIuYf
WPHOMa+dHHeWhekwwxmNvbWEUqUKOZS1+63ryuQMFcsYhWnzK95laf6KfjQLd+Bg
9HgHLj5PCwsbqhU6dMGBXrr1FOrYhnAbj5o0cXOBEzgURdkP2/RwsQhUwwmahFQ+
uMsE3Vk/6BJQddAWjT7T3iPxADSBWXoObcitGWqNqZ2nyuUU3Hrds9TKHS4aV3ZX
FC6W//qwey7jxNBJlbL2MNYCSEFrnOZmDFtFQrDbUb4kiv7OgvjZnWIyyFBDq97m
JG/PavEtsstxJZ5xOm3RTWsta4LZNKTMI+X3f7I+RCG6zHs51KBoz28WdwdqHypJ
C08FuiptQuMwuU/3OyhqZZp0mGJPvb0amMwxHVowDkhSEYST6JSwSeHEQkELYzRD
pnbQcx8nDukatwdp5BC1KKlJ3tc2cH9usqhXe1Wk253Hx7/NOwdbfZAq0BpKlKRs
cjGmGhpEQkBkpdLVVg8Kg1Pvmolg7ZbcQz48yuNjPCaSmFg7O64uI/ypyy5N8sxH
NvAP84C6ka0aGubuqTFMX1kBeUkX6WNKn46w9m8jsdoPcVgTGWlK43YCg5AlgYly
w46iy+GBfZKlCTqkXz74BHAyq6eJVkqSx0Ud4ENduj6tCbhbu4IszLD3ZJ3j7NU5
SsFI0h5xgdd1fMyHqrHD+aYJblrNKLmLonlFudWZQ0A9uffj72wbgv93eoXVHnM5
YfcEkPIBlMexqoISpyS+cj/Gf9Y6L/xnKrxNF0da2sQGGKybGz16QBmY24HyQiCu
S0C9mQWUy54WJ4x9j/SxONhWkNMyOkmMXyeO4sbQ3YGfH7AkOtxSf2b6zlXflg4q
yZVh8LY1J3kPpYB6CVFHaYfOJC8mRA09vWUMopMu+qZRryowvZDspzkJLBUu1axD
2PIL0EldUwfFD+t/uUmsXm6XHT5h6IAZrd6iYUgnYzi64uxr2FBtvj3MXIANVaNF
KqgmyPO2TE8kQ0yDqXzZt1GB9A71Xon8pOuWiEFCT396ZOZIJ7NulaQP0zZ3jKO9
eqK7EVVOxmg2suGK2lnYOk47c+Y2Ja8RkS3buvi+Lu3QhDoRfrQ9fXEmQcW5qPnR
5pRxqncoL6EH/MmD8gaHgOyrR5R+meMVvn0H5MbEM1Rzt/sukm+kvfTJoBqH5J6K
ypsoiBqbQ+vsy478DbPVahFPpP+5EjMI0MKYTM7V02XLhh8Lqc//rqKJ6ysRGlEf
TcndD6667Flxz5SQ6wIZuL9QPy2PZOBqX4bgYUZRUmgVF9DMUliiaWiFQHHUZZRZ
E0VpEAwhYu60SIasiEomeI9RtISuktkYQsL/qiFVjKFam3uqgzw1c6ovsiJJ1FGi
GyfWIFAx6uCJqyJcTo3my8Q53wRIO9yA5+cpdefsezuuc4fLp4WYx2rOp6LZXofB
XUd8rzjNtFYnQG6u5JkGGtI12CNFCUR1Jmw8MmsFOZyfd9ORyZSWrjC01gpKzPW4
hBD/JfG8QS9DUFVLuNJjR4+2kWKf75ZwGwYlLuOnZC1SB4Q3TAMDUe/xkBqVUPJO
oTrd3SURE7SHeMHcof3qiNQnjG+cXNoB5DFDMGLavisSDo+bZ1z06w7ib1IQTHyB
XyebZDeOjLaWdz+qLF6WQeiZUrIrIICLzK+pWjL95tP4iUbnl66KbOh5dFVSra7R
1002OQZCjm3YyiZPaOZSq1SZz6YwJnR2zivJIE3W2rqvwhzWEIwIW4hNDBBcUtdM
4UT7kEzoOELS4rbPV+kiky/IlCinw/y3OvxSwdOabFkeGheagWGoav9BagGm1ekI
BOqnHFJzJHqdrDohK6aBARSHb97g9CaOpQ7hHvOYGZoDKJMsEdW9l4bmhZLpq7FJ
5CL4fObW4rz19zG/kuvu1iw+GZTAmdLIVIX2Rci/npx2zauqF/7HlSVckO9zuPgU
KHw9MHOUNSqPYdU6ibBV/shPfP5wFEqPZMrzl+FcLxN/uX8jJwEgjUSQ+vMzX8cw
2Az16FjprHOTUz678AwGn82Cny9BmKuqKHCm4L1h/qurbhgK6YtJs9WWQa+LYU3+
X6QMqVJ2JyMyc+CesQM/QHeNcU9Sm+XuohE65pE9anRkMgW2PBOKnzdkaI+7PlZu
d9ec266jTmcJg515dCNCtmRLI3B7g0R/uhRxVQySeOoNz+fGvdfT1TjfZSYfmqPq
kCoRKk6tBqWJ5uLqkFbnw2oIk00F9YvEUq8N45zvyLhoQDfJ/yNzB/+Be16BsN3O
y4cZSpdQONk9lrjUgq6kaSQkm2Ccg7E9nthRZnaZzi4QHTyHhlyIIr2U1vvmKT5U
19Dg4BN0EzNPu7OpzrLUr+rHwzasER1XDc/X9xnOJQEyVPWe7E3T602MvFEvNg90
mF+9JowvpWKYNa6PeAdJlnCUOZ5pyogwaaUdv0viZR7xXMRCwPZRkteKxIV045b9
GUYuT2Q7stZlxx6s7repdCwJPwawElFTJcboLzTpKyxc6j5sKuqTldKuOlweJHm3
YyT220NciLRHk+EszNCZDSLjxm6rIwI+wTZx/VfKjWqGqc5vUauSuHS2yJstQ2n6
zfxX9A0g6TRQeAYoJojp69uqmMXOSd29xxk4WW8aTdGAwiQ2Crw92R19cJQbDZdJ
dA6uWQpcaX0noDr2CdZa+ScKSKH9Q1zJmtVG6SiZcxDTU61EwjtpEl4JIVapLPSt
6euf9Vx4QMaDyvIq96ght7va2iHhOElUnWg9wV3zi3NF9XcjzDPSwbTmU13oczRn
hWKvyvHVafUsxChqiEmyqb5vQSaIfFVxE5L+P1FEuc+MqWuQu1PIKtIN+Htqsa8m
7GlktIsVZn3AlGSlDaT6oAtWWrgHOVC5aMiux05Dk4U6WCwNqcKvdZzpWmsZuIV3
wJEeowvv9fU4I0TtaLNM0l/16yopoDCQ7S0V2boNCgA36fuQEyX9LgI+1741ruFH
c5usK7AT0dDdJ/JeJ6yZcz+Sfq9l96tDT48u1NOfs1nTofPoYJzwV9zeDRn/gPAY
eBjJWAbSYHxWkyH5a5rXo8TMvXeCFPfShSOa7DY/g9l1HVa5gb+CHlGtPD7wglW9
Hcq9RuXqAn2ISxK1ecSxsqKhfp6KStGkrty7euUNor0yYdNzVQnB3M8Gwd+1xW71
3pWCMnVIIz8lJrOa/GUXtBOwZXRwGqe9q3kin5A5efwn2YcbAOwZPtM4WjLNyITb
boJaUV2MfejxLnWdDUbHYI7xzNuYKEQCwerujz/KLSZZ2erqi2NtFGCF+if4zMFQ
p77OFLGzi+3VqXP/5D1QQ/vUGyaZbYzm29qFZRBz00QPmFxXpg8da0oT15JRUXeh
Vj28CZ64UGOgHoF+C6opT71arQkeshfKk8hqFqmigQZdE46oupexZOQfYFXraUyo
BHBTCYCNyj9iRZ+Oowr2bdWVB+DpAveql4MaJO8yCapGGJNS4djEVdZmeVJHCSZ+
/5cI7J4RvkP4shRZxqSeroN2vpNhM8aqX5mlyr6US589P9I2NuDUqwQCK3HwQ/z9
iGdzhoBAeelX3bxiwh2bSkv1eQQ8rsAE2/Qj6lvzODBgEueKhFa7TZfqdgy4HFsl
8YsNeRTc6P3/J3X+s4GYIeu/AE8UsD9E8Fldy7xcIsRyM1nJkpoHjCAY6iRnv0wl
AWj64v9eg0P5MnrvoSoSoReqMfXbMQLwwyIri85KesvNX8acUrlUsP7NbYzlKAN9
Wl/fUhvFl8oJVESKbIX7DqWcy4vXEdGb465ariNxZkR0Tg4NVq/oLHGAJaSbVqQR
yoQmLDGg1t5Cv/miB24S1TC4f8o8lGQFYL73InrEZWQsFnoxQA4Wo9NOlYDSFNMN
oM6xbZQYiG/D4HYfT/OV3wq6nInsu8GTHGeI07LBJBwYmKuoI5GO2l5j3gityOhw
2MMQwcvjehY/hyRCPnZinr0+85ntwRCFxlLb858Mub6Nm04KGO2wk9i3NbTpuIrJ
f4z/R6ZqOl84BK+Sq8Lx9IkwS7GZpuH96qmCaQXBxeyXyHQTzR2YjXCrmGaW9yTg
cOE/flb8MzTFhe05fteJXohbP0jiA/Zg9D+RgHPSWkbZ8/zvxDa6Qg2rIBLNzQt8
XYoDDSyShNEjhqNimiM0epV1ENfZ6Q6gp+rU48peshXIFJoch7qiwcKbjxTSaVS6
K8fzIZMXA0TiH47dE6yMFwL6NNzDMbhgi+yrMw4iUi5c5GPK7aBba6K9UNc9t5mH
IIUX63SWYwxoxNC08N61Sll+AVtzCJjBHble7CdhAIWn+23mkdRFRoWd1d0JZSou
ySQfOkENfc1mLoiCTxgOQKrup2jxXk+8Y7DWB4vBUc0ZKM/H8Kd48WkRlJ/aREjl
rUtJ2JeNcQLpH9V+nTrLAgxz4HyNqC2nTqymtfbiKkgV1cTLnmvoqIFpkoKpUwPf
Bl75HjJmjQHGamsaxeXuC0Ug/1hhJDZzpwivT4V84cXsfu7dxn7mPxXbdqucjP3f
8zzOTDpbUZ4ZJka+un42XZ0eYKRgU7AAIAmKRK6jGNWvIR7R0JHaT4ZNSgr5ZNbX
kYgaBvzVaHA9tLqPJEU5pqXoLVDRDiY1xEAtiTX89YigyKs5s7ENLJ+EpHLjzb67
6SQOAAioqlczFYpOAmlZwJ70g/vB0JGTUXEhtBpnBn0PYGOsOViK8seJ6iLCiAPS
kHMq0jeuxc+xBoJUHXWIpRiSM4Z5qEZz+4TCJ3j8gJVHJbBzStjN6wB+mKs/PP2V
V41nA5y1SPM32SFf4+ENWC2NgmouAKqXKSzqxpCoul7wKC+rHaiks4l3YZ3Unl8/
Eit1l/p4girPQpzUF1hWQJ9iRFooinIrXnKg6OJhjtuiVkqk1qQmavV0JEPUDpFH
chssnLzId7TuYJf+sRATqZYBJfTuJNiOU3hqi6JK00HuMYyKnaddNVIdQjFKSPeT
MAJuKAFd2DBknb4oJTlWDp6i39HFZa7uYYKexnMNv23K+8bl2hlZLoRccj1XFv+t
8H3F32N7B+UKQbTI4GgYoMBuzxsyI/5qFB1vtQ/LFUgo11PiO3DI12JzfHOYUoEz
ylEpAYXXBtNQep8uRYyGYCNlBmgXzDbbxievVEN4EEiTiut8WDB7i8HUkUHNQgbj
b4EsiAUNixeOfYistzurN+ZfFgJRg7n/l2HR5u8qkqgu7WZDI8pH3OH7yKdam7qV
A1yUA03socOC3JzNRVQRk68peNK404wm2BTXaQaAPTMY8ekd4r3tqc+VJPgcvmz/
OYrOv/6/bD/m0INb4rthGshpecGKFj7MeJ9SNjj+JmGX4aBwJMf03nP3BmghpDzf
Ah1GzsYzS5fB27+TFEHHtLWcz5RY9kPMkmH42fMvNoewxQDdED4WGaOv5CMmF/qR
v4zIfobr4dSkjlSZNbWae++LRf+9hkDfDWqhOhKxD/lzRXxNJ5ybx1SI4OYUW3M2
aY9PVkB8ct+D/RnMdvDEGJZXinav9zY6T23N8HJsoNZcQRDXEsEHY0Ex4vMSgTX9
/iaax23NZhgCdYUTnlr5vHv8c3OxZ90PgkqCRSJBOyPVVAojA7Ihha+UaB954C1H
d7MLynZUebXSwchjQfUVrbSmatk0y/ZFIadzUuEIScL1aC3GHYP1nVJ8VdUoDXdc
jsS3GuDifWEi+r6fO2LplKhyiVlQ4VmIAKZij5w7EsSy8kmtQEpRYXOnr9xVmN44
zr+SM3pWjE0Zwc24oAj4BbIRwP/LyOzgmkMpt5pJUFpuDRdH5vIbqXhmJyxcJ3sg
Hy8r5rom6M2k14uN/t/W718uyo6KQaMPNU15U4JNkPKyAZ12DFvDaIXwo62Rjz+8
9DYwcMyuhqHX5B+h36Fc88Nmermb588MVPRlEk/zBscKJl5lYumCf2KHvggtoDI7
e2PXrq+D04r/4ftvVjVpyIMKQysXCYqVH9doCztnTYaF5aktBe4CQQTyAAhzDN61
E/DsQ/lRXQVyGNfq4glycY4yRq3eoo+J0h8tG8HM8r8ar8Sdr20CSApbaxZsDuJX
+gQGdC76gUN7Kd1xq13dSTYC/c0z7FnpLjoHBhqp9M2mSUeCAykwuCXbE2j9jFrW
94aKvcpoW+oAW+VoZAxVtVQJixgDyIdT+miAaOMoDjX3rbSHacmIfHatIMk6kxJw
p+8URzlNa/DSkWKa3cXoHRX5aa5RMrRoT9edMmzG9fXMY8imISrHdxyBnaFGuWh/
IPtkZNk0/9QCcq7OJ4ZtscDtOMLmzOI+jRgwPhKqAbKH9cvVRosQEdYOK0AGOD4u
8bpoz9lK+Hb5qJFAUkl9GF8xDZVsNJP8WNmWW/wzg4kK7RHg+JfGm7VhE9rMblBb
bgnnbwLkdqg1K87JplXDnG9mO9yltVvpVYMs+syt0l9Hbz129D0PbnZXK8bqao6i
Q4ott7TLS0pDIBUadZsUStTd/gD5tkLiabSCMSuw8MS9g/bXLY7cgGmTgkcfWqm+
ollWDCpKoqRaXodgh/ZT07X+Gp/YR3TJbRcj20nLLst88FTEqWMSwHYwaE+7ccxk
RSSuUFgbnoZDof9Y3oxSQ1Nc12klQAYmIdAKo1qDTOHtbxjrTa4wpn4iHBFXssa9
jdrcm8IszAxJUrvFC6cUUrLfxiK9nqWdqgEWK5MuGNILhwYe78yHY/+StUFElXo5
n5y2Ritv+TSrOK3vTFCQ8S5usEyZP8Ex0xkB6EhfmEnyik7yQ1VQRwrgcbLLSVKg
79zypaqUksCNo8txs7ZFYWECQV1qu66QWzjHZFuAKbXhGulU/WBk4L4PXaycfICR
qm2mTbHDu1m8RwwG3Eu66GZExKGGKnlZQUoCRbnvQmct0F4uGIZEeO02jjoqkhhQ
wW0obA/reMVB75iQwCg4zuTe5DN4yt4CVl65sepmoLqAPmy5dxsBQte7x74dyr+b
goTi4x0TUwIiTKgiuWumx7jAJKk538P8G8Ydp7BB5SpxpJlSzTOwb/eRT2u+ffv9
KTS8iMcPpoEGVOH/f/ePHrEw6lZD7vEnA8wiUsDPIMXg9Y600VpwTfIJR3sPPLLm
4NN6yPAVdafXWQVCoW8TDW8gy4DCUqZptX9NGoNbILpYSxXBqgfNs9OP49JDRzez
UuIdfnaJo+8zbkWr1I0YymJulHFMUAvPZ8OVp7zJPBMZl0IfRci1eJNFzQvq9UnS
csRbO5GHd8O+PaQ0DACGGj7WxdCL3wkQ7DOXQrLo99+yLRnwTobsU9ZjoklHPegm
bTg+3No/G8LYUpLaTExp+jP/9tWaYCiCwD4Swvlep3p0jyMpSLEzAyz6wn+gT3OV
8TWPZ/8FabEKgaaodMmVer1vFVr7lZePoRxHaFCJJ/mu5mZmkpQ7Sb3a4Y7qK+x6
dLU1L7AZ+tGEhct7nUtbu7YmaFjrwxeezZ6QM7y2/ee/jrLBToG/kCfm0c29E3u1
Cm+uoBFus5g8WhoxBFI081pUTUry2KuBmMJShkfH6nc2Gki21cxyOzJBDr9xSRch
Rpj/k99PbqxPjcGQe2wp0+zU80E53RP4xVBzuXqVBBls7/1qNSr1ZDaVK3II3zMV
sfT/3U6tezCAs5jKEL73ISwFSy0pnpjh8NGxv3Ic9bfYBn2O9x2Cr0cfabeystAu
s4z7sM08DNZ8wAkF0iw1Dgc9QOTDT9Ctmz2Z/WQ/Z8TNcv8BdFGWTkvmlSr6NrUT
HZfWzxC55E85+o/WTwCvv5/gJzgjtbL/TwFCeEYKhGA3S6or53oi+evyjxELyLwK
GGDjN0Fa6Vmqe/m8JEdfJxGiKFAsUcdlT8Tr3mqkVQDLo7DgC0+xhcwCyoyjPq9P
b2mx5HymZnU6NObzVrEcee7cg2T2VHVqSY8mkEA6xtmRNFrS8jdiUWtlGLDGQNcq
/5C72utWBCm9WbpUeVTgzAGH4vGpCsR3+KmWQw/ho6H8HFHy206NniYDFjdgmcTr
lmdpL+3FWwlju1WdZgBoCeWFhCdVq7stwU5bl6jc0mlAZ7bD0BKxHc0akeDm0K06
4bbTb4JVVX4+WpZY+Un1vn4xuUp3kzHEjHo1uzW2EdfcKsx4ywGR96OkOLP03BCR
1l5DJsBedGhphZWnEBwWv1D5+5xiv4IHoGqqK8sylP02+Cl1YsoRwXEgyxZATrNi
HVDOOUshZ/zDtMgnuMnnto0Kukm97kqS2WWTOdqPsFyXgJILCJOyAthAqhmiZ2nm
Mu9w/EfmC22zTudHhMvUBYajQhd+i9uPsGJdJ9OjJqOspPrZa9e9ih1QwbNK43yu
R4gubG10jtT4v0jcIP1iHinbQJFLFhDRhYcv4ty/g9M9ifXjar8lOkW5DSks5qpp
HmP7UItCGP24YKzirPlDKE6muJWoWs0Kt3V0783T2Nmyqc915qR4/W5S1BNiepiQ
CrG2twmPTP8yNZSY+qdMdr09QEBKn6X2BGncEJUbMOYJ2UAI0Qle7J5MICO4UL08
KAjg88VLqCO4DLxtlQftdl2d9V5bEi63NFF3+ZwwmziNO+0RK1t1cXPCDGyVy85C
sOaHAVDqpSOSCybDJothIe8XjLgZEerEHS2NjHKxmIexScyMJ+wHDqKxaeHTyZUX
cH/+6j1ni20hS8QZIT9W4iKk6z3mq5HsO2YOGFxqS/NLNEsZMurtFQQfGoNybnJ3
LFEOf2sDR74oO3vcTf+0F4UQh7ntBkyjUCAzFlKQP1+5R36ZoaON0w/ZpGckol38
Zc8hr+lvITwjty9dRuRNeOeDdzoEjyn3NATO3mJVRd9xkbUXQrLbFIRHVH6cD3AF
J6lehEBElxiygNbz2R9/DdgM7iS15+whtWpeR4Fv4qm+fHclCUiz3Yn4g4iY08AP
rL3JH9SriJTrHGZWosgfhVkPNd4FJY7FdvlMXmd4Xk/VzY8s2fswFkkKB/MDxAl0
MNpY3pY9S2l5E4Jz91FWWzI1e2j/HLTpULjCloDDWsrysP2Xu2T8gbDAghCx9yyr
4+KqpqggkzugrgVgoWPV68onIQZXdShPS7li05yhIfXFhF3PL3UzhCMldZ+t2hOU
AXSml0iTxTNkfIAjMlrX/WeBPH75Mvyd4IoI+RhjFMFpSYuzXX16DQkU3sQBjeiv
mM2RCG3+WFVm5aaEPJSpqxcJtfZ288AtSuEwverI5/vFRD4YpODxf/gPSPCS8UND
z9n6Hgl0EHc4Jl+P9U8U/9ymI1K1nDUcHvZsQt9ekoVvZEfaQ+V7xiCJIGv/U2g0
tlQqVe5wJVtsc2d/URZt0N6LRz0bd4ku6pAWXp/pStC3I1UPqu9COwPeBjxG5uFr
PJwokFYlpmKxgPdrE+G9H4XnT6Ms96nNlgI9f6E5n/DZ/U8xIF9KDKkE3x63nfH5
I1N5J5zHyHiAwHedF1h28hU0gwQCMBR7KxbaSUJCeBc/WfWF6m8lbSaK+JdW5oO6
HuJLoQ32mBuT99pIJnRXuobulIaMRJLW1QXn66yvZEzcd+WHyIYGKmBjvqfAD44l
hYyZ/rj149k3MTU7ECvuYPompWHBqHIC/iWPkm1D1/qPdm6MaUQws23nblPo6vFP
toerZpTCxVMMWhYMOfy7jyncqhH2u54/CClOjUSJiB/saNTkGClqjRnKJsGN11f2
s0rNBluz1o6k2vBwOBcobmtozhbAgMsXGaNTHifY/czDpxZJ8CSaixC06Oy6FQ+k
LHpIwxCrXdNTG6Xq+pukgEPN02QSwXADDotoyFwEyh1URInie5HndHSEm/UBdK/x
on3itpFea8AvpTGwyCbY7LlSAwwcn9rJhZ2LhGR4Wy5iMIIH8ZkR1gnv52IdMRpe
x5pauqbLD18KVGpeSaBE0Ucj8bx3AKrQ/fhH9TvmzG+4c6JQEalg9x9BJr1gF2gk
YIJDJq7hOi50NIFhInkl38YlbsKHedgdsq2SwDjNW7BzWub0jCfwk5uAOdQ73NUg
GxSyL0rst9w3CxTygqPU7KSs42RCWCl26wu7Y2UOseK3mxVpEzH0o9cdCTZSG1X3
fpvUKaQIH0avxm82ElmHtPCR/Op4EPUJFS4q816M6+UZdjUMJEdEz04rA0KGBdGW
BqK3K0qz82zYoyI61aAGuXCpSTp51NZn6ArU55b19sIX6SDZYqVDoAHwD5GGNk5i
tzc6pNENHjV/ngU3cjlAULST+jHCFhj5Z7e7+VoHvQBviwSQssylBPu84YlWdHny
Z3R5+lJRZp42RXP7Uq1q0iZmwM/AZoqLmEhLXMhLEkEqvjY03HyPZwTUL8w92C3y
eODN6bYAPllVB+Tzrfrpnh96bJ9hKMWmCHwRNkJ6OyARCRZV6RCLa3njIq7R169W
o8FaJkOdVMTumXoumgwIp6K12yIleYD0UwnhqV+4dRVoCj4LfXpm5ciU7nijmNIp
AcAftFg3kHiPJYqRokQksKyMfKbxHLCMJd+ww1lIesacFCOK+HcYdPuT42oHrbDu
ubRYPysCrWCCHaW39GKkwiZrYAoL/3fc7jVbZ6IKFECTTruuNaDbItHxGpa79bnp
w6zBA0DrkgTEnmG3g2bJvDCINdYem+FdIS3NiLqiZqH9w4O2jYfsXO9s0w83tM1V
gboAYoGGwocC9AUPUlVALXb7x+onmLUMCjGIBKPEBvt6Ddfk0CKJN7APYp46wWv8
11B/uCaThO+7tquMAX6nB/zpUpc2ILynzLwaTdbiHMnY8gbjJWPWUJpLJKyuALEB
MnpK8j+tLVq8dbMR36pOhOa4lxHNYITb0QnYf5Z1ch36h5HuJxKaCNWVOGCGIjRx
uDfpJXUomp4nLqL2fDLXeiu1bTV4yeCCYWTjwHdHuVMZry8oOMUCUJgZhJ9CH3CD
zXgNAwrksMzIEQm2Iab4aclKKbTsIgHkHQ2i2G3p+oGd69JmSZZ/EjiRMDORWQXo
vX28I9KTgTARmaaYvtDnEaUHdmhG7L+eCNIbfCgxKgd4uFTG6ezCVhEUZyYckoSb
l1DdrBCG1OpqbwkTIZEWWW5qjOgdqY6+17iiln0UfFpQpuQorN35xHgXftG04rTl
+UN8/DXlaLBJlXipeg5rMQrj9ip1GNpFaNKfDB9vuIPV0y9467PK69VcFwEtr+ux
tjTMhRkK/nDix15Y0z5P8aZ0ICHeWz2Vlvsms1psb25PrlvfZB6V0CWdG33KHsKZ
XfjY38C0fzORVROnvIJ6T9Y//oLg7SrYf45ZEzN1idFtwMrrABEjXaObW5clwppG
ibqJ/4H2LO9DcDMsyaFTkqLQmkJkmDkpEqwpFewnintSkUyA73DHYg7niL+Ox0DF
5BPtlNwVcPX3qW+TU6rHT4mxMNUtP2Bp8S4hCdSwi/ATUlzDvnHRTM+tzvONDF02
ND0atVbZtSBrSA07QDDr0QQg27hZGlH+blfUEnR+rCmVQHvJ2m7MAVUrMULFTH+5
5uWrOHnVInrjthSYzTKk9bqsJ5BJ4v8qpl6RqvUU6N9CN3komjoEWiJa3YZfDo7d
PYozDHrZy+PPLJ5JYus45eW0QOdzSD/+EAuyx7j34AO4/MRV3VEya9r1/1HGos+S
dqH2bC72w1pgWjyv3UVdRflVUFWo9BPS+rNcdup2UDF5wjSx4s3tZEgXTuEAJJMO
j/nik/fHTBu49a/TPhS/g/4hhtmYm2Ot/ij/ismJxZ3lcdhqO1sz2dZ6eUucKhmg
wl40sIaVopgKcT7kK86kIqbGJCAxcafmMHPhm7t7r9YTHLmyTuKTqDs4JNi4xXtH
exzwdF8PZtriuHvy9ZVFOgLdRDAXebTKPcvKw1wx6MFfrxhbgeSaRIzautu84ZuZ
kCpVWHkWzgu44gMe5x/Wrx+lMboPntgrJrhGL+ZisJe3cJXmpY0CZy6gdq0pWd2R
CJl2NKYHToRYE3/j4u+EDE6yRZ6eQ6x91lqNHkK4VJdz4BeSHumpr7wWqvOkZrZ2
nuukDI252xTU2DcyX20pkbOkLYNx4WFNAqkEUfiaIwdOMEH3Gy6yZ29NgZEvEXBH
kW4gEzTq5KHQ2buEfQnG9xhuk+qqvS46WgE/7W67GC5pSm5NVxkKT9pmOb5+ToaP
iZmVH3L8Yx1eOD8AurIdBxaR0dAkhA/IueqfuCPZ5rClYweUZk/NoDU2q1T+fTJD
RV2YwefljGX2R9ZEazIuB5eMQl57W5dFLnfjIghUlI+oQn/ajlY98cL1IMWRI1AW
m9QE0clRWcVLT/mUwzjNsEycLjP7QYlzpnRER8cyeqAk+kPN8u121DkcrP21FZZi
AtdSxZJwuBVOO6rWXwFreSz+cA4Ci9dhNCF+qgZFclNKIYbYOYv0rAUXmcgzUrIe
O+X/DgrBbNoIkng5bDle6tYMT+jxlACfHaaO4B2WjXBHov8+LStWcX9PBjcz/m2d
FEIzP9JOsyb+WUXzMesFflCgVZjjzYlYUeqd/fCqv3vCFThmGluyukC4Cd8zA83n
IlvtgxXRCIrFuQF4N/e2va4Ou6ByJf3USVks072rzmvzAzqBnEqRIKYF2NtaZGMd
v49+nD8bxMxnotwxWX5x7GazaxmCAdJE8Jt70/zY8ZovmfiTMaqXt7d1WNfKUsVq
KVC+9+5dR6z1S5PKZAKq3P4l7MTozRiIBNjehqrURa8Vo7c11U/+2sAXxgq1mNR9
m2c7vl2fsr6Hse5axDMgjIwZCChg9LEBkGTYZKukOlNYpofkE5p2LbHhhdk64/5P
iOazfDHLya84zjmHHJbQrupb+1Dbj9WXGRgLS1/p2r6rgYQo1ve7eapRUecpO4jm
/235Id40zVMGM4x3c8pU2dj6qyec+g1BKktT0KQQBbSZBPPyhzQntk/SHb3Hvb9S
L63E0Psb6+etqSC3nKlcUaac9Sg1ypkb+1/nEal/rU7fZwdeFDt4ISp/lqoTnG1s
1I0UvsOikoFiZuAKdrxjghb/4u2Ux39kEucCzjOO3y3yqcJw06zCXZU74g6cAyNz
8/X30R7YN8uEi1yiXrEriLSp4E0YRiKEbzm9Tn9SvBNim8UmINyW5osGlyn+2M8e
8J0qVMI0/ly4I8Sw2FANos9NaKNPJCuYuXhgRIW/uik=
`pragma protect end_protected
