`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
p8mZpIA60zDuRaqNWNtAD83lMDV+9+fKgwVto5W9Z6BKNwrsCSL+ykvWd7pODVQZ
MNi+iKNujlv0d381A2PYVRhWf57lXGjgS8pjoa8fb2bbWNGNS7JO9EHTpo4Gqq2s
UV45r+AhB/49FqA0sB90WZswmfoptAjlQnVSr5eGQ20=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5632)
Odmj38d273Wm5JYVJvEmewcl78b6GCNpLT5DV+td7yudRtKisnOoiVSNn0HY7/vz
Caw43mto74cbqzZhB80HhVuZnnqgWH9213zkbDjdEXjnHtflNY0AhVpR/O8Wxnr/
7DUm5OyJ0g2/tnuY8XcLFP8VVE3kchTbdvGX1/FVe1bduHsZVjjcfzzL0o6R+aFT
YPhxgeOevFurVpXvXytaaF3ilvYtINExPT8iqnut89nBoWQU+5OaDSkttRdOQ7DD
8II0Ly153mytg1fdg891wi/R23VsMMgJGGVdm9V9OQ6+zqyXTRdCZ1jHhTDaFoz9
hRzuba0okrPjmC/0maWOXfjJB7375x19DhTiV+gps32A10gR9pjuw9AwkW62+gUG
0czoMJfKc5sMwIal9i2ZOWSwpmpiVBWZ3jolYTpxxn2gQlBVw1uNz2pjf+Y2XPs+
fkLnxdLvtmnOWu+3qMb6i3H2oubbyCMJw1+blpciRYuO8hTpGiRpp6GNNDChl5tn
4vp1sdBtw0n0bRz9y/2byYlXhz8EdOxNJuyZJLzPBaozw6wGhQHCeOcOhdO0RMs7
xg7T7BZ3byjB7j4hcYT1Ae3LQmNEKkvXZaceMjowhZWqcVxR+As4GGsxztISaE/Z
pXFBIfw1fX8otfCtp5FbMnJH5jwNlaHImfm/97rGFVqifzxaOdVv4vhlVj179cKY
h8VG+sltJMpuEdXY5VRNBSK/KuV9wfIX5uIwuRNZS5GzTgXVph591EdBnEBkX5Ty
5Scr5i8MebJMvvz+FrjYJDGBTIUORYtzbXcTJusHmOkZkqpT95B0HM+FILIjW8Ki
m7e1XpKAaZTSLLoQWwsNCtR0lQOoDtfWg48GU32gB8/9eEz6d7wlyE5eAnSqIFZA
ODwhQHsKomCyzCvGOEeJYn7yBnY9/f4Ov4aRGADMUjEW0B/+NxXizZYEUoq9aPvn
EcNzu753x9Vd7BAMnWfK3tX8b6HTkaC0IILLr9DqW3aWJgnWIrlRR4/ZluHnkQr+
fNX8C/l9U7kAoRGA6qfDRUBD2l78h1NLujDra4J03cYJFeiX9XmudXc5sZoOLttQ
jMW6o22+W1uHDOGsNlRaaSO4xvgPwfUJIvd4PmmdnGL0bgUtTnVzMwpd4pVvKYdz
I0dzGLuXzc6mgSbndvKm2muxussUsOZ/oFWVNDPZ+4RUwzYJsFYuH57NptfhGMRG
ijy7BZbuORmiQTUXD1VZ0z3G4nc3gbbXaFHQ3nj/zswEdl38P3Pz471+DdRI9IQw
ijT2g5bHyRRcNGQFz4QZ42BJ/NpDSgCC9lGwMEsy0jNy0tV43oaqI2vCJO68wmNv
RoNLmp+uJOxjKY1Mf/AG7yBxJ/4dbkIix+8iI4a4XUGV++G1E+AZolfhdGXkv8W2
sgmaNf6vDCL2nX5NibcGtPznAxOSoIdCdqYip8lVsnlIvu8bepIu/ZHf//jUhbEI
fffNEDMuDD+ec1EvGDMVi+Q2gTm6OaS5i6FFygeN6ZinLbSgqlqM/mUrGMAZWEA0
NPuts/o6U43KpBx7Da1Q1goTg9d+WXA/D0IL4M/ywtMBJrcwABhcPehSYbBr9ioI
UPWJKlYsmPLROmRoS4+CxqXk/0JXSa3QQ5/wJvRscIHdj+VS0x5KcbC8vclahYk2
KMhOkgUfuJkB4wu3vqYU0Mke4iP9knM19Xg0a/SJa8VWYzdGb6VNxxckqAZCM0Nv
AtcokssMPCvELX6zb/9y5jIAMhemEsf5fbHujb/EijFCnmq+0HUIJzmqIjWQrDdL
OFgm6PtFLJUhDO8PhUzsTHLWdB8G0kURd32qYc1RuKA6pIRjMJ/xE4T/EBHBsG/N
It3N2wSxsz7MG+v/EzKS/9E3xkfgSOgXny9FZc/RmHmk3pUzBMJO22aA63cQgq5p
CHOsEvBlTt9oBoYRUEXKGhL7QoFtmABn1F3EmWxTvm3YZ5bnBWCcnUdykeU3k6xz
2y5N4EmDKOo3nufLHBuUJEjMNfS/Npc1Tr1SEB47DhclUjYMwXHguYs4CQdM2W75
wRzwORx2DFTI/Ma8sLmnny+cC46y8cMLPAw2sa4QnxdDDNxnEup57kE8cIK+8T51
zpCd6Lm8uuJ7bHyWySfgs0wcELAqAxLvoIee5lRzrXzjmXWsRLSC2zGsGbBIGCEg
fWJ5bVdkqmurFnAgD95vTNNSgBF77jIhoXO9EaxjRnZEdSu3q39JT1ZfTgQYLcuk
boYmdqK5BvD55dCHIKrRr+YFtkK73EWX+TBIR3tFy5Tmp6b42JjZJOnPEhZMdqVo
rZ4k1nSHZKCXwACAFaznCZAHotrIjXNaC+hnzeh5BSuNz0fjF0ccliYn9d56Rx2L
AR003HLYeoiz6geGQ28gIVbxgxpN/cIby+fk7zb/QyuJsrP56qqZu2q+pCzo88aA
29Q7rOTUvgb0KPvA2YTI/sP7UTQZYcOYW+6N+mon6tRCXzPVSpflNojFI3KsPVNk
7nxPbos7KtTCDh9/zZx8HErouLF5WPS9ejNF/0h6/pxrbnLeaKD/xnf0j4JVbRr3
f34CE2GwprhDXrFwQmbw3TAgJ/eNM+LSByM6/KGLqzF0s08jw5RyUtV5slvtsd2/
2i1lbVvoYHOBhen/palkXdEtRqP2FgqpwSzTk9yLefhiobBQiW1jpKrg48MD7dD5
dCtumROOZ5U7lP7wf2LELSQMEJoV0o5g/yB7hMqTfVAsNuhNqM4tdlABKnrHVp5n
r2XJGKow5LkDRYEi1q2m9MPfhmmOfmbH049907ozOHS89+fPtQ2eVhzDOi2GW8se
Uox6PSeI7wTKJ+kX4zJZB/YexmDEg2f9nUyKD4UxWVaDqmYxRM3DSeL+8H9P/OP7
kXzsSP0QDaYyij9kzbP5p5npGlHv/yOsjPnqRsdoIcSvWFgwIFZXgu9sdZmnTbUq
WONfJczmjfDdS5bi2rJ8V+bnEj39CEs7Y5iWF17KlwkWzYdG/hYzNpFtlEwU+9Jg
H6acTtsK5Try095YGgvjkwa34zxq5eL6RbExphoytx8sYSNB7DfjnYqICAI6X+nB
aPLhYrp0RX+MEiVbuAFf9Qb7bKTxj84Dx1/S55Jns8NlqIWnTtMYZUNygjjB+nYj
iUZBoHi8a/4748sWWKggpJHkcb8SMrAHn2cgNnWoPn+nbVeOOgcv088vXgGJAdu5
84vcivXwS08sfNExtmCIrs6gUtWcFlKFrrQE+YtBzo+qdIDYB61BKVtltZiJYIR2
U/Bq/J5JriVzTy0AnqJv7FGOF8f36/hbwrAqIpShRqic693GalYak2cZ5R8+P9Hd
IHoWfTa0bz730cXEkXrbTm7mgH3fLoc6aJyud0lM1nTHS8r0yk3yUQj4NXXGjtiv
TJmGoCDi0d8s+uqWutl073N8aVaV+YLvUM/zWTZtXN88Uzn5LtQOUfMT7t+NpBME
vIzdjoVkEPrnzYU62nKx+myhm6iBAiMCSz2genXtkE07I64ryvj16eTMrODjKkDE
biRJrVa+Cp44AaiPMhs3TLtqddCUfJue8UjR8wHzgylahOn8L3xsetxJ2Wr58zaX
FzvMA3Hb+zNxgJu12gaRcqgKGuVHuCX/6H/vkEzHpRT/tZYq+kqMNIHM//uosAsM
i47PUOebaP+heoll01kRTFL9hbcZbfVCbyYTa8vYwXDGPgeVNalXndWkiaCtYdrD
rXyaKfn/d5j/VyvXuyyC3F8YIELcCg+W2vSP8y5ndDP5A2jI7a1MjPsZmhi6cnKz
Fr2rJNm1L+Kjr8Y8sq6nXPYYPFhXUfr3DoMzMGzngRZLRkNJi9Ezwweal0PzX28z
kIakYt+aKejcDXbKGUX9dYceLnXSi4ylmVUTk8kQP2kF/+JpnbS4oFN2j0Fp1TwQ
eZTpwreW6qzk+/+H0O4DqeAFV3+1Cop6hmYxRzI8E9hb5mJf5a5uvO6JBWj6lHfU
8DfSPwJrhvc6URjTf83yKJYaDlAgAmesgEqLbMLY4Z/khEKbNJF2svs+LGy9vBzV
9T5JgnEhDAxlCfnZaTjXlFK0O4qK6tz60i0J/pQU0+gyeWqjn9ByftEruN8n3ZL/
pO4vA5x+GXF7I4I6tL8phY1u+pBYrY2IopROYdf/4W1RE4GJUYpmUBEFifW2KWiH
/2rQhtQyaViPPgZyFccwlU131aTWf2vE68xptRpilgj8Tkt4CbBE/wolj+Dbf/Ng
tvqwk96HHzOw5yYzIEA1SNitUFKaUCL9lDrItR3TQ2JzhCwqCq0do4x7lkohxhk/
V/F5xxY6x6gtI0r7DKyzl7DjrwgBdxpuicKBlfGutVf2KxcoNI7TPM06M9kQzZgs
n/UoTPI8+Al6hlUq14PAzxO+uZQPtapHRIQET48D6Ch7Havib03yzitixxFRaat4
OhPs4nL22qjON1AnYGaawE1AuU6aclMiRyR9dX8KkOZSFzKrC4F/Mv1DgGaYyYvW
AuCZXFeqRLCKZQst061V6zchh4amUO5ociJrMNtHzi6J3n8vqB+dn7+WUC1fGWG9
4pcbKcOf0I7a8f3dkV3jBCKAZ8JZWWj/vvEL71Oeu3VgHFdbaXfbaljylzA1ArwI
PcNxCD01znmaBoBcq/coZjQg4okBld0Nv/Ph24iY0Xx4P0aBDSxqI5LnFLEjLbb4
v3euHMhYqp9EL6sECBc9AFNIJT0hPAHNsjw2dzQUs9YzK7r5t5HUEPo6MQ07/CoP
GKH63BwhRLJc/Qs0GnrIh3FMPjbDtzzyVJGoUI+6ntCLU/owUx77TOb7Nw0zagRr
pKHPnoM/VHmYaPEEU/bLN5a090Or4zgIXNS129+vZLW6FF3UOdz/5DmptDpgPxQ/
06io4Jj5v/Pq+9R7PDVaFp3+w5GWD99eZA0g9qswGsymyjeTJMqGefdyPthrN279
OcGwfh/HnTQ/6ZT/xJ86WZ+W3W6Uv8SEdc7jQxVikJjw7wyJrnWaumxTDt8XYbJL
e2nMgU+9inU2NBrTpjTd3fFl8hMbmS27+sGRbNJ3uerFFl9WpqNP4ddYaP5V8LyG
GnEdBEWRcA0AJ6GOTuJOPZmt+4bOm7WBlkCR5tD7c93BAEIEgU/TUaLBdLNP/6Bo
JVgWbXgy5oBuGdbfj8wO8UvqEqqDWv7iwdR9S0I9YNNZ+zO0GIbdP3vljcee2r4N
mga3hBFXnKQi8LG49QO4qovpLENlR7rOn4AbcS9IjSPa6D7NZhyRRKWUn9B3eqMZ
4OUsrf2PXXCDYhzjEgwT4WRJTnSzylqaHwpj+LB06Wd/3cuK+rY5Vjvg5wnDAi/p
SlceWLI35DJU8PVozzN0qYIww2QMN9U8Xq6i8/Rxl9WyfAOswdfZWU3WgUpM16Rs
aoR5pNuCDqsM20A2q7zB02l0cqZLlyZCP19uH3XDSdHrpkZ8zqZn1y7K48jU2rVT
IBExSGY7p89ESh8e4K4k63+is3/GyvTYC47e+FbgR0aVe9V1FXi/FVgiQqr2QWQs
nRYkX3NVtfXpk/5K2XlWg/6JxLvOUAojFFvKAx0vmZHggHdk/43KJ2mN9iuj4y2+
/Za3Em/SoeyF4INBKEiuatlXRFdRXCLlj/Ft0AlziZbXR2JFbe25wqEZrBMaP32d
t+ot5okKCZgaM/wTHOBqCzKlUqdrR/NdxRuyyiTG9UV9WIxDUcAp2jaFH69x9FRM
RMHczbG5Mw2kzwg3QYvgxbj6MhX0jyg0mmEo6vA7IghNJu5w0acLE4McS5fWWNqx
fpy0Ymdrk5/BdVaEKs/aFpWJZJ6r2LLSXpR+GqLyaqSJTyy52OkXiCY9uU0je5k1
0XZPNGlbEkQRhE7QzzzvHvJW7psnyHxmViSFO96UKn3iz+StwDOIRtbGy9G3utZF
mEg9lmlIAC2QV1JBG8I+RxgojJAdFbxZ0CKsHJoCUvn4IV1aFzEuBKp/g+Ox3hSu
PDo3Iz1upTEQ9RoyOyGZ8W5SUDWngG8fUJ5or+2v4qovRjZ8lIar6ZJHSmxODr+T
q2eUxhmqitMAR50fyupgWCArwMAfDUTM7aEf8V2Di515O/XWVjFvyHHMNOA6cLuj
CJzxSWQWunuaK0mkF3P7/BmJcyhEswDV6ZgoTPStuytIT7YPKoFYassp56wt++4a
MtkCQyppmg3A1Mz7T9q19e4bZk5e75aHzqEjymDNwGdajG86JcYcjzsN2aTmBbg0
vOBF6pZeLPtYwVvYhBoM3tx9U0N52roi4oDmsJAHeEIhmlpAib609gxNuq22068z
ItUg699+WaXVVSASSWrKMa2ZDjvEl6V3TQiMxD4fo2AQR6dg+eO29q6Omqb5w72p
jdOHo42ErQAl2QidHXiKaHE7/yuyPhdY95IOXpPxgxFd7BNr1EaFUtE+0Jdnuszn
seN3Pr4kRstjZLK5nTQ0FLusD6uEouIcOtFkin4ahU7fibS7qupCmbcd69GCE05L
q/BLKfCkbGEaBsrVPVJCZWe2sfUvo1MqDNf+K/ghjvX6jYiVkvyhLaLx17Z3aZzV
rC3Q2j0/Ne6TbqscaH3PT/zA+AKvFlfoMRqPjBR0MGV2JnuTNGur9tJL0X/E+MHD
ulXziddUd0tM8D0vsEsaeqtwh18WzFmCpawRUrNN3Mg/0nJqW8YcsNRe0NO8ygGv
QWb8H2egr/Z7IGEj45Dpmd426a/LlFejsot8es2j7PjmrKiwEkLNM57pw9TwQuY+
BYSgXpU3GpZjrlQ4PVs9JxxyWpaxMx206D9aNxlJdpizEuKgsKnVCzKWg2xx51VM
4vWcu3hWlcViTA0Mn+7EZdDdVesC/TfO5p5DRo7NAgOfeEDFzbMCJozPTGO1cFFO
4lWcrN75HuCCGbTU26ixVXS9f/vAE7aGcPWeE6/B4a4uSiH8/uU6JY1qZfM2SICH
N3WnZ0Yl2AQUn7dftmmtelSbnZHuLTtarvacwdxKGUTOundG0GAxZIC4i81Y9AKm
WBHwrNOXiRsflVx/qgkMFGj82/OjBAHUrCMqmeayHBLy/QlR7X3Ga84BfOAAoCF/
XI5MeKqOBymqZ+/seSWffW1OeK8DMpShuDL36ZSbIozt4A0OKfB8be9MxtmcZm+s
R+LVXc5C3x6sJGuALst6LBdzO8wXoMklRsiusC2R+uFtvwOl7M+YFa9ZgOX5fEqO
6Uqe24RwxfJoeppx11/xYbPhirm8XfEqPfFkQVxEe300mGkx4YDQ70z08FVan/mh
zhW7+k5WT6V2wc3JXPrMQUB1AN0XHGTL05/3MPGaNiNftYhLNmfzvw54OOouDusl
Sk+PWNy/VHRfasrjuj9hIspYQzooVev7UdopfkpE8oGhNf64CuFR2ho7gJK9B7uR
lt9Lt1qDI//nai/ssMHVUV9wCU2267KCXdb+BlFdzn9XnID/bVcKOifZM4Mkjn3J
OAcm6f8zMGHLpwCHdQnASedKKJ4WphBEaIEssdjxY5OV/VXqd0DMW6roGqMioCy+
6BxSJqM3pT8UCgtvPtQbVQ==
`pragma protect end_protected
