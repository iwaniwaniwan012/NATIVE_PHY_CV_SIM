`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CaDxNJrLgTvi3pZiGfj9lCANoGq5AJgoLm/YpKzV1jCGFU3GIqREUaE+q73EmnML
YznnokD82uCjTmlT+IcdwqkgedN5hqCnuiwSAsyuE4u3O3rEE6dq1WLRMuRTdP2L
NhiyyRkQmBdVUcn9cckBLfGIJesEbgvTJV21WrzgUsc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 70000)
mjtBC2/V7Or25wuku6XC7475mdpAy65U5aluSMaclfPDxs9R4hUde53jTUk7keBW
PHDLKvf9g8aVobgxU/sK7yvYcMnJcBtP2oSPRgMpqYgREY9wKMIlBqLBTRNxEbXz
nZZVOPlo7DUMNugCMzn4A11RsmQeYO/MUeBvBatHmWRm/tkpWq1wtCxUmDUQROKK
hJsbf0J/FLmkPIHECa+CHOr7HDOvT5BkgXtIB3krluxLytgNsfssPb4fHMGgxhHM
oeGkCWnGM06b0m40+boFf5zB6CaGX0tWyHF9D6AszU5e10wcBZGkf/8MIcjMAJJx
HHljwfRmFlo0LcEUhedP616brlcOyzD/3sFDqgj3QoAbwlhwU/D7TY6RiwFV/Jwn
RDJ4LSjSmFwTQ+dimetZscWClGdR5lY6Q4U8LXfu4hGdRb0Aci66oEr/AODKAdVz
WrbJnCz+9REombeYQwdi8joKeqSf0apYw6MhmD1f8KBwKELYm5K0rEd/hydo1vJZ
B0J0ZvLahhv2F9liqZ1oFcrWLbl+lpz+8ect1uecILdJfnkqT3hgbuPdV0uAL6At
oN8DJNzV/jnGMGRuWLnvCSzH0HYgbHO5VuRrP7EU3kbzJeNfik0gVYrhiswdTmNN
WrrX7i9C7vwcQu7JkX+PD0WHBemieA37JASrulNoknvm8xlE0LrYekyOnR9NMbiO
WeR9WWG6foOoO645f09uVzkyK9QZAlYIZbjpujSlRFJbXoKGlIWQwY4B4JEDHJgn
Xp7W2qa9HvPUif7faBfSDDsE4zVTM5YcvECBq+Be+Z5gp1Y/PSTYkaLYNzzORMBk
tfBARl5rx9kJH+MkBkfMd9QQiXoDkXoFv8QPdOnZ4qsrmcUVoqBeV66aruG5VIud
nLNMR9nZMdg3SkgOqXX6wbuH5Bosmh53thsR8EnU7+1QFg/HLR74VcG8ibpKTAHe
X6wir2OPP5ZzespHacztzSdFUv6YULQiYI6BGpUNPhsc7mzr+ifJ2fT+0mWZimZ+
JbyxdZtW2wR7BH6nSrwjWtqw6tjs/rRrWNrwNRWjdGGeON38O22s67ZX5TEwXRY3
PcpVPHoePwnw1GLg8+YZTwIBPDvANrcgQ7LG2I0SHx78dXOBGzP27vUQDcQrCq0F
EHQXIyOr+C6O7/X/AZ9ONR2gao/MhHFfQZRp+OK85Uo5/7XwVGdHiG1orAmu90s/
jpMkK0A+mp1Fya1Y4tI10cAMwSud8Q2lRscHM8mrOn1v80QF9i46nTub6RGmQcDJ
Gk6jWWADuaIZnhwNzgfy3+oilJv6PhRY3A/NIA7nJTLiladiTa3hV5WcmobnAp7O
NeGfyxj/sSZrvh+dDJOz7SGnFp/EWklfOBmoeUcZZ3rCM9x1ekatnDVTJX5e4oWO
rlDljxpTUWaRzPbhXr2TA+TeoN07qIWEotEY4CIMWDsFqxUBAMh9yAulA+oqaVJN
0D9Zkq/bmqipj7fQ7OgZbjqQk4Wqb8rVvon4AiXTymOK3Df13INqKSkJ6BEC2j3Z
8TmRJ3S7RwCXbZG4oPfPYMry8CvPy4BbqSZvzzBt/mE7bcct6JF7P5TGXf4lBz30
c8QQX1c+ZejLgafksP2JfjHUYwgw2KvyUjUKQSnCekatg8Uv9MwXYahfiE6zAUQe
9XvuQde1qYA48UaZkqDW1aE98uDj67mqxdz4vE021ZC5JS5hseRbFi+Plq5Z9K/C
TIxV614w/H2k7eiawV0vxxjWCEeyKXXWiYWEWGRga77fTtltgAJLKpmY0jr3hkaK
4o+M0K6L0FenKWs2/Seluy0zR2Xr2MkHSbZLRl0ClsrRXe7OrLTbYpq3AAPfp89w
De0vqcZU+CBofsyHpD9zwfbWtrog/ecahcjdfsRNyRftrTiLtnDTZXylvbsRQnBS
ZvJEzQHGgpoPlSO7Jj4EjjBYCqMgcRn8QL0hRZO0ZKRYI/JYezda7Nq7NcqurH5V
wGR0Hv1bh8aDniaT4Xz44I87ZpepBn1F8+NqOzL0IaTtZupoiM6oh8i9PL30Xi3K
IV+ugGfqLACfrEGYcSrbwTPa/n4TjaE6xvGjyakQ3PokPfwVbvTdKNKMANCorqpI
9Rj1Ytl4XXCrepI8Cd0CCTLlgF2R0SKPlfNjjW3i7BFTHn/ZMH7fuRGlQo/ZTRnb
BtMPOPnfc2TPYCE4P4yH4zH7J+NyDncK3LFaUfYehgy5uHqo7u0fIumL1e+mci1L
rgdnAkzAAnsJp38FVi3WYXAJWseYYxwhxI6EDG1PMReRtlvhto/3jfrEq+1c5Jkv
vQsNwkWTs9W4GKabKMpSda2tC82XvoZxWGonHnNxXYJtTgNWM9vR4QL95AqNeSEM
paOdbwZ3102FEQe7YjeYrg4dBHOMX6UcrLNjm7XllaVfUTMi1wuWbWpa3LnfQt7o
dIpzILiPz0+d0Gz/i/moEdWIrCRrX0Y/HgSiXhi4GqIqftL1j5VXhQUwiXRAFK1D
XNTdlTL59chD0xnKee85XZs3Y8zjjofKJeuicekH4oSCgCFbJWI6epn+cqkPctMe
NR8aOymK1+MjW5xAEScYH5HhGLWa6NUVTfHLfi0kL1WAoR5jZb9tFPqFrOBIv6pL
nIQI6rYDTBi/OXGFHFUQQ8wXCus29q3nSNoHWFMW0BqOCE3og9CUhQ2T3kkW4m4a
IExhIMWzttZxp/XNgyjK+5MZLMFHtZHTqD5CJ1vhGILR29EiCysX465dJpDxwc6m
BZfXU2pUFmJT3GmbD7etumwxHVHiHe2aoOZopKKJQ+oYticq0m7/Hk+vDixN4iF5
HBUtMb0kK6NJhI/tY6FB0Sw+slu9b6LAa/PInptMmzmKkkatT271esA0J5DYG0TE
T4tS4rOWF9MoWk95gHm8iSD3Lw4G6DwoTVErSR7ptjuCXpB7BpD2TQsrv7NU/BAZ
dzOvlc0PtLFFbwRXsDOk2YlPTpfyenSPZbR20a7LyR2S9Z9S8Vx4w59H1m0stzZO
/thBS7qwk1Z5h8XXF/wOvZhbGDur9wt+6MdNKpU+UjP+Fs4EZSRlC+SQ8t06OS9N
GDx4EWHTNWwPqbJsu1LTbO098SzvW4qWFIWxmeP6UFezN05KXAdM8XNXVuuz+OAV
QDqMQLFuQiapwAgjWEsqrPWWGfK31J5P051QEWjoA+2cHE3Wn5N5/zI5iUS13oB5
YFfZVd438VdI/cz58e53ur/Cx/A/Bkk7Y2MTTmG4/OJIRcSF3ejokTa7K6xPrt4F
IVtXcdY1+kEjc9jYCpisPT2HIwwFzsDT05qs85bmkgpYY6AEKbudnEI8BK/VbbIO
paZzKvyMu68VWfJ7KxDAjGnuYcqyUjP9z2XtfrRYpC6tZNcguFIgonZMuPdypP3T
yWuDO66latSfwUsuzhaHNTtVQFrgXSzxdaQIAaMCsJpaeo5iClJ6KMLC+/GNoBc+
KOtZEroCdriiJzGexwqTJp2aZeLREs+FhaAoMJwwTrHBW7GIVWYYjFwWiPUAJnV8
OstOzi2cYWi5ZDmIL1JiiA4hqH8IuD8u7S37uh5Gr4qz4anPkxRKK+VaHAy8pkjK
MHFXeZAYvnctEdvMDrpEGjDQvegeJ65S9A0pqb73leLODThx1NwajRCKXG1q8JQg
2B2wYiMd7hIzIMX7sqOtIM6arV6XWvrXcegBzFUhNXvPnwT87oTCOeSrA9hFYprw
0dEIHsKAJIvFbeKCzXrapC8A4/oj75xPe1n9NxRTQVG1M/csjOkYiUF9kX7dmGS7
OYe1NLysdT5PnQnSF2J0Y051WRnfGvHW4dIVY/SAa6se0Ei7xw35KmIjxUiCdo9o
qyPK5L9pB7uFsWQElBLj2JWuw4q+I3UOiFwDqZ1G3BzkjFs1QqE24M5twzbVsiq/
w5fkgdZKFzOHRXeqT/qwpeyhB7a0Dh+ubQthdtNSQs9y97cA+gl9zMWj7gdlgEOv
ilBhl+99Wb/i5OsBwc92+D3tjpb3Qfo4PJwkJC7T6ovqht13Ruj8tXdxhU8C8e/+
JXl5K0RvI/9FPWNtzfPHqKYOeNrhAFqtTrIkolyYTocmjUBr2IsW3hMN2Ht2caIs
BXmqGpx1XzJUXmmYGWyMUJNOFcDturSYTgvFR9bOfDHkmdK/NyBaARxBHP1VCa4w
qeWrHSIIwcTwwDYAR3C4a+F5jBi6TiGi61HgXzBFbA6r9U6BSgC/I4D5uy0eaql9
XEO3JRQtxTM6EAmY5x7P7b7ig/IWFMa65w/bfGydoLcaRzUPJRyuLpF42Ea7HEYb
AjDgl5u6aSkC5+DjmHlMLQMXqMzxSSmm4D00YyhNoxNRvufEhgwHBg2msgS7Dp0h
mk5cdEacKzc2pXWDf06xYf+PZhbgOmJe8iCssmu3sELCGeRcoaKkZCwesRy1B9JC
sgFiSJUc5Nanuwt8FisuYcLF0vJppXv7YNiWtuYU8l3ACOzIndwdLJsthz0kZYlL
Gphjd0hdLuSnMaIwo5KiH2y2LRyNmpUIiIuxSUe+UMlUsVe8rnXo0K5WU2IWjlud
5cyWr69vQy6okyitZr8PBp4GazA7LxyxwNX3Hrxbsj9sMeb+1UAZYtR/SiFdBR5v
StFYOrVev2eXiD73fmMjcyQ0B4Se0k8s2T4xQRWcRiIqNJI49Qai2D9cYFhVfZVe
UMN1ybsWACKj6jXGh+d7OqDgiRY6j5/CDq4RgbVghZfQd8+UfNk8EcL8s73IRRaL
9OTjuxh8LsR18P6qsOOtORd3Z5s3eSvzxawjPm1MeZQ0735iJ8oeaYl0hIPmsZU/
dSt95mEjIzSshN42hPgHCahirMtwmxzevXd/ONbg1hLtbmQXRK1H8MkIJbEKbGJX
RjqNG8NIfCD+XCYT460c0zsmaO6+4IYVOo+sAsJLuOXie540fVWjfK9YkbD4v2Fa
EjGtLLKKFrnFM92biyrqRiQ1Pl3EHMeNkddoDzm/ne7rSnaP7Nsw+7OdhvQqCQdB
jw/BIXnhGTA9SVDcn7cfuL5uxmV+XkCUyKHBh7GzA8zDRj0+olojQxvdPuUOJCwR
1k5oJ8RsLewHoLOiy+Sgt0H7Q70810wb3W+zAy+lmr649uFDDIkcH9hJwKfcdd9E
Vv3VOYU5+1R37zaoZ8ClnIPe0BoEO8754vA5DdDiRaxTF9yBp8EfT+fK7F1KNC/m
9ebjRdG8e5jMm+KmFF0BbIt4r7Xb4EB7IaylBepNxVw3h/vNdlCOQ+rtZa7DHjI6
MF4n7gfT2RxUPlA6fWehTL44sa7RshF0z9AFx2Hs1VjOZJA6NLO1JKyUyd6f7JGU
pSHTIP7KUbhxqWGN/1efabj5R01ZacIvo6FE6S34pwBUJ5DnkQSPvnxquGABcADO
Gam8fR8nRbUOCLgEzHKZ0TWtc2FiA/emb1ry8V469kKg2KlxY++M0vob5av4MYZ7
M1hy6+RF2TbpbhW5r1ETkaRUlKNxgP95ZBT/F+MkJIWaqXz+pE9g3EcTzQtuiibF
E/Pzy00uAfq2F1DZLvHU0CPSB7AmAQWWZcs0Q9ZTc/36YpN4+tCBk3YDR9nQrZpk
G3i8jmeNa5wWZwp59q24n7/xRFA4Blbol+ODPseiuGPn4lfxEIDWQtMvM8IdbaQn
n4jJMc3IYxHtIGa1Llwa7Uk8fxFEmG0OpVCtR2aFdDKGAKGJ6xT0JKHGxgKX5ceO
x6VTsD535bt1u8zcM4M9FyzaTko8S0Vc2S2A5MSBBFTIldJlofh84HhZzTTaYuKc
JhcE5cZ2fvzRZgcrefWaaHXEa/N++emOUn/8irE0SGmAk7uU2a1DOBV7+ryR7PqT
jL50ircerguyl/ig/EvGOwNJmZ8wVwmxZZuZgTDCB86Odyz7uk9inmaYFK4DxdAE
srdJCm1nPrf9rud2/axKP9x1bGp8I0d5yg1cbVKwkmfXqwY5Jp6afp+119y21u2J
+iRxMPUc2XTb+JK3Y1v7kRrFN5ap82yRw4FYCdX1ivVPtZcU1bu999ktMJxOvP79
/Dexg7QBj0iUh/kMChSih54e3HVBknob9U2eqckQAEtmmhouB2bZ2U31IqL+qS0d
Q+pZO6yNNreDE+ZLW9biPEZOqaka1srljfkLFXpSnPvbXbjwtZygM3F5cXujvDvf
BuQnzPY1kAP3EVuSpx6Ooq3gHsd4QunoGPMkljKquq2foNux5OzVXDIwxVflI8GT
eOJJp2Rlh4L4UKZmzj/csHbnnjeMgSiv80drLjJyMXARBpWIeHCyg2DZVnFjWxa+
8YcFXaGSBMYmCpUoZIZzBmTZ/F3xWVpPTzdq1PkXsba7xI8K0upubHxMbm7sqCjI
DJN1Vd6gNNPzgpvoupy9EZMSXlygQt4zyt3EyyBdfLh6GS6/aXELxIPz7biCjjxd
/zf2JbGbu9Tdz1ekGlMpKHAF3NLa5/ya9e/tKuH93bvptSMB0QHdYH6OnILKPVUR
SjNaKkEwaAtAfANQh3u9NAsPeBm2HNnLpqOHdYBYxm63q2L2jPJRJCOOw2oZXr4h
eVa/iUXUS2bY65m2SAtUPS5ljl2NfQXgKrlUYDlf/zE1WFEpB0JxMF8uD0W9p+9y
n/2/CidozDzHxQ5H0LT9x9TWSyBFy9N5Ch5Bx5Tw61/JWufxIsIYqQOpegQ6pZ/V
UZhkiwPdPM4Ouq69aLtK5KwympAPT3W4U3/X5fYIXnusj07GlbEZobPkI7M16AVo
4S58AaG4JUihUH+bT7C0K14kP6ryQXqP1wnCzrOOthgn2HdjJWEeVhZsyEgnjqm6
qFqd1YFKE1Br8IsF0ElYbA2PAvHw8pHVl1ayAFr+57UA1LC2KG4ykto8L+qZ/bI1
cBVhGkjCL90l5gWCUbX3ZaPRGpps3HaXJF5KSntfUaCNxCQIT1eseAV6JDnywCcz
a+glgfztChb+WJXrVqJsfdXol97AEVNsB8zBcD2UP1650U4wGaQDVPu9OhA4CRdw
hIen0DRZe1sP6EbNCa9nMqGoz49ng7FlLDzXc4FGHs9i9sIlXCJ932uVyoyE5FUN
dDMd82HJmUPfRhZ45Iq9c5O0Y3E3anvF1W76rlP5FnbVQugAUp3dJ+vh43kVkDwG
u+MbOzcK5+PeWMiDGxwkOvSR+RVQUwvft7sRYydrQOeP1knacNLjbt8ns69AYlUY
H+z3xu8oh8C/JJkyNT9WKIMGBWol4qco2LTJ3Dotoqn5DgwEXG77m0ApuNztcC+2
bIoyxsEhFKy2yopA4H5ItoY6gG2K3ZtfkBq+twa3TedXcsp8P4lxSw2hMhZKDb2z
tTbcIWzuFhO9Z03u7Lkc8vKLNfeS/m4v/uqrqFi5POafybyl9BhatxqbS9p+inVX
uCbij+c/9rRBhmWPPLIbw2ovvEXCSMTpdMDNSy+BOgicJ/1ItIA4gc3em7McxWUs
zJx6P+B0KecsxYl37GXSXSR6dIMQGQvw4THDcjG2P/2H2gQqKdzaRw7tX1POdUPx
p5aCQRvLikqzLYKjQRFcCXluWRbaTm0EdeUwzh6NZeCKGd3aJ17XmPqIfj/8L48y
u2/eCbyyAjzANKBCfA+7wRVkPqzGY6tU63dSCUYRFleFUI6BZNodvYNtF3oyQiuR
nurUPZ7fX+IYqkOSpmSQUcVC9JpM7nU4cPCRReq8ntEPVtLUBPi1il/MpLskSHOO
pJlMGOi4S+VcHs8BwLZy6hGQy/sf5t3dOLAag/I9nvVJro458+1AUa6R+qXCF/bz
b4enXL0DewblFxpfGILZIzf/T0GDYN51s2juT7x7oACDjdKsQygg4/xH6RqdJq7S
EjEuAiD06605/YliuUou+ZJJM+kk7aWhlwh2K1fzPNLl9I3Im6iPOgyYTgqCKnyD
ElFw6YBaYCGvgZSHyUF5Wk2z23Y2wECPLYvIorlWSLsasLO7mGB+vsw6X60iNfhO
feDx8RorXARjwzDklfMpmhhcSF0dDRdP0e630BL2BozodAt8PGqXNHrfYuySbcF1
E7xL+P2Y8wrjO0FxsUtgxWJG34WvpgVrNjEyYOeyGvv4P1kDqjSncFhqoCGceNag
mqciq2RfcEYXqGwYgb995WuJJFc318aO48LZxG1+0kd4sbf+dQVQpoFBWZx/cQ8O
PPeZefPAjr3Pgbx/frqp2hUNnDOKbk33/rvWNxLZgORAtG0CMf6liQXRKHNG4/Tf
pVnVDbstQy5g+O5qMSwgrj2Gtvi9WFf8EQHuHNla5FSSJwhAMMuQmjR2QucnOzeJ
leOIxCnK5VWRNivbhzHu4RdKzI6eeVI9ggDHn7X0dgbHsikGqHeel1NERd9GPktd
tPBQL8QABle+xl/IR33HQViScvMlqXZeSmblnRiC3OfCt0QenUEPgujnbfU8d+uh
AJ9AnDLhGv+/ad4ZMOmC5F7N/PIRzP/6MNQRkp9PZ0YPiQ/7Kl2zpQvvD0//T95J
4jmAuUGaFCYGCImelH/FkSpBXKKMpn7k2U6tm/oREPGt5CcUjK4ncJgHH5nGcv7V
I+pd1CB0lyU8p4ImIdbNC8WAY8yNFMcOWd6bgLCSeb36/nopDWMcdKsOt1c5fjN7
1FnJhZ7k9Ewhgs+cV5csECowHQiEwqrBwfouBBhvw4vT3j/ghOQVTH67alcQjpE9
5RYVigv/mOyqQJAUekS+Z4gR/Mf6jde/3bwoCsRqeLnE+i6KdLxlskDGS1vvuHF7
AKXBQj8ejMiK5UzVfXIj206Mj+jB1dFUCJZcu06Q2sWcbtBQIOgyGMoE0clSj0/y
PrvsP8HwZbo8KaYisCdnwL1YkpG0s4KfrXjNYer2RaXj9yWGa4fmftQOaDN55WeJ
l4AP2FVhkTdaAYgsIHdipAq1d3r5K2W9XBl52GrVS1H9bTfMmlSALefTgzIxfUCS
Tne2n1aBiKv/pUm9OwMyXkOm6DO7UF6ZdbNdNYD4Vid3pjUzrfPmtCV4gJzPJTiF
NuE48I0S6Vyr3un8/ISjz+p0D8RsAsZDjr/b5JSv2s9ozg43Q9CBr6pBhy8oGN/g
uWMJZGFRWGcFSSmZU5KitCiPrKQsOUi5C0mnAB71/5CnSQHLqPEe7a3U0J2ol3Rk
DKmRDd4QRVzcPEGt+FuiTf2Vn8LLza7uTHMT6JPWhuPo6MvxD7lw2of1IhHoWWSn
sLc/TZmKGu0M+hb2Rdi+k8NFK+56TpIlEXdjZ84HWARQguB3fK/+kvEjS0kPwwZr
7iH/t9d1N78tj7cKVv1Pyu+T9o+KeqpYK0OIxyll1Rf3TSM8NCB/4tA2IBOO9o2Y
oq8I1Cv/BnGMY2R55L30FhfoxuBHCRQmb0/IDtQD9NVZdVEjnleJmA9vtUReOWum
KgKfrX5PFxtXnMrsts9d8ieMADt7SJNjwa7hFU0M2/VWICP73OPEKOPtL7bLvMlP
ACencCSfclZmn1vz+SmOu9cS3YPCAsQOxEdXPtiXT4O+9TVvpJ5jm6E9IJGeqx/6
LPyz/ox57VWPd4/OR78tErdJBHT1ZO1+FLBzh9XBkAlwz/SuqLtEJSW2hR6oD7+a
vxLxCqeTLFGajgA9RXTShY+zHS2hzD3kuZkm1FkJpWSrtW6MyH+jmk4J6ulwgpXw
y73DXwUimSmOrZ2bq16OI1OqGwX1NWFhJCoA4aCDj846piuhCI6XFahBxF2SJTWn
UZpy5eetRprLxKyhx0YjBtWkTYZKPSKSC1P856zzzshad1elpQIw58wX0NO3t5jn
MYLeNmOIXQbZ+KM9pvlbw+1xglaXU/tqbjsQYD++pu/sp9+RplbA8wbUOfjgNORL
UXv94j4h5+hrtNEOEzIftsSeeMBTBjZoEiFFeksew1I+P8JwFDwG/9p7yCvH17Rj
KGJwJA2KO3CMq3JrrZPl/wzqYMZlyh8x11WZsF5EPcWCBUMJL9O/pFrQJCRFL6K4
EflHIf/KSw1TG15n+VSrwxR1mGT4OhJIbQtyUqxWnnvFwnYU9eq0DbxWJ45f5eOz
01/op5dEoJdgYj3WHy5WI21fg51mz8/gDjGVpK5cT8hGDEpX/qWeACDIPYiIQmFN
60jRXuThDAMlY6qA5JB+1OcgdcUrR/TTadgcHZc11Z62bzOjqpUf91zhsPlCVtRh
htxwLzK4FLasZYvfi33LROp/XLI3uAAsGGHKQHCWomYts3lzvfhnx1E0piYMmlGK
9iP4w6MmaIVBjU9BNrRI7/eteeEwqedIVR/j07oIX+amzKJGr/8JNaGv1s9ItHY8
R1inKkqZdHg1RpIMivHfpPf2Rk82ipkxRESbI4UWW65tnu1EWbewHzCW2TbPaIh+
O0wBIapTCfm+0eSMm+C4l3bKTwV6G8RnCOOo5Z6G6lGdLpXW0ocr09IqywuM89IE
afYxT/v9y9SJMbEugWGgutQVzRuaYdkiSPma6Bcherhhb87ErGvic7CB9oKHnViX
RW/PNDurQvQsc+rnpYsS5DqasDtnoPEzpbCF+8XV0MxOFCeGRjPUFvnj5sop9fkP
580c66rUws/3ZWR23BLVrLrsqTvydk/f0qeIW9sFK6MjhnCvSaLVVGmvsUSKc8Rx
72gw7NXiVAXfCXx/j31pf7AeJqR99VQH8W4lCYD41pZGxgD39eASYwzryB94zqTb
vf/V+Tr4OyEJ/7EeiLrYmD3fOvG/vK+6muTcWHbGfk5xcArkXfuWU12tkNL8MKTD
SYRlIp5t7/4XsyzvrYMP81qbnIkfn2/v3RYbw1P+tSqtNYMqm44wLC5ODyLVYcmd
T+AUwG/jQHeCh/65cuF6FgQKfmA1roQiiSDxlemqLnBqCWqIUuBznojOKp38yusC
z5EDcbR13asU33C5jwQD2CEhAwoWEc1RFko3QcEkvZ83Qva/cKYJBGjyAEdqZrlp
Te1XA23zn7fKQcSUujq3SrnVhZYcGsYpVT+fLCI9fYIcNwkOuDYjo4p4IPPIsFvb
hcE6jNIZQTCa4Ad5KmTDroZXB0msPSsvONvcydAonl1IhPrIN4lcmiRVXPyGvhkK
4P0B9PkGcFhZQNrKh/DASWTJ8Xw//mHSU6wSGuG09ZcUEZeANFCI9DKO3mMIF/FZ
iYqpLqEDNMH/+YnrYlUvA1wEjy6yDDaP0oE9JSvKtFBZUSroH3S9wibeLBhrk6ZN
uWy2h8f68ih+FDzCE7Z80h8RD2YZ4TMyJS6Fkq0ocVLjZln49cTyeDgQLQ9c6zGh
Z/xQIfIrjh3j/5fYRZkmB2AqyYXJ7KBhj2y6r3I0FHYCyOwqBaftSXdsf4LyiiQC
UvRwuA0+59Q7U/Ih3Dx2PHYzOV3YYr4YFIFropMRKqssAMl2uEx2ZUmSWRsFyJRa
PTPrqflLdiFO0oZZSHALxG2wR4VKHyTsEW2M+sRDsWFiVdid3HVU6UHxfJidMGle
ifBhOyPF8agZ28n1ybki2IEJACp3bqMafnSH2Did6xLZL6TdJgFIcD3djXlfjUAo
PGYyRFkJBz7gS1JEm4M2Dp5YjY2aOViOIZQuBlKWIXqL7M88RCeqqZzbMjt36KAj
p783fkeWI1Xg1zesvZJtzAyln3M7KaFQS1Jm6QTxbSydkRoDRKjJmoUs6FxP9SAD
D+GB5+XJaDYth5OYIGChCetsfAZI5l4fo4jk0o6/xSdR92LK3mKwr4RBEPbuvinL
qO2yjEzqJPLtJQIJF8W3Dcw6GYnCFvL9V8jSMMln7o8MwxV1yP8axvJXtPNL7PRf
ilSthp6Ng5b7wjvrB16ymPRr36oPpPNrnMLZZpZAvd5hlGzDX3YXmpD8m1dnKZzT
wWw/V8L7f4M3XIEAYakntZoMh8WbrzuTnkr21dRm2EqKqnVxYZQ3ApHMYo6JkP7g
rHVTDHKVtt1lUdpsMoGOk3Q/Yv/pgdKlIagubJIgVb0BkbtswIEv89ugBsPIKd76
PCbXPyqJmpjXjc50YIdtxPZAoqVHmZ8G5+2L7rxcH5quY9SHiCvWi1eC02tpMBAd
h8q3OLOQ+b/6jpFth0U9CbaYfLU+88b8Ba5qe61np1RfRWLkeKIW17bxUM2MEQFN
VLJYEI1hJSSLW6QUvog81k5UAfIG0wheS38EsxroHOVmKweQ3fvTL2V00Fag6kNa
Sx0XGtfeoGngLgg5mXt/qFeLDnLpWWW57oAw9OIM6TsLcVTrrJxyMVmhyJm9A/yp
ZWlg0S3ryMpg3x6ojEb899V37PNB+QZ/J3z+eGsRh0mgfW8D5HyPc1ySRxzJrL46
yKGsC4lFOVeyGt0dwwSmrfMy/1qVCDMahF30KOxkF0tcyiPO+IftwRgKMKhOKF1C
jh8M23ZJnagS50JeY4SjgTDNFt88zJqUzC7CqzDY3+814vVJIy/i7y4z4poiIuqK
FXc3QozKIGN88s7/5OWE3Puoq7iy6L97UwEnUM1KDB4YR61CGSli6AUgflHambyq
8fkJMe2qQVA11tvLE6IlXqK8xSInL06DmY+MDJDt/geXdYawgXw2rGfD2IK6Yvyg
Y4/dD2lwlxRxGDYOU9nmtdKryn5e3PiZ4oPVzPK/zqQtrkEsZHl8LtiD0XXKRS9i
FK7MvUjGguKs0xDqTOBDdFxEASzzU4roOYp4x6MN9Ilniz9+zRcq8+8C/OlUjSEl
qmHd5FygV8h4UZfydYNBFGbFh0k1bTSP/q+GQvNG9QWU7WDlQFkhhvtPTdMdUymK
3H5tohhMC5tPvPoFPGeN/5pXGcJjAeqy87dHMljh9IsDn1N7r60iTcBFEXKdmVJ6
MeDG9AcAnhme2u/zNbDEjVu/TTcnRpM4E+10th1GN5mNd6xcdRpq6qD/j6If6c+F
6+12AfocootCyErzWpzkugzT5YJmyv9itFyRN06ETpTyR5scQ849jnHrbUADQhgv
Aj6Skvm5HHbH8Mcz3Xi/ick2/ngiQEAZTsXY/aNjr5wm7TqC42l2ExKNnF2RNUi7
qwg9zNG2Lr5EUnLK9E4XslYW99gvuw5eRwAdfyqBMr+lxis8MMksLYATU2sSL+5l
Mp9upCblglVigsYib5aFLEcFl84I0UVaTrFhalcgeeTFvaxA+e8MwGfx7vZD4cyL
ru56KgIIMsWznMgCRY2uQNTVaM34kY28EQJIou7qOI4bhJpJ8oSjR4+pm6AGMktl
VLfgP6DzxVL7A81G9idcpYChmRwDdcMDeh3ilvU7W9Ktwp/fzYZJH3a6O504CnpU
a7sTpyEptZE15IwhCoH9k3yaV+RLxImg9D+QDyZZvlHZ7+7UJMVUQr7rANDn4Nun
7Gz7ROPIUgLhpgd8KWbc6OrY5oYSZBXVeeUTcxh11+0LQl9yqnzLvlvjunhzlmQq
bhKPoELC7Hbh6YFo/sAOaJkehRXuPMm2qtdyDnX0BQBtxk5hhhyP2kjJxISZlYSY
B/xzWAjxcAb6tBNN2Y6pFwaKL0Efb7gqildQ/tK7cgKZ38RyprIYgJQ39Ac9R6F+
ED6C+IS1omQXlbYnKIMG7or22sYnZE7XGvcFZ3NxHZT+HJSNt1jkHMsEzdukySSZ
ycn2VPg6nr2GSaPCM3bskRQ26E65GuiuaOQU3WLSwv83MoHRB83/w49RuOSm4xoM
arPdNWzFLrGe/Y1vvKWRl5QKohl7cYAI4Gb85z5i+klRFb89W1uJ/H8JOrttuC0s
USGiPiW1BjCXKdS5VON6nWp+cpf+jGMsKwBs+90Cxb1ZsVasCtBku9P+kcAReBrO
d73ObY37u2NNUiDARxJiryzPC5C6xQ/NYOKWMb3M4wS+UZtL5x2Ik/80Z8DZykya
iw7mdW8HraFAgZBXjTgNsz0dB+vZ1dEbs5GTmQJcQgSeryKBgxMGydR/kzpGd7T0
DutOHaKIgwjLY95dFLWBLnBKm2iIP78u8KYZfIIvHr1K6EvzltZCgEUee882ZgIJ
YLxx/XZC/1P4SeSPHEcIm0JaAmJlkpB0riOhNwb2b4cJq9MrHcv6Rql1OSXiRGB2
8Oe80b0hQ67NgQU+WOY5Ru9F6iQoRFyuIyfFr9Ugs9hjvuSYrvIJrSJ9YT4wA3Pt
EZg5OOVZbTfdYMb3NEvMYIsAlnKEDR77xHDM13+0XxLg0WeqGjFRqEj3xInhscUf
b1lkVGbTIwmNdiP+RIs6Z+5bdz0g+bJJKTFsgFMo9/GDvQkqD8g/H5yWqQJkhW3V
HHfkOS+iZ3IIAZRcgVtsujb8C+J8haL3YA6E0FuiWMuTlilz3xj5myeIlRcyjGCy
gU2hp7+5Bcr0herKjLHBesymJoHOnNAyliRU2B9JVsVVaIXm8MHiPk4UF02XVQvV
ZEEOqKaq4pH6KuGF1WtrJYSsk29v//5OEg8fYbestJSZu0Z5t7fv/MT92Ts9QmYz
j2czURMqmMaoUAReq9k4Bx6EdcNgaMjFZHIyrajjNUOJDJq+42r29QvecgfyqKK1
q/0BSg9i7oAdqZJmihxr/8mT7lXk840R3iS0H4FP7fatazU9RyRpQCOtbf7hg8Lv
dnvimTYDlxnAeiYvfH83Fn2M6TOE0Ot57X1XyWynvVjCUU4vodUjt2ZEqu4xcatY
2+8tYSmBMFh8WS1xBy+x/QcqvyBM30eRYVesfRxR5qply+vbkTVwe7lOZv+LDPoh
qeUDLKuTHJF+6Ak9cKJSb1Af8fsRny17pecVEdUCkDJcfnkl1lS5TZLnFIll70I2
UTrJ2YJGC+WINGst/d4oSq+6NlWoRTh9BCd3ZPUBKCcaVrXSpwTmTi2gGyWMl/yy
Kiy6uYi28cIDx/AP2VV9smCqaRTbJx+gCbWvf16u97cUNLQnEutghsRL0I8oOtri
HYlZ8yZtKpDIlnerQWN+wcznD0x5wMXP3WDDE3dI5DQmoT4Nc7yMdnUll9AU8XUm
bD/I2CeFuafitSc+qU12W+xaJRkOY/6+nHmHEr6p7ok8qjKIRBfd4mRlwJsxWqJK
5pE/bdGJw3L7PqGNL/lj4LV4rrNIn4XoW278hPB7a5AUk9TFVaUIWyLpAZKU+Q0t
i7Fh3VCNzpd/xX8nh2VGVp/aNAJHUDyE3VGpr9b53twBNIrAMDhQ/gUbNBNQMz2K
g0VrxOcYwymsTlOxo5DSR2MJyy006x2Ixe306+8XhG6vlTTR2PqyDdujO0MBQF3/
Epn3cJUlMBIDYtQK4z7MIadCP322gF4UwhxVsIM2ZB3WHEOrSw7BmNAe0Y2fGgIA
g+xyQw45mq9aWG3uWzB4fD/eHvFj0bJdO1ERkiOaANB3DrrlDb6McS7fMH50kIiH
J3s8Pbh3425Gizdf5VlrnOKqxwFReXHr62a/duwP9XylGDywyHOP9a322A3WTC10
FtGYUv/VMRCh5fjXOm3cjQHARS8qnHQqY8Q1YpNmMXFIQe6Z+qPJYwjCySqqDUT/
ZRYsl0l2xbG7V61yoVgq+9+rNi6RHF2+ufq48Vfbv3oWMUJLFSJQQIDRA46h2U7n
7TQad4G8uxo7y0tUwAT/lVHkGRPi/7TJYl6GJDXSUkCAzUvTk+stRfXR0626tATD
kWvrSNuUhIeO5KIUxSprms7J2jpU80+mBW9cyHVHsYmof0PsApfP2jAEF+1t4k8n
RT8x3qNLH/NRzKK+v3pS8Q9n1VrWSQh/j2LzWtODPfetsLUF1hCZSQnNwk1z4wlo
wjjXlv4uOqmT/K9jGLJURxcy+aFpNaUjo4tOJCIhu0T4vExz9BDFvL/dRl5b3NIa
SHItZOYq803JUgLy3DKiC1hhTnOSHip/CalT2FsjRb7pgwPItP88nQ9Y6aOdWcWf
THOb5sklu7G6EOyWA60SIM+cUiMD8GJ2HgttVZFMJQpuIAIlSn+jkPcz5osMan+k
vhXAnyrscsuVzhZgYSHxYEM2Q2eWSEgtn+qo1KuCTGbFYtlJMEWZ61LUKprZL4eq
Ou1dgizz8KGaKua8j2j1MErQ93QdmmnXsvI4ax2Bpz0x7UuiIQLK40f5i7pxb50E
FcQEnIwHddIXBA+1iaAOnw5dD6QW3xeRnmwaqgXclWrc4LmrbyI53N5R22bxZPIs
e4r+MGOFiosX89e7cCQ1VXhqmDhROCpOi51f8GfxUrehLh3TfCufJ2+JtDfxsFtg
kVSXviaUzig4VjYCGi2GKXgKBGtO/uhv9ylmXndP95q8uYnFGAiWAA7KScTY4lTo
Mj7J8ny2twTu+s8rmrMVHDpY75YyaEdgbk+7id87xriKutzcMoGQLHOin9PmOek8
vpQC67fXMV45hhGswnukOW/eNs8YSbJBSmsrtywJAf7hdvj7ngAgKxbB2Q5S7E+p
kZY5A/ffU4lqW3vlpjVQXMAdIMUKbHm2aSP28QZFd+TVMiH6GTGn8nlreftms0tv
iYFLz2CEwkJZxZhMX0BsVLsCxS8mdxgukK8YlFyDjOvy4A1w6daIf3roW3UI418/
xykhnFig4zbBktGO+Spm2ppkvK+soqM299Zhpxr/+1rC/IzLxcqs06RvWH6mx+i6
i1no3VFoNpoRcQ3fzmLezSGJnHDnMQckZA8RKYlxyI/3s6EF3g2j5ihM4L13owBm
T3xrc55QC09ya94akl+hRtY2D2AMu9yjQiFtezr6HRJ3J1XheoLcCO38jcBgIlEs
A/p7jiGXsM3Y0xmpqy70F9xIJGiRZHBi1JcDCgbBVmLX3d5mtAJsXbk17Zo3cyh4
tlZXWKALXR+J7JjJlr0gWNr1SqxMvwaARzzVjOcvZJk/cG5h4q6IMcAW96S6rgjj
echsJQiAO7mgHyLV4CfSaIQ5tMTtLhUWpTvkqmNpYZ+KsXOnQhBYrogftJocaaj1
z6giXiJ1cecgUvnl9LPOmuE2swr+8OyDs/gQFJUS7Ar9uZ54NBkQm+bvJHw2OwdJ
onKjEprr+lciABbk0IMU210cq+EuvrJMvus8//JCXtioKbaitlCAG2SAaoK5sQxL
DmYPJgysdMsi39Hmvj6xMsK6x4KQUeFHuF04CD6x1R5dBIJLW4Zm55ALjWmRA6GC
h8SSB+SSTIJcJWm7sAKzVEcXlMG+QFf0dpQmlrpNV4qQZ0ibm0O54+p3s9SQEF8l
VJ4HLkdshwbcgutnvD1cbngcYOenoayaCXeTEZ/nEYML1R3LFUXBG/8tqmjAUG7L
UGSrIO0HyZ35e+ZL/9Y0sGWYgjx3AwpS9Q8baEXC19rOb45DviejgaIeMtv60aDK
ZN7JrIALEfXFT1ByzyUuv5uGYOYABggUMfr53Xv50vIimQ5y+68IyX+VnkmCCqLv
TpASlRvsdtp30ce2qHURZw+1wF7kP424bzVkGrXXBTZJl3PD94QcRPQjQLSpp8yX
sov3kUQsnAi33Hb1UhWkwfaslsbiJCv30LYVnw3qMPECu8u+r8ajXUs3QHnCKge9
y2cSL2uK5A8si3Jzl3ohKqZJiogemjgKVwdwALEmdnJ7aX6Ib7J9hnLszeaEWPKq
kQXM+7OGhyOprY0dlAqAjQbm5ratIw0+BfCJYyhbYb4mrSlDIy4YhU0SOQXC+m5p
yc774tnoOx7dhfmjCGuwUEr539qO2/xh9qB4cJ0WdJeD1UZIG/VYPoUXJCbTNc8r
A+66tuKlmsciV72ISQDWfW8uLGoAd3/hM2yShk2bDXb9uBgVEh5OAvtCqGz5MIp2
cYwAHbgCcZ61c14bJFwNtMjQ9OcxzN0zkM2mvlSlHszAmjxTjxVhEioEMKbw/7eG
aTi+CFgVjJplTYW56kr8FlADJirK5L1Z0mrWnSQqB/4QuERmgK9Xqqsoh9HnIuL2
4ZubfgAyPDI7u6X/MDS+LsVSJy9G2Bx/NwS9djU7PoUJQFv+E/jWbvQjNT40+cV5
ChSV141PjDRUmRIqnnLaKiL4a9xkFySQgk0YXiT71K+qHp2i/W4zDpg+SNw/PUzq
YUSD3pvrRJjQ/7/z+5P8wQhF1lP7/dEDmijYtL7iwZhodPjwpxRqBRGngygRCLQW
Gvtb0YsIkrHySQyUdm+QzYXFT4rvKZfwxeQwMrhB1YmhvC5IGiK1cEVldVARSO+b
RB/qtzcxV82Kgmfe+TTaeLZHA4ZDSGszy/nit6PgIV/Hvt5FQOn5fMoEs6dyfq5S
1XXfon8mRQ4JnbroGaHmfHNKZ2LfjAJFeETRsv9pmYBh/gmp8EkxpUkI99wvR0k2
i7BzaDLGVxQOBpHYJeaRyVysZjpdUFa1AbdeN8G8TCr9awL+U7qCfjVSEku+8lBC
LKGpHErZi2lhqDczIBrf+SMLLMTu03SUpknowgU3F1D95LxdbqmUEfhpZQAfKJxm
J78K0jSSsmgivw+3SqyH3XXDLa71NJNXS7GcmCPlCk4KuXMgRrbFwSd7t/STS6O0
VYFuOXCoz96nJCj5/xwJQD4IeVD8FdNcelW4QQXbPfEiULmbTVWR2wK1eM7oBGcf
+6Dt16wsEHW9yXGcyz9YIneV0sPlZG9Spv7g1Lp8Ja0kTMhM1OVJfgMLFOqdy/XZ
+ZVqT58gvmaRxUotLZJhHe0RBOWKJ/lcnJJwo6Wgt2Y3mx1m5RBMfx4vCPX7tRbj
Q82OVitW5KfjHYeDBNh4UNOD5ddyssD+gRpQNKTHI5Y9dpqmGMhEbBlacV2IDA7x
+OedheFCa+/JKBqefYR0eZWtnq76oJpAFtMNSMl8TRC10ak+8U/q6IL5hzVY+cZK
ck4XC7WUbYcNhuTIfIrPqHIHsAAPYIHGOqhv5RuFrwkGr0dus3tRfIwcxyCO6/2z
imQETfjah/FrZqn5glVlw94az1ieNig9//09Ou2c006uZ3iIU0MIcF8m4G7Wd307
uMSoUWhMTiczF62Kc2D/JuDn4D221z1u61x/iuDBy9HxGkoSC52zo+vU94YA0u3p
/dLNMxkk7kVk4+S7NYVrB4gSoM2YOUcJinu5UJ5RXMw0z33bpMgCU9kZ+0oJnL4N
rkdjDW16CHOxpOXk0Q1+9YCnwRuNvlblzEEKUdQMFpazkQVsN4Xp/9TbyIfrEBvb
+wThGpTibiLgtUuGFCg2SK4W7XqE1Zo6mcvA8KHOJoeThTyesP+mloHgmcOVBqiS
8vzJKUzQZ0JYhoxmYEGDcK1bBK3G0EM2/PYbzQ7ZeYdY1LfZW98esEJ7MDbhejFK
335mMzkk53qy6RGU40S/KC/9sbqcsGQjWyIIlPWTLT3yR9Yjdv3Vl5TLoSetAc7b
Ggldy1oby72xLhmisBU3UDkaXDijMrdsoFRiPvQvPoHmXla2h8dt0xyeTpK7E6Hj
p4YW1qn+PocrIYuzXL45TZ63vsKEbnHxXhJR+T6nVGlCKHheCOdSfpi9Alk3SciT
eh5ks78Z4d7Exztnic56+wOCOX9t20xdTXR5Szs+I7nDwbBLahaMDM+j0SBGeO/b
TugeQ5xVsdxxsN+SMpIboYTYdTqE/Mnu90yxjBatUYN5UnwUeB1k6LKIT14KR9f1
LH0OCwlzYn4E9WpKGUGY+58WfRlYJ4gDZnhd7SkfCC9MjrBhypJwV0NtxidoLgm4
bwNoJxhHWbwUsrQSetLhFe6xErMSDklPcOw67uINiiBWvXNxxRQEm86GivY9iB3Z
jAscH2Zbp8nkzWZgTlY/Pxhp+r/N5mV+R0wtoUmPHzKZFUWDTzvmA9Vp/9IXl8Ky
13LoxY4p/YtIv4OYxRLY1R4yki4OFod8RadmcWWLaffebyt3ARY3RUn1VnqUH/ub
T1VHwWwHIPzXm3/0jN/484pP/ltXgWNx4+rjK7Ux2dIuabI/D6K1uAda49BYPDvn
mW3HKMRVFVxlD7NdsOj/BaSmNi2ztcOjYiLwSuuVgP1lyz0WjU/Kl5ywz5sQGfuV
k+v6uudMn9dymEnV7rGOqbX4xvo4Ym6RIlPqYVdK0t5B6dkajalh17mMnj+tV25G
9fOOmDR6oZ964byORETEAFbB+iIFebtsskHbkZr8xYioTArAH7bpIIHa2IH7N1Kt
/5jOo67gObwCXwAz8DUdVPDlTLbRvw8BQ82Cqr98Wr2FCbsbC271U6lCzAA9f445
trYu6b8yGPebaHecjoIdN6S58pvO0ORHEVUB7deu0f5OekPJJd1XvEY/IRua56Eq
qxPPzeWQJ06XhE4wtrzFa7KxdyyKdF/yX7drVbTHLo6//grROqd1od16XnAOJM3n
IXp62e+W13iEfwG9leo7nlV+kRhj51a5j79C0kTwgj4EukjobaGE/5k0ycdyyCKp
GfStjMXduwgkC65V5HsiJV+HKR69dNEA3CrOLjvM/a4jJU7kzwygrquCencu/oTh
KVx7scpzauOlMOHgPcRO4i0FCkRXVvuEGELm/3OIIHPcVlmA0h+5BJILWSNfkm1h
KdNGwOHhvVaA6MWLpjs75xGqsSGAuf/6UExKdGbg2pXv2z23v1S+T52jZuc82wzr
O2C/FB7MCovxOCAG0A558G1Fw/bO60EXRssTVShwMcy9qPOZduPzv36OFFW+L2oM
Q+K6exr6zH/D99rNREc0oi7fE4F8pQlryuWAPbsI1YYrQ8tfKWsJAAkgbA5UamqH
MCduIkCu/hb/9Cu6ZyStfdwo7rxbOKqR9OMQYVmjn6ld9ovhsEOhEj+z8CTLrsae
BdqLgMhiSNAkGy7+SLmZGqX3NG0qCWcEWwiIc9ed5QXBtxMgs1QUQrZEvv5DUoBZ
gvckjOyCE9LPNwLw5UJEp9LF0YqPTsYAN+ILXnx2kVsE7xT6936josDVLMza79PR
LYK6I3D8U6tftOdDrMR3I0eL1q7mTzpTsEiD+NEjSFvQaatTjCm+Wojz6qTAVeT9
BqO1+5nnvFIRj7colZUyKMeqa0avPcaWYx1JPRExtao3B/3vfckVi39BR1fzGXx0
qq3pF9u0iUwVyPCL1P0kvDaInIkva9JMF/5/MlwbvohsNrqhHrL2/Q3wSR8jTYot
CsCbJkpdnDI2nANcetPEAMy4hqHVsLcf6eZjbaTJsK+xaD10RcSLSyl5k7WefFoo
tJ/0yCc9WWJGCM8mKS7B358gFDkk2QfF4He5xs/jZVyN8P7gkcF26OA74cxXKv3E
/A+w/AOpfNpiA8iQXvKXcjBX1eBBmCh5ea22Tz4KgdhMtV6ZuSppiBCzUEx/4fpM
XqZpQdpXsf51IzgC+fKQxKN+lK/NM+4BLEFGpUZkYN8d7mMYZMop1gItVrerQopE
J3P5owAvO5iL627fLIbX4yD0jsVA/ajWT6YswJdpz5Rn7ix16kPeVmmAiF2ABoII
dDR6R8TG5wf8PeVhcdYzS9D/huTz/0WZoVI7nogJq8qY4t/xKO1KertYoPs4v3bC
MsmfKvg8spsngKtr/oJ+QOHSygJx6V4FBB8pibrcsgBexrkxFhmeDZAb0SHJyTuP
RSkgGebNOt9Sh7hP0Jf5kZgljm3KlClxxAIFtDNJmSIrzV4XcMfuHvc1K/SZuXGi
OvQvjCu5ZVut+ZG0XB06sq/wjqTiDsFL1FqGz+8zQOee/454VombhFM4ZXugyda0
YKdYpmJGpVTjTyzPcOGwah745a1mfHFPqjGlplrKPy5/hCluUuM9hCYFsp77BBWV
19CAZvnPmPFaPcwRXNxZiVBMRG6zpO2DB2pKeaaQg435s/BdoxeCINtuCgA9VriA
3wo3n7EXmoAi6Xlp4xdIIZgqEa9rmb++NZCMsUQa4dnO1B6iT8bpgEfjvkXUzLeq
XDG9WTIlHbxWsnjkEkhKvG9N9oTKW+fqGXqdj5/fyOBQd4cTU/8Lma5Wt1jEO6zk
o79PpNHzC8r5iS01M8bPjSbTOS/Cu19IDGwA/LpibhxvtPAiB+U1I6bHrnkCWiI8
GxhmlvxgScP+gQCkt/3NndmcJMHMkYP8+uuL4abg6ADJ2mJQxBqS3nE95HaLNMHf
br/7IOsIt90fQcR1rExaq85UA/hYv7QnYtYBAwQXBdQRY+U30xtf6RLGX4fipKWa
57/K73Xk2WqblyVFzzqrk9vu2ud+teAWPzPN47CVuB23QkZVfPI0EspVTC1S/mOg
AqZtIPX4zVE2su0pouWACPhe3gy/qhl0BEzmPMCK4I7n2ql0+PUCS39sp4qMyaxP
x/lfeIOqkOCEhsdyq6ufE0cHC8XkBtNcFbQqkDR6rr/TmSGEyIYgEpfS9gS80niC
s9Pwia4RXkSBQLNnd8k6mP5C/02ef/ym+PbP2NJ39xkeudmPikULjD4yLZQOP1uT
U+iURju2xOr76O/JEjCL6BduQYaaWL6Vn1ln7iRq2BAAMs97etMCsZ/mh7FYixqM
wsu5n6Ptx/p/LBNaGZNsnxFYvcINtfsxb2yKQpxurrpKTQYuOjzVJgfXVka88/I3
BE6ok3dca+xfe26UX2KDcsoWERrQkbeUUdvcycmNrAPTxaWaumuVKOatfjhgxu6N
IF27xP1FOuc4BKFkfBJB38BZ5tRqGGIbA1nz3R+M4ili47im4VhQ8OQM7nE9co6E
PxHSCozRRfzk4d3M/q0YqEiyyfFzE2oBk3CArFkj1JlvYJMo1TQnNgk7Si2bOb7c
dzpheiBOmw4dKJyvSGP0qR8Lfo6Fo8pSnJtF1du1SXW7B18F/jKOMU4T77k9LtmB
tokXG54oHxHiN84jshAKTFsRJCIb0RwSd7qGudB6iZt9QDn1NqTvxiIrjFxrWu1j
YudJBD0LqxG9bH1d+C22/7L6kIcXcY1G42nazhgAlA8/zKJj5xF59SM3pC5v5tG9
6DVolg4TPHUelTsPXh/O3mnRTfAiX8t5U7DZ3n2zMKYJhf54O0xBtmfIquC5nehY
r/72tyUOstJAkqRl3b3ng/gxH5upaXh9azZwAONePdjDu68fyHjFym/KmbYkyCCw
ai+LgMiTNxdLPeD/ELdkKF0kqAk566zDAsvVydziMJArnaF3SRmZy83cmV5uf8ms
bkI3MVlVgwVR5uzkqsquXxOrGF1RQeVN1D/TkTQSb+165XfMoCH6l90kGnQn9xJW
pjyVmPqXP/H7JMxXJ7Sua7HIjKQy+gGsWy141le1E44yJWsY280RMJ40mcUBTeeH
NGTPnTIGWpFkXslYBFC0SnD1bUFcbm2ao4FoaxqADboDKyMmZom7NcKLW9dE5kUH
L194pWVJvThU8h69TBRBaE3exFrMpo/P0ueAmOxNXB97VK1hFUUoWmocEIyOgybO
pfRvQcHaali7dxtul9wm9hzUcokcHBD+mpfKUG/KEes9Fcsp6nEwnVCSYLN6H/Fr
abx9FtHYBgsfz9sR1ALPBKt7QHJJjoEbodkvuG3pL97gZBTHoKVQ8jPV5iz2FFZs
Iq27hViOeXLXfHm2zwKA28g5eL95YWAaKQIZXKqSQlLikxxnOB97lj3NW6fm9QrM
qQSKrRM5l0J+JpRUdrI+vPGtJwqB/+j+qw7enBhBa2fvHdQl/Q5muGXrHNwLMl4Z
htwg89D4vdYMhPO1qLinlxGZ8u6tFfKodPTOFa7yCAF3bwJe6xOCaZwV8jpKW4MU
/rlrf+a70aui9SLVinFkAsSPN29DVA4J087xxbmNbvdayfXUPELgplvA4J5St0Ok
5LNnhFf3vORWvWnhsrNhxF0w/YVWYhpKciwq8k2RIkhTNjogXyd7rmIsUeQB3M7P
EMc7BWjYhRnDPfUhvP2qhn9X84kq4vwNl6viVv0Yp7pDNp5JebTjpXUkXRi3x7CC
5W0cQYfoFBZP5eapNJMpmrc2Xw7aSneCRzygs3J/4129+37kkHvCjxrvvMGA6HA1
hbLn4ct2pZsrEx9wzxGC+I9Byl4AZk560G/yhOXzZjp2/fOsD5V8gnzo5EJxs99B
LzFUpqwt9tDdzpDRLvQENJLWr6LOwaOWUy4qCQ54NbOds8qt2igBYLf2htgfRw1r
UfvlixIy2sYvwPSVV2D5FBC/EyooXsVUhC1LWjKIgcKEnsmhcIR8lYAkJHJOI+Sk
xMHqNJD+079378Vsxk1nUZ1+Slmqt9UdVsx9kZRnSVzt4vGPTyxCzFxN/lPCyWLm
wd1NC7619vleO3Ee8r/P779zGyFpknEkeWoYuoQmrI9s8rPwhvoBIigWu911P//n
zbQEuZ36WrZ5Y/kZA7pkY2vVa9yXQssfFXvPO3AnEkaV+9Wl79YSu0uRPmsT1Oxr
8iXbEbxBp9OQJeyO7yM2qv78z9QubLYKv/r1sHWSPUHMHodXr4vV6wa1Odohv5/8
6VryXKhASydJ+CzrxZuzIto0tyxCvJnu4G9+0Fr5pShlYIgbKnM8sNidkSuFeRZr
zgyy0bdql04/TFjMjMs5QCNDNL6IQJ4iHXUUOypSrQU6yT4oVmraATWiDgm/fu7J
fhGAS0BpzmW+h9aOMEhzXXoN5yeLj6Hec50Fe27D6dASFd54/9LD+BMJ+UW0AYpa
GymsATMxDTxAurBm3cvSC36eKCjhFiZ9m5R9+GUJceDYtCIKAAl6tsBHDaCz7S4g
05njaUjVVHH71XhcotrIrggxrihlgQzVaqiwt5ds26D6ziTn/RUk3UREXvSi/5RT
AcewfsRjjGJ9Euw/J0oXGN8+ZWctbBzgqtiFcGXT9EHdpRAoELeqMQ+Fh+9iLA4A
FJPhIbweu13q3xbNPfXhIfP5bxswwdVE/Eror2tEt75dphjbJbnvudvjQ6W6hsUl
pSdJNBWuNcRsuOqf0xzqDcCS+Iml40cas4LTdDTu0HoneHgyT0aGChepT2xfaypT
npHqQhaJaMOwOMh9B2xGS++WP7OPN1rVA5Oens57zDdNmq+YMQoqiMVfxTfKvQS7
ZNsVK7C6eyXF2ibR/ZrgYL7cMakbHlnPHGdMZD7XfwR9/uwnzwZXcYU1aWDgkH/R
F6wDUWD5QGXwvGSOrViccU+NZoK1xWVfxTGV8/5qivGGgK0vYViJQ5tODq91rAKP
Jc8K/mbZzw76mW2oYzBaOY42yoZWX3a7UFMPrw7GB1vUsygRaxzCBZQJdoObJRre
kwEuflK18XrtZFic3rC1Sz8NY+j6L6nR7zAIkgs4eTNvZ2fHzJSf360zDChY4fEU
vPs2iazo0agXA5Ut2RS/6GTs4VcmMk57KeJhH6ZUK0JBwQj6ZuEZ2vk712XUSDBz
8S2yxEgUjISgv9I4kWUcmt50wV3MH1ZYr9dynk/x9+OvClaBL2UEpX+DlVs6wzpW
iXBYL+3dojojmle7daqPOwsEyJBvk1P7OjhfpRPLfYGzBexGdjlhekyLnzK4ghdR
vpBajj1Yu43gFzPSaKhMCq6qGr/MnEHVo0nSkhu4ScUGdWmZhViDRxpOA6SD+RZw
qSbXmac6HpkSfAdypxitPz1Tl3bnV9S12HkiJcodS22QKqvrKDY86/jC1CQFNK6n
UwpLtIj2VAW2hMMkJMihjT4Zz29WRgIn8x/YA6eMS0kU2hbOmVAR3SViSPUU2IFB
tFpK3XoDoHUmOh0GDgrF/wH4Tcms6oaWjTvQuFVBiPmD6tCcOfAIXFsa9mRzv7Ar
Q0vIFNiKm7u6GCvZdqlTINHO6Gq2b2CRmQpofVfWoLEOl+8EQdV84L0ob3xIN0g3
QIjw8uyonC5KEOWCKtMk8ApqFi21GKTIa7C+94wDQIh/5/nYVMZiCxm5AZyUH/vl
0Ubfk2Ty4EbRSF6YgfcViEGrU7/iJRzciQaC7JMwS7M5vsDpqBPVRVVJgAkVpaHj
qmmNmGhHgAvT0Wcvg6Rly48S1UNhnBrl4GMs9rLQI620aeQpJ80ae4/W/Km7Up+d
hbO5DlIkt/Bes9r2s1cT5cfYu5Nb89CHez6rMKCNCV4dZsQjjyp7/yQ5wpGciFDO
KvzodWA2AmtKMlEwNWFSxJUrB0beeMC4VGDQZImTWpb3JIGs+YvsUxvt9QWLhsuE
9rH196XBdMxVoHyQs9VxY+Y0C3fEdUOJ+GuW8KpQ3aNvmnsmi5Cspc5i9kZcj/JX
lR5B0e8aWYFeKnLUGI8fMfkeXIAsYLTkdDRkG4dfiVdn0IyTe7UrOYQxxutl6nwI
hPKK2+PpBqv5BoMx02+NfeCWQ+Ke7PppIKaX3tOrPWtwtYrVge1GkVEZkMAIgAYO
gL9Myl/1R2VqWEmBdbdLhA7OtRCcaPrVDBNM3qHRoVQuKN/4lGy2OfuZJBN65/15
uis4OlZLqGBq9GBQbXQPjuchYh+BoK/ZyF8QBHPghW4Xd3R+EEmNye4cytkHyVCF
5RntRlF0/6O98XBXqNjT6ZVjXwCbK4P0Qozk73QPe27RMp22kFpCUABW0YIAaD3h
N6m92iiIU8qQ7NJ1nTEHKYixCQfPx8cRAzxWEMUwYx034QlcEwoyAGpU/Ua+wnX+
8Zbzj1+I8SW4FFIMpQi5PwPOdoQBMjB8wgYk1oYjZlWYeijeIyIh3jSEwHCLTRKk
/6AGrJCXczPdROrZkRP05ahPxsdZk/Gr1VdKfNhnrqsVVitmK2NO2AznG7n6X4r0
PQmBlCupy1wZw7P8R6sk+d08h8EHxa3+2TzNvNlb9fHX++zNOXsFxnGSyBLOzvPZ
2OJLLVlK3l+esVmVeZ2PkJBkyaK3K7CQ0KqUR08YOjtJsxnazfkwaEZgbxcaTucm
5y97LIVaScARPT/AOZeq61miDwoPzkk8ZR+AFCLNM6vMz2tvP8ruYBYGhOQBJtA/
j4b2IAQg7dcRqwd2zvC5rGcCn19Gjn23A34zJ9+GxcwaTcYRwb+Rc6qdwpA0Ec4V
r0aY4Mc34vlznUECY1AaXC5NP5QmZMZnsRe34aK231XWOTr2vwLSHQJmom4+JsRW
GR7T5p6TfZhBl90RqymA7c+IyzJhx5jKejvrUDhhxb9SpmsApI5aRifetzgxFr5U
lyY/gCUBsmcPpA5PBke4Oc+pqDgFBbxQNIOdjseJ38GD7VydnbWSOpQU19AJnmcJ
RUerD6MPJL/kn55tNYjyNOuUEkdkjyfT+2Cd6vvdvWsZOiZM4QkjZCLDHPE4X51Z
GRitIok5Pzow/L0FYf4U6yEKSAp7W06C1w9fOzoq6pua1E6AhY1X5zgjeZqSPk8s
Fg6kvyCg9LgEjhioCLHUu2jM2Ou8aOaoQni2bbwfAb1pSwGnY9sAqXwMiOv1Shaz
2esn6+l84TXOTY4yH7PjcNqXWkfQmpTb20P0idFO9uuA9HEEw/8wKOzioWTBV5Bn
TJq97zy3IuVTtLTo+hnic1JX3jOSNIBnoQsxeqRaItUihL65Woq80LrmlPTsEZZk
ZrWKnd9oPjmjMcbzYIw1fzu7/dQDRzIecRyrPjoncYDcBjLs5T6nBRdQnU8jTBff
yTOBRe6nM+mxOEjXWF4tl46JC0lox2mFOsWvu4dRKB6srBquHPvnm/rxfnwv+e3o
tpdHeRIW/XlxPJhlVrOxc/VJtBSMZVrEoHP4TrCI/leGFgp/nZPa1EUMu3fLOF/o
0THDbV/zmPA7zrnxxbhAJv4nIMG08Z1whOV5yVrwCp1ut7inA0/ssTDv5tbRh+jn
PhQccUE/3d5t9u4NTSuSYmHBX0Fk0Or3/fYNX0nJ1uQeDznY0uFXfVkx99pENPBg
B4vB62OieRauzsmBEJJINsaD1Gf3kSQ9cCg81QrD979khGy33SsXn60lEmIs25pI
tWkXVLJjpbXEPpokEI184dv2CJV6G5KqmlJZpdBRllWnD18PXnIvuRqqNzL0N7Cb
JNH71cgiHIuSpSg4ovmD/V7HRbSWpNKWcLxF9xKRdzNlGAHKQ79j8GP6bq2eldTN
Xi7Cfo555iR3WsEAoOzmaKWWzX+JI2TaPsh2oOLK8y4Ilw8oXFbgieGrJUozFHzG
3uYWPiToaOd06HMaqtSDIna/4Vu7CHf7uG9710w6rdXxV2ABzGGgdSV/CkdlrgLk
YPON6CLWtAWPYPGhpxKwXvJl53F/ll8mTiz/BdX1XWc6kuA3B7xoynwdmWQgb+N0
UCzUbzT4XAHJNRFyu7BJcZGW9ZsxBhqy38m3MLBbmpUhzsS86DU1xnrGU8n9ChQA
SSLW3cS2BZCBap7VjkLIfZ22p76c+4K6fExnXp4HdDDZ0js1/xVQXcGsIWveN2KE
nsK5tbX/FG3opcxb5r/jmuCsfVW7ljyPrOssVdkDV5SM7kBSnmCAA0cmNwyNn+l2
VJ4r4jp8TUH88RLftT2a7Mi3aNBEvBjCN9+ky4QgVYcHyE7J0bnCcatRcRgzKH0M
t1JoPhxDWdxVnBqcEYhIMi73dzzqZRKZ03khtrD2z5GOTDQ5sZDVppSoGqZ19soM
AHyMzmcbyUE9/jDRsVKtZFpp97Gb5PBAOLsPrdHhYCJ3M75zHFdK1j3sJRFxM9n6
Q7J1OlXNeXg8Rup6HqFR/XX7Lut7yi+gjp3PxZGSQ3S6Vmwjyi1k548MAweA4nd3
CA+tZtH8VWBmr4TIXDDb9AVYcYaXJOqYZwjgBLVv3R1yscwnQ5ruyRJbzW6FCicu
yeVEj6ZxoMD5e8rjtKARai2IH+bVNwi2uk39039ywRBQIbMw/B6k8ev2WXpmZaQk
chr3L90obwZSd1MgMT6M2cj0sYB1Q3BpLIAlrbp/gbKWFB+B0B4lPBTI9hB1flEL
1p3lx/9RgRWLsWinKlSn2je9mM+Nq3LGqj/JnmEC+y/3Yo/Jz/mZ7DLmPLiuF0ff
sC/XmGgphm0z+ezq9h3cLDRQlyY1piJOCHOKsNuQFUZY9gwuhc391yYYf0dCKeQN
NCuo5bCloqN7E7tlpy6uyjMdZ9ZsTrn1Y3GMeO6zyO35hRp5D2V1xpHSflA7Fgy5
2SLei439cRrPM2XxIIPJCuM6kKO8QXlslE4RA+PO4FGY3uARWTxzsPeECzEZLjCq
Kx28c2ZRnIapijvcqaQKx30D5b0cJaDUQGqctZJNDlRWvCejw88iq/FbZX3Yp9it
1PDxELeqMdzr1OzAdTeqfiLFjbGHjmwXsFVGhmR91fppxdoNNKiUvdAmOe7Y8Wg9
yVg0pkr3QIWbEiw1Ca/i2+L8zgPZH5jVCp0qYCNm9nRtkpWn/cTNf+jRK7ofkSd4
Ft1eud9g+DAYOvB2j5p09wgUmoccYtdGB122cTfqBoYe4JCX0hdMK0CztOGfyMAV
Z7gg7IxlIu3tIeTtALxjKxSYBrmsCLgN3F40Nv8pL/8YqyLrDyUUvde/Vev5fRzM
SCmsHmKWQfIF8aPfiy4BsMDTA7N6AsHYTzKEbh541JMA4ixBQ9pqAu6BCzWCBwpD
U9dtnWQzJrSZIAyWfoC+yaLnL13pjWX+ofhRKN3SYHEWeNjBoOHEcD5rZB3wZvsO
aucUuW8XD48+JsN39cks8jsBUIH7b384bWNplFJMFokvSFF7S4cBywmGtpo//J3U
lg6BRpnOKpg6UtCa2hnD1AlWUyW7aorK8WS3BAj/HoUZLE4rGJ3YiHlkqdddfk62
oG+kDoihyWci2R1pgj5zk7Iy0hAukiVD7qZf4L4ugl6h6AKtA/qGKvHrMwc9iRHK
/JbqVOO9G4dw3B0l50wjHwCWvLmTUtVBIECcxSe8HH38VRX/e/3LJu/7SrZbBBQX
lhJbNaylT1+KQSCzRZNDuHRWbAcSA037z9mK0dPBYRs0Pr8w4mTiZgDWehHmV2wP
rNOLm9CmCEI+6QnCdrR3GwNj5TY9F/E9NCtB+OpKvb9D0jZKVIypvUojtJqbNWNu
YCkxURJGGuTIvY/T2punMVafrMRU4gf5Z+UT+NP/nnCLXKo3lY3DFJ9yZ8cQb+c3
MjFI1H8qoLFY/SzMqiaXX8omoVlnCCDSCIp3Mmqt8P72y/wTPa8o6/E2rB7gCeSR
f3AQxc/Bspu4yBbO/9HbOiT7VH1iOCkr/EzYmVrfucVlEdoAnqGnLtv+B2SPU7vU
L691lQJC8N92Ui3NS84Gf35DSREq6iS6SOaOJ7UAIDuJ2Ic3v97XJqacq4oZF5j2
ZzUvMsSsL2mKl0tLwRmfZM/2kawvwFQBIEj5jtem5w9Wx+xPF/lXlEPm409ZcRyU
/Fn1tKKQv1a+WcgxOHgKFMbLjP2e8RDFnDp2o0EcTlRjJ+uK5RTtgb1Kc03pLrXF
qgV8VXWdF8Tw9/ZvP+C7B7E3o1al4G16gurol+SwqORN6Xit7p9Th/WmEdPQeCu2
ooG/SbjHweO6dfjp8MWMGlz+fqJnvj6bzXoB42ZFaDuUgLgWLtSZMklNpuhvss04
OS2+m+gKv7qofJMUdoUQEKaKom8TkSR1U96dvko0bZVOlI+ZQZqiPS+pDfvommwW
ufOJRg1+1jLZRlVZecC4DGyB4pVX1m28jWtQDPYMnBcaRzsEYjDR12CDCzLssrTW
RD+ok0F5yQwC+eTj0QuL8lNwAou3LGGj9B7/KcYA+p2Zj6PFLcKO/ImuNJv5VdWT
ARw/mtuZa4JPkHBMjB+e7F5OuZyROAmb5krtnTy2i4Okw+GqAXIas4fWCY6H5GOl
u/KR9QixwDDvaC3z3O9ilzNbCpYDXi9rM/0iXdI3RbbGJO3Vy6EAgtntFudOYTNC
ksDzNQcmXkpkmonidZSMj/ADYSd7u2uzjNTg3pj78prpaynsreByT6DTjAGXpuKa
tuaTJmwUJPbyt8+RJp97wv5bLi/05viXx1l7/qRrXDKWUZLIzmgzUB9EfzWWrZhI
spa4Wicauen0CnfAlByD9haOxtYTo82KquWgX6H7Xk2RADJMQDkavaLDYXVR2lDS
8Dp6Y6qUIlpRNplfnWvvwOn1ZjaIGq16JeegHG+ZsIxbHJQKKK1898/PPyZHhg40
qoal1R/pS7c0XGMb73POTIbx0Y+r9BScbAlaF2+sdr2PfcSh8tIc5M1AA8az/SJC
zWc1i8mwuWxqcsYKNWWotx4vAMbPsmY+ITR0BVxcC8VPL9/C5XQ8bQ5ZUW1GdZmV
Mx2dqKA+NLGZedZ+DUYAAmhJWXvz6Etd0OwDC2cjMRu62FFxtQgytJMJFiuPQRQ/
0ysfEotnC8ddXrAiFJbfVkPcj5pRFQPagpIM/8WCivAK2P80KbIUVkLrzZziPmDp
T/b5BUSLSzMzF/tnxJVZ0ukGZEghEswco9JiNueOMm7r0huRefnvT8BW9bXSliuS
tZ2zylEv5zmy+C+V6i1nYj3FEaIA0tF3hY++IubUDvK2cREuCbnqplLSLoFh4tCF
l7F+sFaeTe7CkGZI6E6fj4p9wfJIcT9CFjPUPIu2VMG3xYxdCFO+GtARm0BvKwvf
VX/50UFmqmFPx9alxlsYQ1sQEfUsRMKaq7DRsVfQkE5fuGpEvrCGfpyq+ge1VwmT
nXNgac2KYagwZju9Fbykyzd3+npjd5XXvxZx+BfDyZUvxKozcCdTgfLz0E3q+DWv
XnMdkxJAoonUUP5+/kok5skSETgd4vzIKvryrHmAJW3isKDmAtMYjNp25anMYpny
3AcBhTfJbm55rog8sLLYrblk1CpU6G3ZNxYZ24ZQhKekDYUNOzsZu4DWLCmBJda6
4Dy6q4b6ep6Z4RxYQM5fnYMT21mNwVBcAjK9eYN2GTEz9DdFaGH8rCNplGLL82zf
KW/D8O9vsoNbsBXbx5GSjNC+Rzw4l/MmXptyRBqopznvpfHUg6/577L4jt9BJqkY
tDFJz8R5FF2BgDQlVdQqIBNADFgHlPRpCy52WAkUs6v5Fb++ut56GmPx4HAuGCRP
e6jpb9L3R4yuGdd39CDQw1MpDXKQ0ZHZAmhUeayhgrqGm9kjxaAvba8whmmonHY0
7H7anmRkhpL8Z7/wl2xXg7KJYyCNpobeoHUQi63fyzaLKcUp6a7DB3RB8DVG79i4
i63SnJr9bZJuEF1q3EZMLjK2v2viqLa1xFsKCjqYsknPOXW4nt3q54oPNXs+xTUk
mG17A7ECLupZTCFZlFA68wyzE8eA8ttocHrMA5X+nGc0o+nR5+6huoT30umzNAns
QpuExX0cfDrLakJXCwaAHKtKpc8unC5DHtRXHQ3qkoEcTvKrZOnoRT+Lahqk1c7m
MDwltfHOwk6y/WbwevESg3VMVk0K/PfPT2k4hL58gzvZ2iMbzI8uFmbMOBC7QTpt
HzqqLVu2+jq4/Gy/7scPwmRUEX0UxkKOtZ7na/Hw4vq6z+0CMlynPDPP8eUbiYLJ
ezA9XNSTt74cp03PvGAgOn0hR3KfWtyfbu1pZqeyYAYDkbBAQOxo0Ak1NoRYrXYW
LwAHsJUDOfyVnu29EFjcqVcFMRotb/Fmj02Q+Mnt2j3bHYnDkx9Af/rmh+KXm0wn
gwzA2O1t/UBSs3uWi5bFblKkDhmLc/nD5tqhKduMr4oU7i27oKMmvG4Tm52GVY9U
LpVPiiwr6crdYhuNLKFACtOJLEtIFMMn7bhZ0McCpWXJ3xTQI3d3Qib1M42C4xco
A6YZFYOCmSxVQuyfMKBjS0sW9XFu/w9FnSOn9fZqWqG/jrkuOm3YRwyXSz23due3
3k5E82aGTvtV6buM5+5iXw7oTGrWPZtNhyx48ZEaVSt29ExVNOfHKTMhlb8DMkDX
M87UNvm205Rfuihxa5Dzvo33OO7HK6ExHUKzoCVBBV+dAQN5ZQ5kYSpx7NAcWvaP
lPKqPhIjF901FjxbjxggIWJ/XJpD+nK76ISg7EsfqvNuFF3aQmSgGLyvXeVr0Pt2
K3piidbW3tlbFMFxwc/YBnINI5cZv0Woaga9IDt6ytemGVfw6+oVZFz62/snEvDe
ocb0L9Jywdt8ptU7FnVSCgIWJnSukjJvriT3fnRpP8Jj6JbMBP1hMouc35u0XwmS
dSDNuB2ke1jqG9X0Wt+LtPy5Gapn7ibBO08xWy9khH7WFoZ7rDZ5vvf7IwhVZOsr
/3nWPNdQhDYY0ZfbEWHBTX0eYP31XHuN4l0bmc4tdZiOdYPZXLCTQe+aJ+6nScU0
7V8Pw9USJjmHogMZlFEjcNyZBRRkfe2MB+us9OwxW3qqXffq8ulmwS/fFJPsHUae
HBKYqfFSMAxy8JAak3TqpYrGUbGFuLAUOka/Ixy3Jj4PMATOkzqxwljVgeanL/fn
mgUXHPEC7iiFjTtnPbZn7ehXv4mxO9hzuthULgqKkCbuTdh7obBgz2+nOzzp4ALz
5aBWQcYXdpregsMxKa+N9oV/0VX3kXpro6+dIjM1cqXPeK5IX2Pe0PiT2CwAqF2X
DlUO8vI3nTKGjlWwKkumKD5KHaJNk1YMNqswsmzjoiJEQm5fDoc6ZT2cVVLKxdAu
rlkW96pWKWx/d6hoLsSigXDJD8QQvOvhjmkvURewntqRI0dwjRZbWX0K4CxVmTMu
6b6/ltXkLtCHoz7VA2yq+IWxZM6Jecm6DSueC/mWNqgLZ1SgRfzza5/KMKJF/vYO
BStMTEpESJA1fZrY2EIaWbgOKy4QqVySZ9pdkZO+EfI1aB3sGpEHm+FnD/2r6J/j
tayPAIHOmas19ud82jIkyL6nyeltgNMLVJ7ZQqczj+w5FYmp4g7vZ8lSUXXrcYHG
mHM1SKPnUQHptbK/7OX3HxJsuWL9Wl+Pl0tDK3ur0h7ZzPHoEIXBp7YoUkcjEOOH
KD43A+LA1cBlaPfu2KGPhix4GwjhJOAsUruWNA0jCM3Tk/86rXKxqAO+yBKsnC1F
fNN/Pbkvu34KIsrgQoJXTnf3/xiLQLWyJs1eKeyIRQYMeytE2VCpKaPGyWToD4wx
WOVbmhjLgaQp5FO5ipdoxunXdlZ9QZg/ti7FoXxshrjYa9HLFGdteusk4xGIpEVe
kp6A7H6wdqjEmV19ZF+OJ4g/MFkSqHBUILkPBrJxLoqUabmyPclD4UMIOINBYsIF
J0kk19op9gVQKzJ8i9vBi5R2LRsMEa5Z46nl1Tw4IFkqesImxXMpHyxkfyk8OiBZ
49HQf2+6hRjFhzKADE4kYVXVTi3Oqfibyh/EHkS6NrPdT1WI7jILpGUrim2QzxEW
iofKZJ9Sc1eWlVLzvV7H1UO70a+zFilwetdj6cv8PKNmITZPWs3EI1egr7NR97ea
w45w3zJ6WhZKq1WizMr3Yk6DDb7n67j4tk1OShoxJYJiM3OdrKDF7c8ycR3X10Q5
QO3ptZTb5ZRlHb3gALg3X86gnCjJchnSIyhB0JDbZysRTqxfEnSNai6gCYc84lh/
zxmf7u9V3c/6GRl4rqIrvF2fD4aIkBbBzNq/CIiy3hH9zgESFRGqFnQ8WagbnxtU
V/cqIWRMZN/74mzZ3eUMgyvFVdJA70fY5vMhLMpZRXA36aWw4MrbHHifEulLg7+c
FYlyqL/2eysVYWPHOuXARLSlAPise5xKAxHwCLVN0hcoQZssjp39wbED0npPjraY
pVgvRdDyIYHybopInyy1j1DZCYe6nT280VsuPyza49DsOkwk4nwndvufxOXQ6ICU
9RhyrYSaj7g4SXe4wuuxW6KYM6cGI10uaiXh9P+pJ65gDT2aVpRcYjWQSBoXLbuS
IiYrPxIQwxWeM1WW49VBe6+7Ju0Z34kJClFA0zGXXK/5+A6f29DNLOUs9UwSpbKp
GwOVIDgD9Yb4biNwC2KnkieG93Q1q71tquVSHQTUCOMMaql0vEoSUXqB0bWR4You
yqHU++Q5ZTUjz123QPhsvw+lMNEzGaBQshDpykeP2CU/rOOMR2zpvS31Ee1j2whQ
dFphImOU1CDuCdQqyLnSqpzTKi8q6ufUjyinTQzeLE8a9NwdQQZNCs9UbpBzw40m
lZLZVzDMDhvJKI70UdbA98PpaUJyNB9Z0GXJtMtNvi5q4DQWZVxvbzYCwUcj4Il5
e2jLPWxrqgLLkNIaJRX9VKWd0hwmI99sdRuBNdKa2u3KNwbEuhQ1UYrdBDbq7ikn
NuOcSkqIng8ZIeWaPtX4ehuAOtWSB7RkOVZgkw5QRYsYrWdEks7C+mpAp2KXpCS4
lEBDpMUCJB3l6p5YPzd3J85IeQGS6A3KhP/OmWQlDns5QiQWPQ+Q8wyUOQb0m8c8
RXT8CMLbIsErkWEX+HwoYVkmvP3J3KuoqIgUPAHDYIlmBfkzWTfu1TT6Odth7qYV
8lUlq72+XNIMq+raoOWSEqyKSzgGnTKlM4fzW//ABALCJPZs5R0Nr3lqC70FhYhs
y8Yvbd5+8bfbtDvrHc1j24958ALoEBiTtVKjeJ0fSm7ojIiiQ1LbtQXgfRMPXAla
ZZfa7M3zzhjFj4j4AX2swTmRFAVUy5WB77NJruk/MrCErqDdddJI8+q1fGnsMbYV
t+VAF8Q7DhZIh627LcEYqrO/o4XhTOCiSrkx26oTnwLXjDd6AHCDoc2vFHAeqFoq
WKkmrusi3VtIcQDjMkkugyskuuVPsQmFGKjNl1FKgOV6brIAlCUn1onqjKEGnU2I
WZBEae4D/l/J8/x0sPnNjFZHx6SH7hKpl3keqF+EfIpVSnNabM9uqT/8ec+lY1c2
NiM5Kle6BMdOhGWe447FsCfnaLPSWd1d2wLbl2J6YoR9oVm89db1eQf695UQbzly
sUSEL545F2mpk2Z6XBEhVOqLZSXg8tGXkIjPGcecoorggSoHGTuUgdW+ZsymZ7dD
y4NG3SqawvQKUKpC9q+xCKCq2EXftgTP882QM/pFeeB0z/QvLwMvfFpgbfbG+BXd
0cZO1FsSS3hficXkG3/YX5RXwI1areqXZx3Y7wzGzSlb+4sx8uqvA9q/HBRCjyMN
49PKNAJQkzKb+RLlTxzQ7QV0pIK5pXp9WpJS9ojNBt9rEUT8zEARd3kCKAX93HOs
r0vtnmlDjcV+eDbtcIez2Y4WUOBZOGtpldjKPFu8HfSFy95Tb/r71ArdXScLdldJ
Uv8ETpFyYrco2mdHLUHOpVN/kL867Oun4nTSNUtCoGpLesEJwDsXRbOcz3gEp2Ff
8WheibBeFKlPKoDPS+/pYxBZiK6Vxt7xLWcRcpAsJnX8Fni5BwwtMBvxA4jgOXzB
bIGMFjMpffmJYy14I6O0VhCSHSFZ6wei2n1d7lSn1tFNQhBReWVZKKUAl4OPvsOp
vO+uVOLiGPZdsm2yMInpxQUwFwob+xanX7T/H5cad7TbrBSD7l1osRSDVNdlHKX/
BWxnsWv5oL1I2YIs42w33qz+ceFw/dKFyfzQl4O//dR9mQBARKaFicDhWRBoGx/v
h2nrL9BVWRYZhsVlW7gGpIYVTHZ5EUeIEX+rmx4u1WIaBYIAfvNqqVq4QCtzVvTI
2fP5yCeWrnVDh8xLRU9aTDKg2efO7bIPp660AWtuMsxPmgkYhVHBxSwFwb/cx3ja
ztRMFHYEN5jgmMvK4bsEDMLLuduBIFt8KvKzUcPOCD8uFNTi85ryK/W37Lwfyhwr
F9E6AmExuxTPNcEOHF6ieX4w7nPJ0ut/Z3OAHvXx9/azzFDgsCrsbz1meVWN3pm0
0P/WzQDjbMFD2C/ThhOVl02QToQii27mO0kZRazBqZAlHGyRYuENdD7CsoLUj9fb
1lPca8f4BIKXaIGN9pgvaynDt3V1eU/fkocd3WuH1P3wwHqpHur018yhEmAe+T5+
d6aBc3K85j5kdkUp9XZFWcY3lKNP6RhtaEGYWVHZJmPPignAbkfgT7OJ6ltJ3aBJ
Ws4d4tr5e+gwTJGOJdD5YsEx64sAdsfyGUDQshQ9qJ7nvDhehsbHGOteRjor/7Qo
LV+IxdCN1ccSpiVqDwe/ynfUl4vkepDgJMipr6F48r/oQbWLUYqHRixufsElgKvx
OpVvdyzIL+kPRDR5IW+N70vtFUn9gZ2iqcXms4ppmjWnlFiv9//lAo+Oahu+eBPd
BcVpCo4g00NzXGug54ZpcvpLoyMNOpOzT+Qyxf4URIgWjTFEb/nyConKg/HQoOiv
nR98pwkjB0GkTDKnUutv84wut9id3py1pAKkuQetD7EMQDVb2Y2iKgLLr6iFKIwf
XZgjj2cTgLHDUN6MqmdNK9q9j7FIJT+IBSqEIodNPgJJMwkTBQUk10iCXRlA+Ojc
umbqp2cwc+FEbecFgjOk+TZwkKUMWpajeRJYxqyEZa7b4huXzS9zwkSuICCKM40A
CYSyFE9ZeJAAYCnJfUshY7p+VWxea9pDf3/GPXirtnGTXTm8MF1aQd7476e6KrR8
fifj4yfPa1meSYWFJnutp4vK/ut/tXUQgGBLrxVkFjZ6JhTZA5DIz8cR+lj/yu6/
LGZII4mpjoOVcXIPxsDT3EJQAUutIPKE8lcnC2PE/3VyIHSr7+s8UFRzwYILjC14
O+UunX/S8IB0x03nkjyLzCHmSdQOuEZvf0r8q5vpjH5FezFY2L5BTt1q5N5AS+YS
dktfsOjxh3nKvMi7AqeHd+lPGkr1iQxAOZAr4t48670H/CP1NtVXKLBxcDy0Jciy
5coB3E91HPjW4md9upRZWvyYi07dNS2pP3P4ifqP2YkEFTU+Ojnl+7xlZPMUTz6N
ifmlCd95gefUPfxlLMTRiThCABtzadlvTi+/Kb20ioPM8jc3yzG0tyZCeYmSbCap
C8oPM/92JPoEljn2ug7RuvQb6vwWYpijf0kXNpCsjKBtOV52PBVXRE4k9nZ00eNL
2vxvRrd8zXgb0nJtn3vNXrMXbn631Zp4wD5o0baDIx54dPMyTufeEjQQ08QbFelT
FRdNNrZnl1UZZrub4m44UQKsD3Q2bXn3A7CfS/nACawQ+3O+uLJU4NEpjhupPzLS
2f8bDTqjhaQzEMGkDTVhDiLsQRqT6TM6VmYN4R5dEGDhPR71AR/voamjZK2ezWFI
WTH3Ztj8nyQFNYRwK2W15DZE0fWdJSMz9J9xpB79LC9Ck0fLp67k8VwY5cYURqtc
1oi6Ky4DLkmpjq+pM5ET56QLYn6H5CxwyDuLk6JLFsAFKVgK3vlPG4d5WRwSlLZZ
Lcm80FP4NbDHLLCkD2ZlMvvDy1t2XF91TRl+iPDzGBGP0m6JIRBLkukgkLttO/k4
Kuo2rjqXFLrQ2h7zT5hSPoNNZKgd3E69hZ/YnC/2JgRIVm4bll7wW3HtLi2idQdD
w7amDPXfFAS3bBUTJ/eHhPmWsMdzxmkIEE+imuw3+qKhD1/FddZI5PvdtPEXy+Y0
u0TI7itKgItd45GyF0UKkIffRT6fFJicR7i6ggJ7XT3gCiPDoHlIsJd9MRz1rmE0
60uq5z/K8CDSYkgQHjOG0RWAshT1OBw5YGA1Gvqj4JekNa/aLJMn/XnzC3K90JRj
bcw6lXP40uHetPwgFJ6ZZbWjbNwpUYg0dvf2ubN/8GOH/dCDq9TjngQndPfli3cx
KeO0JhW4TRsAVrerrKa0Auya/0HYo3QZeDh4IeApbzILDYH95nFKPcqB5UJw9E81
nJVqrVpIRKmn1Nk6xDuepDou4Qq56X0SVMp2LCCM66D/Kl4IAeyyE1Xx87st8O++
g420rG7yucS5Pk8fU1HjZF2+Yn1MRB+LsAyHGYVwtOXyo2Wv8fK79OA1We0Cyyqi
6e04mKg8ZHb4Nv5Jyr8mAlmpZjUHHZTx7Re35oWxb0MQr+PTCGyZv8xBF36zw9Jt
Ngtf8MuhMo3v2gnPXDVCv/p35sI5ePvtWhAPJFjxGGrLSCS4ZHeuy59yCfxkkeph
5XpqeKfIRuieNdjIUBQOAhk/g4FmR2kxQsRakl93IjBFxRkdkC0r1hSSYZqLocAp
zTRVh0wTwytfsBGylB1F4UNI+Jhmcm772aN+6emA+NvBqrEb4/cOozzDPX/PTBVp
HoJryr25HEBXMO14JtFLEeleviLT5CgPEaumTpL+DPIPGiqGyOFkMSTjED1UOBx/
WyGDS4kok/V8jMO8l00FrPjn/AfBta4yVuBrlU3aYs43E4rRxoT30cxBAK87+OgN
Oiqj43pyG8Mma0iGd+0KjJZAvVqT1dwPJWOtStevxnSxZH65RuLkUalq1821z2kA
NZXpQhAIUsSc8QU/Lg+TAzmQjoojc7YtP0nvK/eL78rkt+akWaSzaHGYlndTdAS/
Fw144XAfAnRd/3WR8PVAf6DpSnGb4OUKFbcCFBL/j/VNdJJIjON5hlSix9QNTBS5
lUmF01ydONJUM0z5nqTTYnhc6tkWVcLg8oYSGZ8eg2vzbl/YdHulcFeKiYyaRcaS
Uo25Wh94dNON2J9aQeOrrsWre94QNc79zE8aYNbz9vCbk7drJlEsATeqyYa2KAPM
yEARScYpuoRpQQXMqOYFXqR4/VDgKxSVIaw+9BIYqKODIN/piT/7H0vbzFBkdaUU
ne3e9kScovgl0ouRwhg0gWbeI3K164C6xzKZOPobrJK/68MboVD7VOIhjhBvl7RN
VlHkSFZLjEeTolQTLKTQU+JWBYRv+FkvQ8t5wFhuReycf1LeJEGCxEfso5cPxrdL
/5nfOYWo0gbAAUuf09YZQNA64WmtQ1+AtOJVX+2OEr82W8ruFp/85sMVlozMJWko
qLfm9/OfSGSKq/yxyx61wFhXAQZdqhewyRFKuzY9EtScH+t/Fw83x5AUFRnqp2uX
nsdEUz+ye/P9TiUt0lLJk9hyeeE0rOxsLE0lDXLeR1k9iL4cHDOY6Bif21Ctjm/5
kGo8eYO0Q29FMwKgatD7ZAQ+SYrBb7EFIKXKek+1LRPn8zXdCVtMP4FYTpXfbeJl
hZRLSVzkcvR6zYxia0PphEunRz5ekQD9JYLnazrvqzE/fF9g9oaz6+jNhtu5bLab
iXsPRmtgFHxLp5m4mEW50wBw5dKpvNt8pv6JZCh7GBHcZE6QT3dy3smTzRRuJtHV
l4jCeiX+TjjET8B3PtMBnzNH0DC9+QUl5NVprHl/0pgPe81RlfEPBGlQjxdnxQhV
TX8NgekR/C7uq+M/aSiXgZNeAx0w7N0tz+kKuBiRSU60D5voTUd+9jyfsVFQpWHg
IJsUZiZfajfAHcw/rozwBQHswQDtCxUs/e5BaX19YaH8xTCE2fGu+Y6ebmtrD+DX
P/cAGkpc+SgH++H92qyT1+bTlu11LKAWD0mGu88D6rW3oz5WY7VhBT+ds6ZWdaL2
IMPMuM4HVEjFNrs/5u6KoxziDmO0bXydGLNNM8rqnmQU5pKDv5xCuuKMX8tX2ca6
nb/e+gkWidRjIA331A7QaLcLb1tCfnW4IV/YtwbvcSJM9Ct3L4EvDCHfLR5yZH4u
hG213Btpjmc+zKGfpcPjYw0OJKhSbuiYbFstHci26yydLXYlJvnHsWkw5p+PrQc1
P2yQArFPR4iyc3jAZmqsCCkrc5k+/U2pRGvCbtcA980rjGhx6PtWmCio7GjoMgDG
pYg/vdMGOu/Qt7SXkuTqIDV0wmMGFCIVaYFAEE0Ix3XKYS8x+LyDpEraYjsywSQ5
RDuGTcjseTOHoHDWZ0TlHlgOmjHC2jYs+rEmKrYI5bgK/i+1SZrXi9OShujem88C
excNpH/MlWbH9pBd7ppGSUdMYuFgfzwp/Pl3XxWpERIpqPsWE0WiH3WnBNj8h7yH
+fQAGdcYaRyrIezVmwyfqIRNnr/d9QiN/QfP1p6Z6e/5fFA3pCnbjIKaYT6D3YCf
YTI57Y7a/hedOrZJpjcscd3HMeZF9IXrq+QP7WjKEL/bABc9YhY0M6kIYkTUgWRQ
1L+VgpT59ZjfaBl4ViXK0A/mpC1ixQTtdqkagE1cTvetoadDtivyp6qKQ9xASMxZ
O7uvmQMVXn3LiypY3HO3G8qmOJfpdwL+2qt66ytH8rFq/VSdXEA+NEdH9tmqbB7x
fxtditFx+65zb0zEXnBVe2WmTHiv+bpB9yYowXOVFiN+woqXoT+sE+N68UXKVtVM
UFVq3qEzpOsrYLYJMfz2yDNjex9GL/tB05jtytnxc4nRWq+/UL1mQN0q3RLpekOz
wWA27lXWiSZapHC9Em2NZBzSYNMCVBPQ2BfZMzznJ53jL90sho3NgPmnL7E4loiD
Rvgo98XXN8ExdUVkkvt0bmmM+RZFrLhjX0+sL164LlWGcmw5unPZ5nMWxpqjCyOq
q2o9zKqn5D0OJ8fKOhQpJTcUNzDamVAvM+y3vbCwyEJcWyMtXM5QSgeaLc7bbGlE
8hDSFUKfbZYqarOKxE2sIFeqr6LPq/D/W8SJudL1+C3+9/W+WyucQXV7r8yBIWxg
26YwQHu9wHSW7nKiVw5bGgbBZXaib9nu/qBNbLGPLuLLPWaOjvDsKHDRjhC8jhyZ
r/4fM4vhLq1xkYAP0/0JLvHKfddCwOk79XTt+/oebsZ0Ycd/SXTpYIkcLzdxf3RI
AaOx2h8D9cmxkoHVznuzMLYdV/SJZ+sD5nuYHeHQHi8r7Kqkgl8uTcpeixC/D2lo
ex/eyl3wQZynLuiUI6kEUYAI5wI4LxNevd6OxZQWhKV3p/7wfR20E831yMW4lHlG
mtz/TbzmLxy0oSK6U+Ti5QDP0OIpM3UkT8Us7yTMFNHtaxZRQ0Q2KA1mANtD2NGi
MLcOfmwa81Ag7q62g/GHcLzqaObzjLbw2Zq/Gddv1FSSukmZdUcx1o3FQtek82eo
/ZAH/BQkfEsNeD1j5b0aQf9WXWagG/JDtViN5RAItgaSFpq70xEZMfBSplkGIjGY
jaA6IoQswiqhc3TFSd7fxz9Ka1EPYHXCa/ZE7upYJw6qIPIhC/Vx0yjjcmf9ypGg
58tOd4EdBMCACqSda+sF2WHUp3FboPjsmLL1fiuixN3dZtMYPCfmV9ntK4kMGMn1
KeB5iIZADkYKXDuHKJSXVee69eUvXdIco0V99RLbTQG8340L8J6ljTIIblkfIDSI
ApOWbLAEIS6cD33r6N0P7xZpDBiCQqWoHW+v26kuYJ+ssOWxBmhSUb61Yyhm+yaF
o8da5J/fLZneeI4ELXov2U1uxlaNDGXUKNMS8JuVsuW3brHdkS3Rj3mP3fYgzzvN
ktzfD9Sqyccwlmb9qOQhz1cZyMfnWMoEN23zf/Y3eJMbBAoRFMJF/2hAmcGxCQtG
Y6kVWmd20aYzyDnum321rmJ9GOjt+zZJbpbgIyqbE+So7CXKU/fYoS/NcBLB0i9m
4FehXJCQhoeEDGF9AML37o9hniOVoQ+43/NkJTxpVI+D3GFx1QKhY04ZF33N/urX
2KvzfyBthUF7OkHJU3toYZaYeOc3g1uqr1TVH7lkM3sKobZACWCkzPhZ5kqb8HYy
N/trCbdHpWehac3yJeTkac4zHlweJRrIptP1E4u96n55LjPuk/ZAzFqu22bvE6na
TYeQboGfahady00XDbXwDIkdyyH2GuDZ775GarBq1/w3jTknA2BfKj67FYVt1ttt
vn3MCK1atze53MGax41kzA33QikORjiD7evUEmjAUwquGkK51G1bU4o87u+Cwvl/
jzLEhkS7TDAx8z/rUIJ8GWmJr6Q3a9uzHm7jg7Ll0+jOb9tFQhovRJ8k8p9WjvDL
g7L2I7V2wctC8M0Hf2V13DNKnYiR3b/ggMuHRyqE4gm8ar4ue5P1aWMoL5L9WTDX
5hZlzLeS+LhPSI+FfE7zNWInDqJ/4iADOQfRBYi5wkpw7qez/XHFkKMv7gsjEzPE
6fIkM3kP1jygvDF41UCHEOiP0p9qP/VxNvJkMB2HHcX/embzj8+1nhPNn4AA6uLG
5renCg5qp1lrBSX73OcEDGmn9H9QuX4QymOyMVCR2oO+DjNgHu5MBmORUVTVixjN
psW7gEN0kK5pcBZvZ15gTiCLOQTRfia5apizvaShiG5WqG90PT7Bpb8Ya4FKhkjV
3ausCbv/HLawrQojbV+jURHDIVjeaL/EmMWoS4rVTAzSvfFKSL9Esqo1tPazCmqR
t8nr6CK2RHwgSUOWqWK62eHJ7uAvMwYNzKgRpFoFPX2FSL8W7/twwL4mb5K9KzRq
L9XGqkpbcVyP+i9Bg9K6YAcVjl/OwGuMTgj/QYZh7x5c2U3x1eFXmesahvWLnN/u
dcGCGYqXq6yYQ9IPMASZJd4NPrkJvU++q4X4fElmMHQqK/Mv58pqF5odO5UBgVcG
GhihjCik5L5EtmojSeR5KNLgdePnr+oCw/6pf2bAx1X9jdz5zdeMuqWH5D7jzTJX
eTxCdhkTxzfdT3/ZCr6KKcLOOnmlLe5s0wdMTnttc+TAOSVLE7mUcOmMwOp/jPkB
oQu/LqUHAEyRN9mklkVAc3VonNWte/xbFbhJl3gNBHj0FCf8w3+q1s3rHJOdTuuM
bwXB7+yYUPsUcGRXJbStRWst3d2rYQF7uKcd9lKSlIFmuvgObsQ+ri/flfZBFc1I
rPxFO8GM2bHnJ+oOJ9vcRJKnOPcyNouj+I0we7q+bljp8AnQhlL5Fay8kk5Zu3H8
qlUk2RKO0Jr0LSnyvYQIpQ1KYR25aKIC3xfBhmlYv2BOLE91+O28VSXHWcH5i6fF
yg8BEn9zHU67XwRw9W5XWLKXYxgx0f6D5wh3CcNnNHBXKjvdLxclzDI2zpPNnE3p
F/EtFd94/LlFZwxuFZaJ8g9/YIfZI3HCYP+plciOOBGvoZBMd6ccTlTw3DmImNR9
RbQOvfBSQZny1Nipih8bNpuWCFlgh4v2q+7xu/x2Yy3KSmKmfC85nN0EKWQiFQA9
kTMTwGhPo2na4aApWsO8d7ncWaSgGO58a+yLCIqK7+LVkonLtvwgjU8/3T9tNep4
QVNsQN40AAED6JZUyZ+emmoznTEPFCECGYMZj2u86CIt2xxqbhiYGgSLzJvwPBtt
v1MwC23iXLgHh/eEBf9oDvtHiXZ8E6orwNaCJpquvIDe8syA/Tg851ZKxKZSg1BN
104+ZriKg5hZ2MwqhhIs92ptEm4aZw11q1LXcahNB6cZaoBQ6skgXOAMfzmWi8am
Fcw3yqyDdyEv9yfAcXl+giICwhFzX0xqJmsqPdgS38Iq1dfVMAQtFFv02kqMtDNH
1K0kInI5bIVBhoC+L6Rf/r1u4S4Cul+1rnQHrWFzafKfo7fIlTzX7tMo+rLx/umn
XeOHEuItaamhX3FZ7GC5W8JoVWezz/vAHHV7QFf8+VXjkscYwAjC+wMNfIMNpvmb
r8C712AaVT+nu4E4Q0gN5i2OMQe/NTIGHiiUOWaTM5yZAu/BS4n9BkyeUfnbVkhG
HwXJ9lqtWHW3DeUBzU/CCLEz/CT3PbEoeIbxSWI35O22IT9XBFf7BLBtu6ZDCX4+
XFKijtG8ysSZCmKd5xyNWJFeHi/2S/AGqvUjkVXcK+m4JIEy61CQ9o2Gw1EJNZGf
lO9y/P3QTkuOjm1g/XQH6t+CZeV6AuooSPkgCP3wmVLmvnr5WDmcsLCCDCCSoqe2
nyCOnNvIqV/T+FGFzuVVWNLCdINUMT8Uv0XQXdVNmlA9SlCwKoDbEyZbpnZqK2xm
ALgnlzEI0OOCp9n4PnTlv5C+r+8+I3HPOkADL/7/4p5Yvp+468DapjrldhcJHVqS
MwEFo+TvEVQFiIlm/+9EI6USUBbwoU1lKI8tp4kK7JWk1kn7GLZZ0s0K/YBfYCF0
XJ3b8c+vZiVp0T4+fM+p2g/nFlZ7mddi+bQnj+2xn4GSjm8cMpe+Dwktt6zWv0pu
OCO5IWt7VivC0PEwVe6i4dsCB60n36un2kUcQZC20Y8voG9aE68LwCJDQOy847/G
DL3egqgx6lPbabpohAsiCnwaHLfHWy/3PG615fr2NJvBVdz5DqoWcNSmZCmIX9kd
cMqtmdPttVV2d6UkRhomhG6T/b/6hieWS5o+Pqv4LAMzQz3vfPvROeb6C0GGpmqi
sSMar684LtM44VZk7b4m3amkZjCFzMUPPN4SUQj6lzeqEPfiiJZ1im4Faknjhsxq
dAlyJBpI5LwO82CRpNQKdvBKRW3jfAvx4KiaSrSWguNczAeHQZ0FSpmBHCC/6HuA
zRzwdyagJj/sWjo5NYKVOaVu8bgV5eGOH1TJayyoAnlhYF5g3AO4/e11fymEevWP
l3ZmOz28eItWaKIY1+an0CgzpmlJ9jsVuD23i+Fe8MiFB6cO6dfZhJEO1almk7Gb
+46ZBwTEe5LQECCCAnk1uG1Wx4HSJy6JNRlBgRofLnVsRV/lp7NrQFQCRp3MVScT
vEensG4lq0mqmO8nlqQNmclwvYiZqsBveaDiCsiztvPutF2fxmdoHF19hjb4InTG
TjjKPl7IMbZt4SB4WghQiub+uJsxG0A7ZqMMjfoqDK5kzInK0TmBhhjBCE70Y0h4
NLa/FfDyXaxxaG4c76H6foDZpF4jhVtkElxgwF9Zd+1BpguX4a3O84mn6/FLLstA
OIFAYjgVtNXBQi0TJmdAEEaL78SSjon2PDgBFxwm94sLJcSz214jx+2js1g9j+DI
BS4Oc2t/xbXpf56XbbX2sQMkOAc6SZv956Ie4C3hnt5PARALbzphgFKH+XCH9K0m
dcOkSaez2IfgRJmeRIhmefYJFxTS8cViBuObTCY59bQ6K+1/sNsu/m4Z519TadWp
81EoHW3eiwLOqJwwQsuUHLPRmzkONBekLhVd1YsaNBTqDDl2GZqIf0g2v8qtfoNL
KiznFWRHt3/FRrIhsEhjpCh5UnaohyXhYKZrX1/e2QXuOFM0jv31jFKbWkRFOP3a
Hih55YY3Ov8uIfAJA7Y1kixQyh/PqZ0tMgc5663MBnoWCjt59ncLv2bR86RxL1Hh
5NouATZ4fzvSTx8bCKO0bp2Oc7kXAnE6lP5Knt3mFaTpA2KTsRMngO0o8C+MrD3W
b5T11F/CkM0E6qBGBnMq491yluA/hYZz810RbUcJ9M+yj5TA36Fa8HC2kPcs5+O6
qilEiBcQHbX/j8fI1cansPQ+8JpbAhRnAszo3CtkKYKF/vuY4d2l77bfIVzOCscb
m7BAqZuROJxVCwjGDr28e2ytSDWmJ8Jte/P43rUJgOI92pQCFMvvO9Qc3rtfx8ED
T74kDMUYJsuvyP1BbQSphJFMFICGAmtcr6oimSa61Jn/YxW1e8l0NOmSAMWw4MYX
yga3yAhadJlO0lqfOGWMzDfNkrqEa21F4mmp3Jg3yHgfrkREriSP3SqDHscZ3nZm
XvZixE20FHWFzRDKQXZwjzTfg20/LD/Sn+zyS3rPeceyMw1r2/4yZb1QeXrJt2uA
duQuOECfnNTU04qZ03qnWuIsj+1GFqtnjX9qnBvK7Q1BMui1GXpdiaxdTK46AOc8
wjFC3SK/Yi4gv/b82ixeonUD6FPCaFbnrQ4LCavWIiQffo3R5QTE+17E2cRrdsb7
pHCZnkHPe5ezqBUNRo+Ren3rDq0zpGsIKubLG/0yuhUtxlcEY1UzEE/zZdzthMyx
H5wy/FH/Z/0AGFARjreF6Wk+1uzlCM1ey1JTHgp0lMl0f3bwZm7tQOe0HM3p+djT
IXSgtusFv3HTENc16rEP+suWqrQ3gr9tIvhnlbLJS1a0sKJlKLg+yWdb3hu+0DWy
esc58GxcKWAh3hPt0J38ZMZTkNIsC6pWm4C4JiXwioEzIC8bJB2wT3Ny7b46yfMS
FApHTQR4hJZWEp3KztcreWlh6agZbXMJgMmfeZsg7ymhOlggXsS5ryuHh8WCRPYW
SfQ5XXtFkyQZfv9B/p8o8qGBNynvfpYb5WyOePqRs1hvcpUSZB2d2ZTUhdOgKdF6
SPP3nFJA1b8wH5lIXjRcV4WTm1Z2jxQZtqwLeW4QgYZhehTRroeUnxmBbZuL/zmj
TUXBC7nHB7DTUvCTaDs5F4p7IaxD9YZopB5304kWLzfp8KOB8REOVGM7MoXya4kJ
u0+CEBjWL+voQmRhwyqp4AGNHYIjfeofjEfGsFRCkOPWGoeLKX8yNllCektwvhlp
WJCL5rUU/JmJ42oecS1XtSuiD8Z1le53jIN3Kj+/DeVckcm7X/gSTxTkj8jG+mxJ
BVG0PI3u8hnRvGqiJseLkAfdpeIafj6Uc3MJmaZixfKpqaB5HSeuIqecqqs2qwZK
DI86Eh16XFTM51xsiFpaor9y/qRXjAtp3U7k9dxKNTCCyNCpdi2QVcnva3/LcWiE
Mea3J41xW5jzMJx26Zg65RAJJ1VUmgkjiLUEI0c8kfyrJ9Jk2LeZHsSwwiPq9x5A
qd4zKTirLqTdfSYLiFoh3BhHyhHnGp97jmMWaYrYV+UfxdxeenewmWvuF6tbi7rO
3V94iF+8iuPNX2ZFJMMePKJGpqStX92BdhdNxAqznTsku67mkdtnNXt9H3R2Qp9w
rBDGmB7QABNd6UiDBdhwVIGF/eJ5omaGQNwJkrfDVmGBvOPGgcSthyllAEJoIcY4
3n4TZhR5rPARsyIBUXubcB1N1XEuUFEsSANriab2uj2FnDPezXIDQlaFkT+hpjJu
sTE+WaEICr0qSkhX9bk5AuyUMEqHSmRcUWy1kVEWEiUxugq50cszAaGuH3EtLBAT
c/jckmdfOvA2GkqOF6XzZ2brO6B5owqU1oczFxW/pIhyyIpPsm5VOyvq+mieNjPY
DreEFkIsGeBQqLztHiPsIfl1T0ezjR4Z5c81pYK6jaOrT9bxzhtzjFk2cYx3aoUc
dNUSgWONCNGkMAMBu5Hfy8KUHX/T0Jk72c+pCxqaEmz/Br4sd2MT8A5qXNtV/wc/
TyfkVaDtyk3mZCI1Iw4tkFJ8mjxOFdkAXeKAYSqM5I/fGUjRf19dtLx2cze1wIfR
HL/Da0opBw84ADwOcgICZaOamOJYoh7yh+E9Lg14UYMg5lKELJHq9fcTF/6vvH6v
0gMsDZRX+c3Wa3khZIlbpW9ohSXvoPdZGdo8OLJS8Ou0Yb8eiZnVlsdRXHwnjaa1
7dEjfvqIeJuNb4d4fnhoeKtXJGzp9t8T6KKIsG1eIR8bM6RQGVO4jX4U6H4+9GQv
muxsd+crsNhh1mthw2ore/7wP4RmsOrtlU9Iw/lsrU91tTI0iUGPEowcHiuWJQlt
Nc1MASr2Rwuimda2Qy2SrAtJWQRyF6q/cTF+sHEQg5GXcy0sh3+6vPs1lu+E+xvQ
so1scF0VilvP5w63dN031JyiPkwmVhrY7cMfiwTL0Qr41rfEgZbZaybDvi1RK+29
N/iBIqhcO0BoNiHf+J1FXCv8T5XtJfMIB/H79AsSZXkzSxFzh1X79NTtiavAJrpJ
aQWpKU3xaZs2Gt0co2PV1om2Vi5UzOU7qJ4OyWR4ciMMK3r3mCEWbk4gOC135nws
htLl66Mr5kxAB/TFiuTwRCmQG0m5TmSl4TW2eb4oEVjrL3rO/Q/PabJcbE1okfnU
dKrbry4iCUY091hJbv7NCdpWv2u0TLSg7JLuxcf1tfmKerK2GN2QzMCS+NGqyEqB
tMzpiJchnExvOMqSCddtrvSdjPSiyhmUgf2cisU44286LO6oXabiqNnxwy7jGILZ
6kD997KGoTdxULvWqjToG4PVtIl8zD7QhNtKXT1xTeNcKyBh4dr0UkHXbRmZ1xn5
gHfmckruuPwI7E1kZKN41DHNoO94s60McO5YiC77juAXHWD7cTudfqCyKMGsnBhE
PXIL0rSr7R2TU0wkg9u+hyginExBmAJPnOOk5X6bosEWprZGgWWomMeT4t9IUE0W
O3RClpRara1OkWWHdWfiZdTc3fa9UqlWu11uOSHbrmCvHyVjRH/Lm1sNbuoDpI4e
Apz2MXznAVqzodldzae4epkTYCdYTXDqXvU0HfgUUOckyQ3qW6mykZFFgzXu2n6p
NZmAb3NEhZ6q0P5SOjwuWKKtfKS7oOJbxFz/XOeCv+B0gOzdYJJWi5JNTwc/hvkX
QSzyWr308awMGXmIU1uo/suPMsf6JjMJ/L0bnuJFNyB/ppUByVKOHY5esiU82/0P
tRLhP3/tk5I6bCpQPQyO9nGAkybZkK7uzqhJJPicz2lGVcbHnnnQxEtRbISSQNUe
WOTbe/M6p79UmtSolbDJYDrYBG0vvRq3mdUBcMyAbQq8HoP2sfoGgPrgnv/ez/8r
k2U9SncxrWTfZYK2pLupdkXez0jRNBVbXKXZAlOF02FE6rhbHjdt02wZ1kNZeLhu
68tl29TdWQza3GCr4oygbGC8CXrmM4d2jv8SOKwWz0/WMGSVvXhDZcmY4hDtdpDV
hjtzlOI1Y3kDsDKuZv4kJR060dS/gSLcbwUApC2HwTYWpQ1PFUW9hOo+JoP8FX0A
1ioCw1C2RfmviAQViGB242E89GmBiKHLNUDeL+fbiDkpfdpNwiCudQjV6cGPtVmZ
v4Nwa/znHVESNc94H8sVjJ+nt/SwBPaiV1FE47xKHE5hq4HPEIaHlWLPi+yqXbqO
mxJ+p9+XOoW2oJqCgOxx1iqItrn8nDfIFAtZkx2YYORz8JfMDdclFfqvhHR3S7ab
aAInq/ei7xzk6zsFdRRPfHsatjtKb9JfF+oxYC+Wtv63RXdejmTwi4nVwFnkbzN+
jmA2X3DJcX2XV97El93sSl/XZVahPOWIK8x3Qbd8gTF5Bo/lzJC7uuyhTg3z548Y
oVQc5EoMrAj5VCLogmwvMKZJebNHEJKps6tLPLlAiru8rvXUyp8+cFmh3BC5L6iu
TXMQwRI5k80XyWrtlwP2L/my7BnK8flsLKF5oDZEBgMvcm24cw/NtF+qxafCJ1d5
dH5m+x/OYyA0+3/r2yZWM0IHiCGifSoo9NrWzmRJl50h44kZzm8vRSdmolf0NThn
9U1uLDCHKECeZCXipkjQ4R544cWZOuQonGcsLFa4zFEVFCKTibZS1A6W6xLNYD6g
YnQnHVQwfPQL1hfdLV+IaNSQFGC2iuHSwj8zvF/qSNTDtVSMdPn56O3jsn6IE1f9
MMpSIHP5xUbmh87Bxuy5ui9i2Z/1uehO+Q4ITSHxdTnJtvfXZwnyRGQ7iVVmbZ47
TsrqH/R4xlhe/Z33DZmEcN2XdTwtCMMQzxxXy1ajngQURnQ/r3E6N+Kuuh4IoW3V
zffOtr/qWX/leM+HHxVnzLhHlhJzvFshlgMotATU95SNX4S8xhXwTIBZ7GD45310
CP8TkRGln+zOy1aQEAq5Z6saC0dZnByAk/+9XWj8xGs+ccni7Sv63RIynQJHfeVV
CIk4qJlAvJTdRlIVIDpuO6KpCBl9ApjAV+uqJgKaPCXNO7adzZQlahpeDoPq4JtE
JSv3VqByIx1d8wLHutsMgb6c+fzvUW4OMyj5+HwBRc/vbdFgb+VnuH6yDkSPDsGH
Z9B/neLewz+4/iBFPTwbpxsUmPT+n+bSJOk+MA4oy1unIfqSy9FIRFfd6aDMUyni
ssSWbD9FW3P/yZE4OlndSnq1DZ7gOWKtTr3HsNCCSO6BR13hR54I12Vl2QZdOkAk
ykT/TEG6Vla/2mrZc/dYTedf3TpsW8OAGp4QO8dagZT6dytUfcFlePw/F9VzKXe1
BNt4zbfWwG9GcK4MtKQRuOFgjuz/Rtz83PMGbGm+/huw3AzOo1yMHzIfTogguKlM
KZplY3APAgW1RIYXLF5fAngTbJtUF2iqYqFzOrXxNOOxz0iYxVOBDhZAp22dA9M8
LhLvAOBM+WQAtYctvHx1wujM/+NleBuhgdoILHy9B+qzd9eGXtRwaqlOy+X/H0fy
crpGz7SqZXj7PtWsL6k5X486G+74LPr3VfmgfCn1z4EsbWhBTsmvr/9jW//NRm3M
fCM3OmNv3ZbV+NxdiNBgnbL+PgkHbn2Poryz4ORbcwCKf7fSlsOx1aBT8tLuIlrW
+Mt8JulTXvtdXvSihwaQ8PrIQLHbIW9ojuK/3vXPX/0EWM3GuUzUrU8KlroxnQFU
IDYbZ7xYLPquvG6VIAvILPqod7WHB5/ZKxzNWH40JrCaYmfXhakaXR3IG4qa11vR
5G1EMBOoNOand+UjIkT4uQAVPA5ztYttLXzFI07ulznd6I1MKByxnefvmoGPVIOg
8fUTPFV9uQ/K8QRQ3dvKmMS/nUi3VSdGuVA+sHuSyxGlrwxA0au3Dn1R3wgnVFXl
bqSnUqAF9Le0ZGz7vZGUM2wi6DcvlLfxDEyeQV2rcCOy0iYe8LTaAkAm1k7r8pWR
A6PytXq1HjwM/+eSpfekPuCeoEWWePKe+wj5/47zXFDS5h13ZaSiUJbNqMXdvH4v
+YpFaNKEMqEvGHbXlpQjd52qBSf9JHr5e0AyRBPMJtRl71qLYCdOwleTezGzX8ZL
QvRAB+H5RRM6vFT30u5MZi8QOF/pp5Nbe1EHNHM1E5T4GogYRbzOBZF0Ei8DbfWc
j67EZBgcH5qSTvdzmTDH/Ao/ZD2N1zzGyzA4CmzvC7jSWKUOahUCgv4zje4kQMh9
8w5Ejvo6Igys1SJtFLbzbRByziIfqZPkTmTiqOay+L1r9qF1cRo4behhNYl5///2
Qrz/dnuNhN0Ax7tho8WXI7UqNdZASibOaBd2T34qw/eFF72F0HtBI3dJHoPr5rsl
8BnGE6D07NwJ7l/rwdisoKFn67pqhNyyX9WFV1oHqO1cUOjo4F+JZZlypX3JhDBP
n8+UUSxY07FUrhaPaQtbE552k6W/3wlES0DP3/BbFLhuFGOJkA1Zjuz3rzpee4CI
NHoZZxroPbfaLRNA1eymapjuM1mBxhfSNldNk/liAIQ/ELoiKDfi8Mexw+l3Zxec
Y+jyLtbPf3EneIpEx1mZVngIMCzOMGitqJADW9lCi7aS7ZpZVnvTc3Ger/PFn/8u
Oouz2KUI6bXsgoWpvd3MdMB/32NyOBd4AjIOElS4G7yPs5oB+OhZLussrmB6XxlM
2PI7Qs7Xd7U6UyYVX2SNZCQnZSTMG7DwBQd9CLUpLn6bYUcwLPwz8JbmmrBh1vW7
HvwOEgVv6sCogPq85eVXOHOrWImKPfQU/GKebI/x1eL6lcTC4bRvqjbZqupV5TMr
AK913u8hRPDe7ZEsFF4qyeGJb21nvt5HQU2p8uwkwe/M8oztSJoGgH8AIVEPrNjg
ryeDaTpyAnNXf1dnIkBfpz/8IkxbF476lvaip10v51f5mU3mXfKnPl0ryhA6tWJB
aZ0J86FpxZFfKfIzlkKPaGfpoGtCAvevxFKX7uPN9BYBgDZwSvTvugFIj1CUe8ja
8ybSkhd9t0eS4xKaQi/5eB+0rDZmDQ4jzS3WRxU463KGm7XsccAr6VyWaFaZlLeJ
jAMp6CxbJW3OwKOcV5mDqkP/fw+N0d8Dy2U2mqZgezt2ANmV8zxHdUY8QE3q4coN
dVeyqvjCIktYIm5ODhTQ4JZpNcC7IbG6VAEjBHn+QGWWFaMWXF/+aV0Y3Dl6ilu0
cyg7LbTiGCKWqGPqv3mtpFkonpYikAoosMX93psnLMzPBv5c0irjqWmNdwMKNlRv
i4dKecWmYzADHuCIu4XltzwEcPVgINmy1uxxFaaYfffpCt0ffzMqjE/kLLHYT0Ee
iH5xJhHoip0hFIz9h31JoiWePXAiZkIYGMRsWz3gVaa1pEhBmg8u/b9gu3CDFZ6W
PQCL/U8YZqwSoeKaZZY4xB/9qUdUy0hm7/h0p3dFt3KE90wzgIJUEHiZRJF2RcH8
fMllr3T9zkw7FwymhhJsDqV34xxEKbc+nlo13bs0pLjscEO7YfRvLqF/9/CKxT64
k3PxT8w++wUYJU12caN8ztHt0W0OsvJyTy7dsE4sN4Fe5R4dXA+2ok+G2NqjVoAh
a0dTwr11Urfmnu8M4iuyLYGDZEqjpoeLy5TM99DmN6QkG2lHO8ruXJb4r6omZsLe
5EzH51NdDB77tk7iYuo6q+YsYekyRM70v8CSShQZ8XUwafxK/L3CxEwa2DJz5fHJ
i0dLF/6lba/qt4zP2Odr7l/XMDKHCg0oGsHfP6qGFdbobTEdNf2UTuejArg9tqYO
pvDer3Rg1JF2PCO1MUdsY0NFKV637ZBq/zJYfM0kZ6maqk+7UEnJRtyy4HZ/8snB
s40unpN8vDoc/3e76Y/jQGTkXYsti6m1qAauaQLG+kLMNeIzNKpcUenbNnNO2MtU
0O0oHVgEQ1YwLRK/QFEepqUevG4pQA0mGijcgZfvWN5lMYVrKhiFQUP4kZPeyGwp
EuuHhCYqfUsHh7qdAZT6hd8RcSt5v4506mTI2s28iFQWw9o5D12V0mUFW8PtHdG9
cBbifxcqph0Y1BslOBpGJTIR3+K5sPIC6ZXH7NEhq61yCJqA6iwnJvAuFE1ja2XE
v9wXH3qKYCcRh31unCFUfJS4x3xMlULrC7kWQWBj5IdNLH9kQZbMO9fQTOFBFjMT
yDeHoynRDXZrMZd96sJf01+lrhHliFBjpECDR3l9D5n1YFeEH1RhJQ+/TWO5JQUE
mrZtFaCCh+L3gBb0qHpEj+QrYtBJHNDB5SKjB0hRoVKV4yZbmYupQKr12bp8xast
GLMj3G3p5MBi7U54on/N7cF/MKnrxkaH6bVv1e3DZkzV8Tdlxo6L4FW89DMJUPW2
MzhGyEEn6tOj36ZHP34vXsXGygMXf5bCXiA3qfuyexNjwMow+3xP7fVCzLLRt+18
JaTClIa6u5XfAHmnz9ctX0Dzm8XUBNK1TZgZGDi3n90/MAoxr7hakx0IpCjEaAB7
W0WwiC7hEqGfzhcyU6NNeSCgqWE0tiMH0XBCIdyR6EHQF5hmMUwj4iUBk7NiHtWK
rE8H/qb5CYDskPImBx4I7y3MCqSw/OjNuFvLdvE3nL4B9IN4SM2E5sR0x3futBXU
MZDjApRfQRDBMAXqtsMWp6G2bUfCsbLuURFrowahOGfbCQtPrNwMBXrk6U+QizRl
WuAEoKN+KpnCZ6idK6u3iX1Uahu4MP026q+7ru1ZrsjSFYo1PE/S5+Z2BpsoKF2K
5RvkQkf8f4DDqG69bD81zTlgW/5JKbKTjaultxT4244bqhu9MwiMHUesEHej3tfT
V1IP5fMawSlXumvyw0HZBy/P0vMA4L4lAJFT0g8E2o8mTJVK6I4vUxOI2JeMpFuL
f5cKbPgKrLiDQ6e3NrXU3vmGV05eJJIo1tRVnpaRVT51SqcebSmLS5Kg3CBFPsjz
U2IgHWh4P1To6bVrOwvjHkCxBUYeWERaSF7SEZzXtz6cLto5OxE46VZmHbunry8s
teftQbL5QCW6LexdXlsTvOyhzjlH+9VeCrTGSNl7hfP9TtdwDQZarDL3esOOE/10
P0SL3fSglstQv1J9EZrfTd4N2cL8/LbkV3jf3KaJwOZGFb6Tk8tPONBkmtzD6R2t
NBv6K7wSiag2/gwmiZZ2W/vovWFkU5ETYqD4kgo0FQZph6vGETw09Bfyf3PesjaH
CnhR2HSR80gZOX2ROKZiaDPUWnUZ5yAAdf6NQGpR0DI5NZU30GPfJyJKMmPOg0vV
5lLNScWYR+wpVhNAnCn/DUqt+8zfmut4IvUqLW04hguevcbWDSZzFIqPBvm9oO3i
1zNk1pbWZEk1Bso15JOUUhuDjtBuU7Pip+XVHonfm5Clu5Tkv3LU7fVrPsUGhhR8
K1r2/TbFMLhBuXfMc+7lbPMZNGC6SRapvoPn3GYr487YTojNKdf/aIR/NVkFD2Yt
HeAWw6LjvA2M4FQWBxWGBP4lVfcKbIUthnqTCOp+6QkZHc120DLFY6Jfs5VEUBg6
y/qzhf7aSszLIw2ol64+2T3zrFkQDFti3SaOX5JEQtKAGQ5KQJ7pTg6En/Vuki7K
Gv/Of/7FVOxSejoWTh01HR8oynK+KKlqrlkRalUUL79av75tFBx/pTL5dzemzpo5
pJuGNmhx92PCjDugcqO/1fepMWfg0g8jLXzuvAxApTglIWkDOrFqSnyXHLgzGVtu
P9bxjKeYDGgi3X4dBOO4X/AHuyEeYWB/cphY/SiYGlDL2zH9lema6jwZCvJA8uwE
O6yTzk0FD9X/W7HTPC+M1Uq9GrHchcg5Ke1ylkuBOKAK2nBOq6DPttmlxbgSobke
4/zOkM16ChfJ32PAUB4ri5ega2TtPGkt3rLI6Sz+cEwyaUMSxalxo5gjtJTrpoxC
eRbSSyvSy6M35w+L4IPN3enw9GrRkjewXBerE/QSHL+tubm9O4Q4jDzw0S6d5gle
Ml3liEES6d79LExD92WJMyFf94NAUUR6SOQY6rxpK/6KjqiPX8ZDsi40BMZwF6LP
dvhB0VBR5X7jujR0BdWFeA/7lj1NOO+qZz5jdqm5eaxZ2PxmDW6SykPfzjjyqiAA
B3uUYiWJayOFaXMXZRv2b75R+9aHhzr2wN4z3VSp+UCF+lqowgq+DiJES+aR4ixO
kVQ1l69r/Aa0Tx2KsxmrMeSkYE/8J0D+LWHe0SxCS5g2XQ1jfmtO0o9zi7HHfa5Z
T8ehsI2GwibUdl4qhHNs7DEaBe978vT58Hj8PW1nQrDyCPbvdHpYXLVZ4Ctc8N/D
VtHEyrT9Sa6FmYnQDxGImUDlxYn4qt24xP6Akb++WNJxWHIhuDcDxYMW6j7bxiMM
bZQtV2ZXIYPJXizzSGcp8ZC1p2+RwPEZ1+Z8JGoIIDsBnfwhniFtJoQGSQnH27F4
jAgr+wdOTwvYSuW8X1bluqvG6C84+i5m7kq5t+rknD1QWhNCatfN7NZJj8wc0efx
yPba4gGgrDvsqdCl1HN90WkJo31R/wIK8NWkb6oZQoiWW3YNK2u2rjEHXnloNhJk
wEv55L4Pon/N4iPStVQlEQ5D/xDktkr5GNkm1B03+cQ8dbxzlwR+9mN9qo+MjADb
dsb8ckL5W5PHfNbzCydftEgLbtEPljL2SwbshNZ8I3BLtDAQqD0oqlXl2fy18wSf
45pbbAH5jcx1z1kiIfDr00wIOARaS5MKJVpihLnikMWGVWHLgqgywJ89RtbxENN1
rJwueeQqnJj1p+Nk98FrpyuzLIGvCBjVera1jH2ZFEsJSvEl6Sg7+qXS1hERLAzO
P0UxKm6SCH2RgJiSagDA23C6F7UVv6TegZQ+lKQg3CooqitQ0KDRV4HXvnGd7g5b
XjGbjxV+DW7Dgww0TfKe/c+yUDqKJSxxg2TkjVChQ4E35Jg0qkoJY8lpM+GANWSp
EBCqst+k56aIRuLt1BwPJKxw06XoPrRsJCNnfeO/7Y3MJaK59xYi92a7bxcwMic5
MRYpuqs1CtRh70hSrXFOMfCkcg64LLkl+Ec0Z7JRLgwW/EZB88QqPbcctV2BEpXF
VIshnHQLEjaeUrCK0l4v7ZWvOZAAxnnckOtPYcxT9bXmiMs1oZxRqb2bQb8WJmno
rEm9dsGvSeXxP07oZYJ4Rs6EMk7ILF9esB+nn9OIazdOGgRYx/laaQPk2m2wTER3
fOSZLFS1EW+jesUTBtnKfrljawN1YoEx/4uMJQnv6mUWnaYQfrN4mdi3u0N3LwVA
N23S5IXlvaQ4/py1qXkKT4ecWX7bWDz8/2lwVv+ydIIt3OUuHa6JZJgnT2CK9GjS
Dq7RrHgL8LlKRd16iNX/F3Aj/itPVh4rPvq2rhOXXXYKPhjGUNs8q7N7WulZfm+E
+LyyhUhA4nHRtDQCGh0i9wIbTEzTCW/ICSpx/zEtNU+G1aVnu7Plzjz91gfVNdY0
I3NCQvFI25R5K06WuJEwUQt6KrK9AW88tMPL7txZyV7AfxkmrOHHew9CbgwP+xQm
wrOXfA1ic38L4egsTaoskYLKQTCFXzZmgYGGcvjNVSYekWMYadFCMTyX1fzEG+co
i6rafGN7zibih7AOg/giDZ3yx3UMiPR86Ep/J+BvzhTb4VjPVwzayPZ3IVgPV3Z4
zfSM6il2gTh+6fJoq9S7DghKHYmsBOAHtsW4CsfMlk+Orzi63u2O+zSdlAXk6sN7
mAoYitN2ZP7kP0J8UJ6ucfk3M6tzonI+PDi5b8oXZhrIR+8FDGlItJm7dK2mCs1O
lZV6XAR9Dk/M38baYwDwoDZ4ySSYqMMhYCWxaHJ/tuZcjLFA/UR8zUL7Bqf593ZZ
2vvM6XedQ8YISk7K+XeU0Tdw+Xb12djgGRowTOs8bS8WKJNbQ5qi1fzk+4WpS0m9
OzuoUZuaw3xrdkXbD6qKiDmDs1aaJ5hBK32fX9Yugx11AbmDS/7eLUtwCTcEpMbb
XsZcVbRbkH6GV3MLdhe7am93WhUs4BAh65dvjx1K6qjqWiZhJt+rwzksEFVLqyB5
G+EojWGmqD+3eq2igbNorVo/i5cfD4urXPrIfclTV9yvuhHjPIAMBsjL+ZhjMc0B
sEB59CLwtSe6V01LJB6Rds3pjfLcUZzmw9Sxw8/mtqAdXg9qQloL26ud3a0V8Zcy
qbs2dZsqkxxqE/SC72rEz1Ahr0+dT4mB/HvOLVNyv6LrHTO3dff+/IxLyfW+IrJg
w3sRpmpYA2t6vzpfTcuWECHiOza6A2+qMSVbnzeUMEijjc4QkRK4nRsx9K1V/ej7
DjZrsghDCbuoGYcdHIxEd7B6h6sjfeWp0Zt1L0adKLA4LxTUYP4+1CB7bwP+6cjM
6+zmwArPmv9Hi3zthfcOEsyD1lqqz4/pgmlbCHKYvV5sYeUC9rwrEs1LR0shHmTG
6yTikL5tr9aqeZ1GKIu/FdRG/PdKgCbt59mtQP+eFQMV4qfbp+kf+w37sLNtEruH
r1l67HedSOYWzXxVjUVM3JzVbEQrvVVtJGknrpGAAbIGmhzw0fbyNxg3uq/A7GHl
v5GGaa1EalgpUPCtP520/n0kDMLB89y6WZs7FYxAXd2gyFnMuTu9pS1Ya9H/1m1I
I5wFccopXtZnKwYTQqI0wBlMfIX6S95Oz/p6N1EdoiNBIA14H25ZUP+mvAb8vt2I
YA9g8qKbkC0N/BFllRueC0UuFq1Tuzn1IfA1p28Wf4Tcqe1KL/sc7rYOjaw0dH5U
6HHh7z1wf6XP1jOGh6Icq5mWvUJbwdN+dKvK/A+acbYb9UTkCTxBMA5mH2MQ8V4B
kWhvu7p6IOXoEMJG/ZcgWa1KxI2BLR+Su8LC4uy3A1dNtvTYfd7WZIcD0F60JVL+
qaxHdckOPHPmOLF0oUX8wZoHoiRDgZMQFpvFvkUABG5naqXuInoHubaj2bH96jWv
t69KbKsxguwmtG8WTrnkbMuWtjwHlcA5kvDTf4+atgqTW+8Dw111wqBavLXdR7W5
vP2aGe5qV3tZSIbWKUR5LD+DHskDqstvdbWQBVkmYZ1cSvNtEG3ZdLcXqi01Wh6z
68BDBFA9tRbu3HHIIYQzWbtC8aU7Rd14+ATCO+id58O/+how9p07bI0nawtiXhud
dEydmzq5sx3ncF8Ki5tXSmQZbDH4oOt3vAS8Ju2ghs11byRdX9RTmA4JmUYAZjDL
Dz1GQFFbOP3PronlID31Qc8w27O8g/IDHXX/C4KygQC4zKbTWXm5ByH3Ks4mWUS1
ZLPpAzDlS4mcbrZGLhLb6bVLzu784gkdRxFaW+URIctpHdoyFxzbhZc1iMr1uWrT
+hi3S0/HM1hCyVvVs4mGM/CMETgu0uHFdt36SPLPDZZ1ts6jzidXrQiFYh8zjFZr
neC/D6ogTlUJPtrwSnrj8Dp/YYgHYaIr0EWkPBZzRq2eGQ/pwmVYaqlBq4/sekT1
iAbEXy7XVrQSRC6OxcH4Yh3djmUAAodPSpB9nUPeVlBu2WqVgXj11EyZHPdruXtR
mhmWBk0+xSmns+OQEvQQJ85VMkY6mGGujNBhFE17jn5YYGgouuhiyUxfyln30d3o
lKDSj1rNMSQDFzBKZQYCZ8rddp5qwGV1A+X90KEFtrg8qX8sKpypl2bdAYSWNnIC
t7bnICahP8q010MIOzO4LOcCPehJ471QeSO2kNzK2FW+ZJ0dA7ZaAmflWftDf6Ha
59gGqH9+dcjHlCNHvhaKviadBt5cBUSLfMj9dzesM0d7t6uDrVsuMj6tFwgO7YVF
JoYjNpuvsO8IbPqlic+EHXr0nwJgKd2jxrzVqnhe4sjAea1rrWqTaCOv6p8jTq2j
+UBmu4BYJ85THLQ42mb8gmIhSLWJ1hrf+d8cpJ2mSFCZdfKMRIZRvitfqpzdTQ6P
yQt90b8pZ0zlRzeYgRQ/aJe2mSNmADUT88+8vhnW2dFOPfeaOU9cHAlzaMDKeI0O
q/xlNuYIzsHAgkyJMTvnY4XzGKAylEkGxP3HnAjglc6KfylXSgny0x/JG9q3u06d
EpTekh+Qrs+cmHzdBp8YpCP1pQFUcs2EUyhh+igKpPJKnP/AnKbmEAclvZnyP6lz
Z4G0iWRn8c3gK/hAvcyN3/mff8330qN1f6fRU5POQlp86jUU8Mjfe6WegqINS2BL
L3TD46qz0vlCIhwMERxhlvHcPA1ZwC/NM7IAC5Y1O4qI/DaXmm82OsgKfCjRLDQX
xRx4y7GbRhq1PV780x2Az0bfSpzaf7trUA1hPG407R+9fq+K1JI7IXzXYyduzBuc
OsLkuJY6zt83Dqpyy20IHSzpPiyr7CyAaEL9AMqOTCV6VpSRwVY1Y9yb0wKqs2nN
cvpw0ADwvga/MhxhLhgvE6yMFVIagSci8ZIUpK16JKshwHoF3U4+wSBU7FjnLDYR
e+l8LFSKgEJT4xh0Ii5bMXKiceqIVVekO+PGnWI21aTsQAROk91vPR81KUc65IHp
h3OH6907d7im6REQfyABa4RL/13SVSOBh4y3w9/bMN6l1We70/YK0Jrq+VZwygUo
w355GDg/XasUC1Z353VR/5n1jxZ/pD09cOoYwryyTbSpNh0ib1Lc3wxj5PGosogg
s566R0Z2J6ZMF4z1B/5guXXtpzOm5lBfOa9jQsRsQUCxFm1XCS4eQ+a+7gz0B41J
f9dWajSDHdFLQNu7v/+hd1cxgD0zz5xwQ8Bw3k7ZC1Tab2ix1GFrQgTn78VXPNWx
h0vWYePC64ycw9sPBy/5+s2C4b/Zp6Elhclj6qg70pbhYfGoTXgC+YTZ/ud/7I5K
XgojrnIiN89YNV2X1LzgWBkFrP3/WtzgG7L0NHM7f3OQTDXnMwoFD/QO2Jr5BWIr
MTaWY3XZE/HnD0hduqBmEQPHTb1TJr1VJ1YKyTHZ8AL7ZEcfY7WA0h4qRaF3FOek
FiYXamYTz2q+IQyD3jrhVza+MtYmyxqCCeliz95aRuCj+tLuVX3b3UzcVdb0Lede
cFRFMSaM2IhB2RVxBdPy7WpH+9NnqKCKNGbfL2qdLB7bMoF1VUmbN3s7XFqyvi0p
eVaI4azKYTdWXQ92KsAgpdy/ejUcb0ENXpyDyi3Zrdk4Mh0hkwoMtgW5gVSBr1cw
Mu04A5VdrMNA9+AnwE/3ebLopkpzxrMry6GYD7OYivZeUj1Yz/nufFGy8TLf/MwR
h4GNwCswc6b3unaAfGZIt02E1X+YHsRKMctWW5sSK8okBupaXEV8tx3BwbRpdT4N
iXVGCdUTFGwFkTM7Hdl8ax4a9MxWe8X+AJoVZmLmoD6xYvNeYITKH41WSTD9KAC1
Q9hsGJt43f6wZPoONFvNgSZkw6+0DzcZN0dwzYPvPbpRL1/kJ+mj3mMEe20E2y9d
KXOGRIY39DXOqfsj9d+vlOFYiZGHmrTihXkhfvvSdui/GT8PLFbjY5VOInhDx2I3
V/mEqCXa3DZ0JL4WdPYXz0ZSNEhxk2wddGlFzj3ORFWbs/y9FEWO/ccn2OZ5XaID
iEoYUuPkUqI6o8XoqmzmBTe/tcUseoZBaC3HmNbQcahUQs/SADVi+Mf+aUCysTpM
GVnk5Dl10a2cwzcM2tsiGU8/FdVyPXvZvYUaOqb5YCA6lG68AnExuyKlAOIp6Sny
DkTjN4UND2YKJEIS49A+NHlt+xDSCWiIpATk3/af3dTMuyfVFuFdVjcOK0I1tSnc
gWYPcMqH180J9Ce0dw0OAC+WCam9RR9YmCGq2ugfpU0mTHbJBPbveZzIjaXhZAn2
ATUgL4PBk4d5QgSqXB8a205bECwZBR5dZ/eb77ea8lKFR3cJ6gT5Wa9vvDaLzrcV
zvI+t2gt7QSZ3XbynHxoGJO/2REhRnYmzjLKJCi/0WbJeUtsxLG8QfBmJerYk3QE
lkHuy98bnU0iHSvQKZqLmvdNJrXuZp13qAjRMnhgN8/k03EvJI2Jlw+olKE2tZX7
PWG/xtDR2E+ZnStDNTySF2qHTSxXNs5B/9AlDlqfK493kANw0Q4IS48PYq3ocDjZ
vUOZaWcpEkVYVwLJPNC9PUuULZhKoAt5hVXSr2BS4ZXQeuquGLxarix+UyYS7tmf
qW8qZUjYE0X039HyfF/+jeCjeB77X5iLioxUv4H5B6/6Vw9dbYK5IoYsQ6+PrmGv
bWFjaL6YYj2NERB8Hk0dCCCGg6j5CigxxNkZgyvQoh0v9+9oTObFJzR0oseNy2f4
hmZAfoQEUHZoUOlsfRt83Mj1BuRz1gsHj9uMMlSrw5EEf1aRPub5CKTEgmyxh2a7
vrSF1Los6p747LOYuioY+LeKW4J29qjbavPC/K/T46BJbh4WHdvbHPuhkT5VrlXl
97hJhn8iYgVI0CNQQ3KSBXshir3eyK0A0VE76UpF0LioLBixeazJYOA8CoYqJBuX
fArCNV2xsK2DH7xJq1t8Ss3lu6tNvXBfydualnsURA0jtZDG+hfSVQ3Mqa3e9S4D
wEVsP3cskQlPIOdlL+lJER2bKi6HOn0Na5ChH66OsPM9fx3SwnFaE0MQsZ56PhX8
0OQzuLiyIlIAkCgHGqaO9M4FSp/PK5JEu3x9+MI9TYhNAvfyQKLb0nk3MN4jFd4v
Me/+pqLhzJbHkK0Vids9WiUuJeZnFyb055C7pxqHnNk2+PmPcalYIwjswyR36dO0
RNU+OnYoDVL6bNcJIha36psFhWxJ2QWpy5+rcbEpJABC3bTqQkzU1AM6f0CWgtGX
y1iscqAm2i51JF0Dgvl7V2gz3IPDou8v7Oo8BWacQKEbrHgeWGIifYhWuGAuEJHI
jSKaUosCgSon73jLA52sAPKPrdd13TcYvAr2VdGq9yRxd/xaN/0DHKCMHtbAB24Y
a0Nyai6hpw1oG+6POvrzT2D+x4k6XWXv2R+tCI85DZMD93pJ8NGxwmbner3sZTer
lLyztPL5g0uIpYB3NiXWkuNcZb3WUeNw7QPqmToW7U2B3qmCsD+Ta1DBYa1XeY5m
sX+5hHikyhBbIL1++rQSLb/UCZJqv1YVKBFlhNndFpVljpreuW2Gf6JeYwqSHMHw
hJevJ+PVTGSZliOzX+tY6KeS+bHzRsMX2v3fgfK+ZmHJeCgYWBXM0O6RCR+1cHQf
USMDgrGYF8KDc7NiRF3VxBZC1X8+xVpuzuWxV6gGNZ+BjZyZis+R0WNH/C7q8mcU
AtuuwEhULQ6L/iVSoI4E5k8QMCjFf8Bl4I3+ZL9iSNQd+hQGPH+XBox7Ynlaunh0
f3Kf5293K54gb8ESnRb4wA4yUxZ0wEVE97EBOtWqMGPN9M4WPByJM7/oeAM/tAHV
fifLG7FbAiqpqSqqgBu8T8DLb/9OyTpk8lU4+WPfiytzVoa0iuIyHimsv+24MLIp
Nsx+nk8/hekcZ0vVkzQ2MSNMIruc7r36KkGYh08SLgME2ibH/3bpbL/RKwzS2dda
MukdgKwDYkAKYh9+9Fltah0QaaBGoCEDzZnsjYerGBS1+VnDvdzpSsrxfPXgoFTe
5+sOKryWl7L94rE3TZAnrG+jbfbwf7/5OOSGwEobZdzXmX1gH4gXDtIbn7v3Es61
74cNQ8vNlT9Qwm+nO2vnouvK4W3uGv8hLe3vVikg6klw2EF2RCLeqciI6zGDMtVw
o3mmOIZPvklPYxO+3ziaJGLVjbQX/GHDCWXm7M13PXMrDBopmwwpRPLjzagMmbyH
lusRyFb0ELFxm1OEwb/ly7GBEQydyuNIMwtZzVB35zTB8Ue4Wjsq/HbXwBN6KJS2
7kwzprQS1jex5RjGJxoigBmVydjIlDTbiOfJcsgwyxvt85zOZzrYmWDuo/j/RnSi
ZKpIA45ZtpEb7C9S3xXSLlmiSWwTN9kVLhckmL4DJ3XGpp3aT9WsfEfiKs1DX8RB
lrxj6EmWj4y23te4PjI7WlJpM4w/FcL18dX7JaMX7OCZVP0swvYxfKqPuLpGvY0r
l5Kmx1xwhSJtyDeKzglxMzJcgZSV3ar68/AU45mkh3Qr4/wKbX1CvnlJ3zrrOzbj
1GTNDoX5oBcEWv4VIM+nPAcKPpsFUrFB/NCeQ/SD3fsnDoKVcuqsWIvl72GRxfvS
Z/XPsuBms33vY7iY4hpWlsLaUjLBGGMM6IQ0FdTi18XdwZZ7DYdr1qBmWKI9ualf
V4egJvdPiTCJOMqhMY3j53JtvggtDi/elf98gGAoAcDlQM6qE/mussV5Z7rWIlR5
4s0UUEin05zmpu+Cm9C5CXqQwlCKTpbVx4UT1SF8Cn4LvKjUfkGPygWXoJo9mfSf
d8xGyieIEMciB2+YOrzv12876CXVyvCfa0zptx76g2U5r+T471Qrltue0IZ74e1e
paQv5vQh0i2uhhA3de3QXtpLXO2OKwSfWuPr6r7KZCRXudrKnWTByNWDSri5xdN4
DOrQqIeVkoyP+MG0b/LuT9PwG5HtOCi2KQvUROwUMp3ST5PCNm2+DVP2MAsi3btx
f3lM4Npqg3Er3YCxpQSbhx4LLTRJHT0p7jmrSbJwto/E/3DSc6YgD5AbpSTAZmdA
3/1qeB+4JvZgeqWbKzXtVZ9VTF9OFKJfynsaWRLtxD0W7zi3lu3oIkrXxQuBHUc4
ZQflNUg64CFLv5xF6bBY6P/9i4huRiEt/XR39r73uwhipF53zSWi8jgfDfwJCy/p
NspV/BgAquVEYKdYfRtSXyySJkeI4ilqpn/kHLpAC1nAHY5Y6M2ufJ0IX0Ni2Ulz
6l1JMPKFPiBRoqq4YoIncUCYF7lGF95ltNGae2oLpWf2Y/Xw0MFo9iXTr6FUMHf8
oeT20B1D1aA9P60kSsPHPvwCt7/VPN2qBe+4yx2vxeakC6BQes/aycl2RjIYIdzZ
y5fLYSrkguUDlhsjdQ4CyzC8Y9HEW5tzHQA2fCYh4wVakmKsgI+g2AsICqX8ANzu
ezR/UxdBI1jqT/5C7+womE8rPIBeV26sk4S9og/OB5TW345Lzp+fJME0JhVlQHtu
NseFSjNr7oJE6nf8iM8era0wO9XvtLgMdBLC1dgk9KfyJcaq5i0iWW+AaH+159ba
r2XEk1YO5qUynloRC/zw0/Sl9dU7LdoOCd0JQoG9gvgFSIx+Sk1KbyiHmV+TKj6x
9CbpaFefDTRjdqKckRbYp+sNfpcWS3ArgllJDjZ1b7UO9dqbjRBrfP1n2Kyg7nWG
77+wN+z0Mm55iSC2IX2Q263Lb46rvjj9+IyjqARVTCpGBy99LLWlXMy5LuLj7W1J
+iSFmEndfwUazoroQNubYiRtFjjNlM/WmIBNnH7gdmCVhFLeY3yIpgZNb70MVE7j
IKXsf0F4yZ0JTvekesKFg9GYaOAP466JCPWRFg6uAvp6570vmcq9uKybC/EhtsDq
62KTJCFzEcYr/0CuCM/9bf86YG2XTqDJj8miejNRd/LZsNYqTYRjkW2Jq3d6C9xz
XhkEoZFCcYsML/XIFbVoL2+DS04UH195Yu7iffrvIH/P2/hNbm17mB7ovn9beSR7
djVjbc1asbw99Kn7a5ybqwXkOugsKcg4sXHuMOjcyJZj8rYgvZ50N5whLPr2cD7A
QLpFLpODt2MRSOtgPOX0qdQZaeHgYxwMnIs/SoRCSrSE3T7Ef2Y2+32ymeyjiDbF
y4oSdu4V5CiJtLqwpPl+a65QO6JZD79lAmOij8BtHLs4RsnoKVM6X0abi9p3J/WY
ZzPpilsw/RxpcSwIP7/AbqTNVyzaqDE0LCmJcTZ41bf7KYmcpW6lgeG8DMxwHkF2
JnRsRYOZR4bGUI4um8fkGcorJworciRXjl8+NDAjQAfs383LCkLT7WLdGmrv29+A
Kckfmk0kAU9fXa+j6T0gPVJ4/931AgybTkcFKGY8mJLdPP1lSyV0gId9+K1eX+N9
Rlp2goUb0exZuWzpYxcRrC21FHfzwP/XXTZud9vP+Xg1KySAj2ralvKp94S+gR9Y
2rqpaN+PC5arSvGCRlk17PHeLa7LjgWuFqFmfAuPX2pLopfpd/17tfCxhGyQJevi
nWOEu8cMWr+3QXmENVI+ZEpvbWwX1laLvKEvKB+1wqw6z3Lmffqoxnu46UQ8QwS5
QNf7jPEVXu1BGFRql1v6EtmyoY1iSqvLwetZp0kC2c26fkO/6D66rK+sM1LUkW1E
fJP4ZbGJANkL9KEDZVjk/lU34sF/xC92lpnGqgKV66HejZXadvN6sRvbU3jv7op7
7GfMJzjntcViBGDQ3Q+HpYOERmQYGEzBouRCLyHt2YP9eyiiLzgg/csz0ZjWuZZk
/pnJbE0cTx9O+f63Plzn+rKaM8FI5yzR3AKJ3qqXfh38YzW9MaIFQeKIWCBkmyyR
lShq+OhLSQQ3tieS7qZjX91q88j/ask/0BeMItZ6GrpQyGYI3uX0piWOMLmg+Pga
Mqw3kSsJMuG3qmUmy1J3yRJLgeHtFh5IpzDy5KTCQ9sUGuQS16K21Rj+QxTAr/6l
2jpTSCj2JAFlbG+SR/oNhkmcjLPEB5eZe55H4hygaW9Bh9wKnsM1VvQacIuQG3zM
/1d7UUtjTrY3ui+TL1zSPqYQ5YxGJWGMzpN5k+63ZM9sRXDVYmx6fAEASczauP0p
i/tpd2p4fBkCO+91J7be6g9DSODcBYIjrcK/KyZIp3CUm/gnTj53b9tf6RkH82zw
Uq1ADeR4hLCSC/LnNg2kQrrcoEyG4v+89bRs2wWHy1VssI8HZbYciAjPiBiI+qhW
ciXltqZSM+/DeG9aEvXQOWvZoGy/TYeUC3JLjuX8/Iar+HukOxjLLdH5gxOHbgAi
RefwNvBqce+fHeq4+i6mWeSao/eLZVCu+T8gKBbZrh6LxV7OXTFE8CN+1Ncsmeyz
JTWkZYGR6aJNrEKQJfmDyGGWVcZPN3ng7WxBiG/gby+dxxaZ8LVHLjzIjEE7Annv
y1VFVap/SBPvlBw5TIi+SveF9eniaiCEk4HtQxB5d/bP/axGRb4B5G27KtPqWFPo
yRoVVYIhVpXI7H92teoNvJD9T8WBiluRjAZ3p0CDLBNZWG6as6Y56vYsbTRgb+o3
L7do3ao0tjfIB6pg4+C5o7An/o5qqw2wI94ary8FAJKz18Xy3eDMnwOT4iVerrqX
B3x9IQ1UjinBtOUH5Xa6EhMwrpixeRdDIPM2xRRPNCxtf8O0BzbRaL6VfQcOA5jn
TVyLgfvcmyCG4Rybl1BOnPoOM3MmWLBnDF9zhe0qmx8oRZ/WMlsWUL8APioJVwzU
P4DCBBtOcKsJ+bdg2A1sDwB4kG7ZCmpg674/zG/QULUJd05cDvqqa4RKtprUwjlG
/tnOcLUHDYrrX5GcKvpi04wfoNQUq3cEseSz1XAeT/d/QD72SldM2f9Ms9J+HoA5
A3yiMBJn/zxGnURqrqRCKG3eYRsXCBLR2LGrm3snyfJxsszIwOcvSXXX5e8hc+XI
Rx8r84ISh/lRD+ZFVfv+HCVoy2Hxasn1ZBz1GFYnbZN3cesoBwM96po3fN/IrBTv
+QgTyFTlD8eM+GbLkPrVfWoa+x7jD2RdbT7kTYJjSPNDpL/VDAyNAC+qWiDAu6kW
8rbneyOrAZv9wbHcp+SkUJUCa+KQHcZ7UIN1JfJDqxRhWA+V77UYOUJdYsfvNZol
P7hz1SncKnH/1umTmk84kal2KGnkGTV/6idCFKtC3vihollESo6DVZljjq4sqM1a
27OCuJ7LuUlj+pRsbzvVPgm7ut1tldJiR6hj0WRr0hSNHxZK9gJzf9dhRQWpEGd2
ByXC+OQEQoWVU3eoPzv2WbRps1Uuro/JVKvQ2+fVB7gZ0SCiNIfyLQTyEy9Tw9Cz
KWWWDXgWOpiiBAI6c+vexgSt5CYjo0RZyevoVtDoYpHkXUtstJIE/y01bmg1+Juf
DvjFtr7dt/2YOphejtNhTpAwm+CCgK/kOUaW2KZSYR785O2jVNjQQofY9DXEm4CF
HBnh5vkgoG+ggnPpPDYLfVfFntjyVnzAPlXVVORrbb2LG3VQgAts9HqO0rzdLkpx
m3BYLTvHvrT/vXkvYe1m9Cw5gWiHWX6jSJvtkWD6raAmyuMzq9G5WcBahB7QuHzB
vv8hGyYZU2VQkb6nsAECgJMOCrb4b2ACZw4ttrrK+IMmyP9jCZbcRt24I12MHRRI
uD8I3IJfELaWzG0WITzh92aoaPVH1hG++Sr+3RdIch5btxiiY0GPQDcC9wfPrHSB
4GnQMqPGvKPeqdcEQpUa4qVo7djg5eq1/EeAU1+R9QsRyTcLWpx69msoxXPSLZdj
BHwKSqmvQrg6Xr/aYl0iP1wkqig/tNP63cGixOCK5tsq4hHfstR4+7PVRLDGvdTG
ajTmnwJ90PqCqo0xqE5YSgbRl18xpbEmow3Er0wcv4VTJUkGLyk/WphlSQyTdcYM
CtlBoFJ3l/OJrDT5YkBGKVVb7JZWs6ZEzV8OVyY0ueLFaHkHmnlvO2owX7d6OL1Z
9OOg+QM/KwQGusTmkolVznqHUVApozEFqXN9GTMhE1gF/Q0j2pEbgdFxcMsTyLRk
BszCwMPF+mwTCyaptemLBQVHpY19hP5r2dUAWpApKA0PpuIoA6CcVqWkHjgt/65X
ZKREeS4+uNIM0cOxDoG7q3fBQVsxAbmyY+MoVgVja7iSCTdgF2KzsB3hLp8+K6zK
KoiNXkWSxDJg9VU1OKwewLVA8ud6wXgY1QMI5zK3XISJ/Xq6AqrVZCTHxZ7+/gfJ
TnDwWGBLNBPMLYpzBVbTIvp1RoTHBS5w7GinVSyL0skbsz7d7c6xum9oEvtmBPPu
HCCeP5z8SFZZqx3sn4fh9wnKysnr/qrYQWn1kdZhazPp1v9hFiW1qN/GQF6ZEuh8
mGor1+VmhxILj31SO1Ntfha3n/D8h4q0al+fG2wzV6PcCd9cpZ8Dz0uHabj1k1Gj
r824iS203+B9bjs9McfzLxlJIPwG83MLVjb318JqBfKo7fg053xPaRDzF21keS1q
hnPrH63XBWQFWUhCiZRsY2L0QL1wPIHKebE8SbRD3krHIhdJUftJCn9CsqIDRXL+
Shwx01eIo9n+jrSt9iCghwN/RYaCllc2iBmyjGociQ7J2+8hvj+4N+sxWV8ODkZ5
6N8mADF7xIFbJQDqIZB/t0gcGSLcMPi+b2009kp/QZN25wx+dPeCdjNfKO+RiQcP
4uRROBuPOkryppsigR5CZ+C4qj7+s4oIRViCHd5r4yPKMC1Ozzlbav74N2z8GeSO
sgvP8me9w+/LnjPyrWnhwN5KDJg6GsUNoEfwixfJlwK3jl+reyFLBndAuv3Jq8gl
Y/76p8dKQe01zPh/mo8I0zglVtXYTlqZBrI02h8bZ/gFy7r6G2tXmjaCA+xoy1gV
/Fmvm+SHNcYaoWhHTXoSJRmkUg5UAXi19Q5ou3eCTJRg9Qtb50aYJeXZ22rMaXrm
VI35JwZ8kZIGj3WX+Z5gy2g3FHaqc/JlzJqE3F23mN3B4eMjtLGFQ82mDG8AyIBP
bbBerT5+cAFlIMl/sgs9/z7Z8Q4+k2fmoa7VIPhUa25s7fiDDBdsiO1RFMlg5G0h
h6snOBDILt9ROr729KfBQgO6z6frMsxbcDJWMKaQ685NnImEvGSKbZBLzoNe0BnW
tShN5QvNq81qQ4kHJXRfQdMxORXttd6f4mtd/lw+S8zC2Wvh6JRLL5V5yhUDT87Q
ytWrMiofgAXMOEr07ZaoZs5WYEXEbBDOi9JNNKrO7c1oNvdk/iV/5mc7e7HVyCiS
9phb3PXDL6VhcAuk5cI/2ssN33+BiXEYYWvxyLHgCmGIMh7J69Jnker0eqOH547T
R/Q+07PhLve+1ahvro5k9Ht09LAevRWgr4KLvIbeOqHc202+oyWnelU8gCIjh3/Q
zlP5IOWgwbZELUIO+/Ed1bNDeXOsRypKMGs4n84XJl+4RfHMtBL/i0QL2LKEKq0f
Tyh5BwIEgvLqKk54JJiKHL9xGy3s6IVwktT23/HxlCsA2SSS1NJE7kfxAjyP1mU5
Ng6+4nc/MjQ5eDhKuldEdgpJmZQnmvsaE4ciyetyxdfl1rJeMMQNUm3AGCb/KfHh
iuF8dRDBymxRt63T32g4Q/wzImHnhk06tRsJtBtuSLGyCe2GGgksz1EyOXxrOl7b
AMckSDnbOK+bWjuE7OqnQ+l/OImhEA7sBZ9SgjQOTHLbXJzpQ1bovkh9bfJQT5/2
T/JEDP00XuwTjQaoz8g6JNc4ayFu3VeiE15nw5ap/GLbiy5Q5WXgzyy2PMv5Xfuz
EOnondzA6mEoLgbg703fKU6VETi7xcXoao1qD/uRjvzJ3+CItM7lYOAKLYmniOhQ
wJX/uCdRR/202lcQAa7TGGIw84wAgCtgBONXqm2GNtp2nfye4xiTkQ/zS8KK0OtR
0QnRQKesNSqOiDer/7XNoEjQtf59s4KPpDToCWig7i3cxukePq60mlpBTvrLr8ty
kkykIxx4LEWrxzgyBCjjVKGsYj4rqjdFseNNbX4HErxoJu6a3OmONBUFqNPr40sp
jdh1BLN+cUncXmoybs8aiU26LZSQ4NvGwn4q9/10UBh2LFs1H5jbbjDi6eK4MUTz
kN3HOxdJZKOTa+rJzYyj8ndfy5nv9ggob+DyJbJ822KZ9w0OIecCklH0q5WPcvFX
cKcZ2XJeFMjvRPLadCJfVkuhCltyzuIvI5cS9Pvl0E7fLbupOk6kuhyYsg/MxpIM
momVAD20AJjaRXxyh7JNOELeEjlRj5g7imfCfb3x3mmHzLMjXdXnJXjWUaPl71kv
HP+opRA9oYnOOE7iSXtm4Dz7rFY9afjoF1szMGlO6aW6P1wb4t5arXuX0kY+s/fp
ICDrSh62r0fwwM7PU8ffkG92ZJWkUnmcXIT/WoW3338DyjazZuVGKL810agoSru2
GX4EE2JNg1opY1Vb4pswkvnVwzRFg9i9MELvkaKfdIVfSfsJ/uTBB1K+/Yhxsm+r
A2IFp30d+dub3iG1iKyF94WU8Z0fiHgKczOFTKY/oa2RWdOjWmtKq5o4DB3Nl6+5
2BDyN9Q6kcfUDrI3TFeRU0Mttp8B/ndrOepk8iqsqscDPMw3F3rzwpGxz9smHA5R
MyPDhLV90OvtcaW+sLHZM7WuCJAMCWDXyfoFVMv/1DLyefSNlcCp5c5OKFNRDCqV
b/3lVAwZkZpIs6GG4TRyjlj0HrjWYiypdI+VIuNcPezwEqjdjG1TVsIdDitZux2u
8b9S//6NbBFjKdlAEca91kJNZjlpND3H5NqZivVmYhXJcevvf7w4Oy9dlLsDtMCr
Lkg8YyRFKxnsYFpdngOAXgWpSNYf6sJFzBFsRANjZTa3wRvypO6Qzxc7SOxh5zzc
MGfObPSdmYokDPtp7y2EN1G2cZuTRs2JxvenEF1aDVr2NOFXJqGij5jFmWip/54k
lWqhrTKKKcubOT/zzjvkADNl3vvQ5FZXZlCldZ15EO/cMCyb6rUAURlJkvvj0nCS
XFSnLxXfUoKk6nUt0OJBuj5aHTHk9RST3/XcBP7PAseq+OJogXnetA+ZrHLR5kVG
wsWNq8+jb/qo+2QTjyjkXuuBEVorae+yWP7OJOjg46Y1h2LHYJt8U0if4HZyXJO5
Ly1OS5OGghfUnrBrTDkVAG7QpCfb9ilgj/W/SPIp04Rsk2kQ5C2UaDHcwmDjVnDv
F2fmtGt3SV6qN+3xDHonKRufc6Egn/3waZ815IAaCHljDvNGXluZddk5AeylvLrE
ww4/722XTaIQP959+EczqbWZ6Ojf83Oe/W6b94Bx0MJUpa8EZk8o5/OvT7nNMzau
ChbCn/XJe80BWMALdnjgvWJjZyRoSEuAqmFNak20mluv+LKIwL4NxEE1RlCcWMRS
1qUhnNfvN5Gra74BzLV3aIOOrDxcBUT8et9N+epOIt2CVZkPyUGLntWvMXwH4/ts
JXzkbqCLtQyytmKqnr69qPLFt+m76o1TvhF0cWFo5PRNbnA+6zLT+gDIjXeHnuJF
V5ZtacRWbhXecv/RKqktE2poZ8+S7V1Yl89Bx2+7gnZD/bkAzxPas/GGW9FIkO22
LQ6KhjGYVLdy5FSEXmBWELNh+tjiGHF33zgjuUhNJOZPI8ZOnC6lsNthLHEVMLm/
+qBqtPpCntxzDKmTuhZE23AGMjTgFVF1ZsR9oawqFBv6H7nFg5bcv9cJDSrEXPCr
neOw2a2/2UliN8RRAxIBkU6pS39dq3jms4nl4b4wP4+vr5DAc9G58l1G6h0QDdHi
1CCMZ2feWwD5t2E+hLYYkMRYHpKAmfHR7n9E9StPHE4GufiIM6Y71J/kp09uwsOs
OmSUUepzu04VA1caADcE6naQ/WBrNCnk1Mq2ErZosDMxmT1FScig73/8x0f4x8tM
vAXEovKQMGj5OpuTbd48J+7cCg7282CP1Aw5XQIV6X3PG+ZzgVoachP8hzh+VEYt
abSH+2l513MbaP5QnaLqOHsZU4odyfr0Ma9jadLcj5PWnlt4UP8MW4+h+ISyL4sj
NbY4eFGu3/9inX2Mpf+VnSuL+e6iue3SWN14e/mjoimOnpmtE1han0UxX4rI4xgI
ugFjKGtZPXJcBSi5SNblegpwEa93SihIzuzwhx+mAE1Sf4OsGq8Ob5DyRUAmvPGs
pFQRQyPj2sgRa2JyAKepBtAKsTzTFqBryjuIkW81KTIceBPEeZE976Dpfz94fwfi
Fb0QoSYERNaQz/RHOO5XEAVjeTuiaibFl+n4yVCQVeMK3dZoGHumHc/BTyK4jmUG
FKokruf+/f/l4QIRRonJ4XGPI2LIKVHOnVt+pf0zxStuSaCNbLcB9yfCGoSsGyXs
1lGagwdty6ZqJMW8scvFI6bzc50Cf805P63Am3Ysie/urk5EJrBajCaUMD61qiWP
TonLIkPBgQWcpDoN979qrtajP6fU8iHsf1/MekWeuNSUlzayOCCWLf8TLhi1LCoF
I+rsxAXq/EUOV3kpuY2enOIsnjEAL5dpe6cQR5xQnf11njIhiKZa5TkKOq1go0Oc
m/GFeFfOnZWbhuchIDS5cj/uT8DJX2vQiBeCFeX2BCZgSTpyNQybFffIdX8iV4AU
me8n9xNLAJfh3whBkZYsMa4esuWoY0V6XGJhPqDH76U+GnVmmNXcCi0eWSy0bGXx
H1XPd1z/3uSFdkPgdLlZgp5BGAq2hbM3iJoAM8hbIIqouk67yqEPodRVonKKC2iR
cRxrPB8ViOy+xC5P8dLIjqRF+1k3qjQpr2jxDi+cy3f6NRyUT2uuxB64gQn7bXzE
F3qoa7lhzQ9h//Rahg83pstsMA8nuiVTIgtdzVazceg/Ae8hlTWEP8vKlfLjOXBE
LzEIyYrF1WzKKCL8KZ56ZUSWhX8Qd7M6zLfgHUwzxve0vSqAVvGKWxA/yed7VLRD
ogfnCXcj4Ft2jG/n6aFcv3WAQLQ7HfHRzUkAsqRcq6fm810Dp4d6b06jH0fJEmbZ
BWJmWQTQAnTeZJ1vHrG1ZOEakasMyHCGRLhT0px/9h4gtN1BJsgXUWl5AgQTHq2i
v7MnbNv65qNTXqOX5Z7benqe/f6JbWkbEG+wiIf3YzHtuSW3ddVc4ji+TZSfbYui
Gkjmj2WAcTXeW/xFR+yST66YjdZmiSof48srfY3o5g3I+YwecIcX2Ln0jR4TjYC/
+OxbDAP+cBgt4m5Cd8Xuz1I/TRwRKeehG2oSYkPzUlbt2vGtOGY05EMgssppSppE
I0SZ54QqWwyaDA3YgKnbrlMcyCDAqaYBhIXYQ47cNnLJAen0Ovx2aNnCx9UxVXXw
o2uULBkGf/qqI+ZUUdzkvBIzTvzsz30zhBR8t2G9YMORO4nofWx9EfDYiRaxRplh
EcF5gSeq28vjFgHamC29Ra+tY2ujXUgpBp30J8+Bde+UAfmQcGk/XSgzy/7EflT+
EndmE3UogH5DsC+RIVHFeZLcxZJjezh6SDHJNwQPbuvzGydcBBsj5qhcrtIN5n7d
6sViiOEKM4Bgar+/hmG7mcTAxv110oIxZlsKJ3RrTEqFVSswSouLHvx7CXIHvluC
6tLJeqyoMf1X60R8SmNewM53l8DAHXrey4P5B0Fnd4ipows9HCoekOicAhmTpjhM
3k+XG3kMu3foGWfrTvp4VRroSdWsUJic3kbDSZeHTcqv4RGFKC3hl83Nrn4W66c/
3Gfc6s+myIEkjkXzT27u51ZmSpwLCxgtriq9Y+w6b4aJqR6fgBMeKtn9Q0zd3YaL
TVecics46/c+08zkXoTJWvcsmCEgITNRpaujknNKXm1/LNFsqfw3+c1iw9G5jChm
GrNELSXXAUOC6o1/IkziDagXCPw3OfEwNvDjbSK0pyH3xNOgcQaM1N2uw+L3gEGA
V1x3s2/sRSTKbV9aYOcDaG+a2r5OGgma5C291AViHY/KGZ/+JLF+8XimRwNRYzgu
XvL+JOjBXIc1Wsk7cL0BWyA5AOhKbC8pBzl13ACUYxYtK8GHaffeG5IYtpDib8pH
kQigHcJcG7Y921DU/f7yV/M+yOOsmuUlWZKgTub9TGek4lXpb7Dsh+cJxOozMVSU
VqPz7L3zEGl0LqOZpMRNHeareCZHwVTGcOrSUXw8hdQZ9vEtPvqseoxoZMb/12WH
HK+tSawtJqqbsTRALcrgxrMEkufQ/C+TayTONvx7b8Ea/sgH7jJ0QUe+VVESwW5e
v38R4rtRi+nXjAuZsyv1vrBojBk9On962X5ZYRmjJ+qjbOoAJNYUSES2zyLQ9a12
XzzCLXrggdG6gEDXc+jXzgvEQ1W4KcWgCZXItFEvFxwv9dvSLoXTFo1OH+jT/sdm
Rs+VVsdIi1nRuZLoeUNn4RO5JxrQ5zC3X24qI+GrQtcYO0ssWqAFCzmHWdcwQMpi
HkDVntgy9jUKEHLzq+3lXHd2zFTyy+6HExFRlt298yvv7QRIIHO54S3HB2zV2uQx
a0Z4csGpzAOIzcM1JyaHATEEPPg0vrc+OIbc2Ls/ziSnxRoKFy8GHWNXUTAE2S8x
RC43s8NNuNJ9BZpoOIF1mzpwXzhNlz7y9ZbiRtfr3dcwCYa/bYIwQZq6NDMa8iWH
s6SYy9nfXkJp7iI9G4QPFCEGMXqc8DJXqlXsVd+xNV7abs8EGbXi+YV/wNtZYb4C
bneNf2EuvwHiMLoXvtS8qkrQOn825uANY8zcABRCGzC7V+5Juy/gdR8zNkA3PC9u
gccH20hUOi8jPPvSgbJ2kP6IcBpt6Ex7bqnvM+aEpkrgHLp2MVp9fc5wgnSl993e
afuBwEld0z9n4P2CQjVCCk/Nub4Yp94ufXvkDinOHiILpKJNlayRxlIY2HqLezyY
5DWk4r4QDOOVTJBpOobEEbabspzGwMFtBX55j3QHBif8O0LupgyeudxeH4UKPinf
gn9V4M50j9A1tLy77TQgCtXTLr2yFYCY1MoF31PPjlWuJyqtnZIV2GFl1Bfruq2h
Od/8uwgrw9AUU/uRr97KI7ndfrb8cHA5EFlnB9UEQA08Fddpav5/k6Nh4fUckssW
OE7ttKM1I95zdC5SeGHJmwb+Qd3Qz5sA5O0OXPIBoMxNVOLIhSwLwZAf6B7+ey7x
e2KxEj1qQc1TXMABT5qfqZMoRq6LN2OVb0zVEKSecpQG6ePkumLTlw8SQhVFW/Xj
rnFj8Xd+E942TZI5O5q83J0uZE42qAWQezkSv1CT6nUFoTeEknOTr6sjOEAAguj+
ZgpsrHVw8oH8JTnOglILv4hjfqQtTdbIMqq9ckNmQsPK97ZzRsFs18d4MMiyrjhe
TlfTQrkZR0a78GWASeh32OhqUdLzFIERSmgr81IYpizgTOgd9p1MekQ2fM4A0s9x
Ey3Zw5Hlovuw1nRxZpz/yi/M0uCo4PJ1aZu+P5u52nxA1R7NUEhy8/sy/EEGsPSd
JQvvM59WU06cdKbXaYfXpnLxWDKTkqBXadOq0wrPM0wxn9Mfsee+1DJ5C0HWjhfn
896HkWbbUv6rD2HJVrnFCRaPcAG94lLp0xJv2jwoauBwDSflemgOsjk5ad9GCw4v
G4QDB+KlCtwJIw92IEh1RYcMfNOJ1fLnDECdK0VjOyDF6TCwAFifPBCkEXc1aKkj
ong4itEDnj0iAz2HIvjHZXuLvguIWHmTNUWUcZI1oAlHa0oVF9MIOF75NHUKgjQh
ezadljky8Tlz4Pst9I8BlaTTVGQp6VQAdQk0r8RRBrv8RC0bkDZC78gDcTebFehj
UhnH6yCMM4I9gXI+fQp3z6YKDgTKWvEUWnZvBdzgO7etRWpkOZqn90hHg7guytYB
CjqWDHKNjlI5w3DUr7rm95qbHOYcnJGKG5uj/VJ06x0ElwBCGeXdbWXq8944z8YD
4i9UxKBCxDHRhREjktHlj5UyyBfKhpcTmTM94LlgfFCH58O9hkPiPtLIOZ14XMNq
ULwbvGXAtjOzDFKll4pwlvw6G8S0+ms5a6TNlfZh/iRHvWnVGXfYsEvvdibiWYVu
wU1w1ex/jnPhacn8GGWp7z4033SYRLjU4R2TgKAIBrkVZIighITPR6UZ3eh2w0eg
1ldcXEkaf/qerKMu8Qp/25FGjgQuWOiGOM8Q411gVG0h7qZxtEONmdPOIQ8JCyV0
KrMOtuRzzSJtGoQE25bpkxoSbSAUu9Cm04URI12xsA8eN2bTDfrbl6MHDoeAcXDj
mSLSzu8jiaa+VnU8eSI9P59Y46oY3AGPPHR6WnMvGk+g81BbtXYv0juMIlaKZQJC
doafj6UokYvJoVUQhAMggx1GLen8GWqGF6O1gKdFonPLP18hnsUJ6FJYdHzqqHH8
xiE53sM58K5MhKpjaUPJj/3xyXr7/oSO3raQdC33fG2LcqgXil4LE6zJDStKeHJP
KCd5TPmQxD8S9UJ2UVecR1lDN67c6m2hssqfKKJK2mKmUW+MQ67h02N1SVion8w0
EhV6gjmzBtIwjjbC1r31ycZbVTjlkxEa3isFGIBCnFHBxdrylGpoTaj+drhamedn
zjCilGQh6jvWS8SxuurBit5/vxeOGIfntMJxhCys/qIWVQEpNnPtRjXSR0xk6UGe
qda/FOM+USA7fd4N7V9Bq3mopkDMnvpIE+puQ2eqsRRNgfs/qmjMVuJ9GLiHKjBs
8DszJ5eFeYN4CsQpS1wXa26MqfuKLankNo1MHBSwLmxK6kBo1AYivXYa43nFpKRE
P/FpIuAv5s6IMjov5Klm2yvY3puVufYW1d+tqhM6o6asKMzShhQ/fqPzJFdyi53b
tV/3zqT/IfzHVeH1V+RQHk4rU29CcAYoJ75tVgQYvD9g6xX3Ep0/HNe8nAusnagH
dx2HnZwsKGUR1ChSeO+zdLQu/fBfj+dCt2J4pgHvH+gI1zxgEDu0UVqOxEVBLpsM
L68EfAZby9OPTyOyxWfMrfzC1aDWWo88c+qd8SIaulgxGmvjKn8Xc4PCFnypVlt0
mSeWM6phhahr8b1bjhgRNEOYdSx/F8RlK0Ajxn+0zZlT7L5/pliFXLFg+elFiweA
btjiASZ5+sB9Z/kf7cwrxET+0/jAPBgLmjO9mt+PZvBuZCyb+28AzMu+hBSkhHqV
PBYFJrO6lYaVU8BXXOI+zHUjDKPpfNxmXM/SkF3X/H21zceNHtdzbwZ7MHU3okIg
/SM3of4KDNY6noeJU+ezeuNqj7eun9JwiClhqCgYmC2/j6EmzQkpXqtgqQPUYXMa
mSDINs3zwSwmG9Vmeo3p4hkvED4ve8nJ4sUfD2UrbKwdWG+eqJXJWkjD8svpRK3q
0Wb0cgYqrjx9Xcc3smoWinxBf7WO+anOvQb8MI5AwSohJc18k0cXUjbESBx8NEl1
xexWCSsn3EIMoPz6FqmHIr9IOD9jDoCXeo47P21RdX6EaZK7fW3b2l+noN/sTquR
KQQLnX3DljiaQZvRARaHBooGAaVNMKQHtCH2kHUJPzwNJNZ2b+Inld/5Zf7VNcUM
kIkDW+YMldwS/ghWZYIh+GVx8QWajNhwXBvY1FTSNi29haYzMcH+Itj7mYSEr/y/
u9nMnieD5ISoiLI1gYeUO6SvMZfXpxWd6Rvxh5/X8dNzV2t1RESSb+h60pw9KvJT
P1ez2ZdaL1/R1GW9qTZLbEuS2mKv7cyE0xKAu+RIUVOyWIU0YZLs1HWAJrQ9xT4i
cW6HSz+AKHPQrRdJiTsfeLUjIm+u7DLdFCchbPN2wM8y5k8S2UnEQrtn5M4itiMc
iX47uQbJcPwBsORgM0/+jODAuBe+JXEI0GTB96OSERiBsqpjh/vLm/WPjq9Jomdk
eeSgR27a7U0wpfT9mY6AK7QbBCpekM2VZQ8QBsqee+CT8zHc91a203JupSwkIQVL
hfpi7np/5rPyJcny9Wq8sr6/cxurdrB+QuUeWFGse8aBEoMWMA6AfV2RcBsnfpB5
UaMGr2VjOcIXNQ4L7/b/4NZ+mpQuv9gER4oOikQ2bf0jeEQY7kLZAlP/OG0kmqPC
nbpVvJA2evwKecvVUau1hN04iqrTPJlmrhn6lgu+5rWmO9upcjIQ97JPy2HxnNW0
RoTq+mhh5aQiUTPn1xWMfi5ghs27Z2r3/1GDkL10CnbRnvONCMRopxwtvqg6k551
zACIFW0P/AvU8BmIaHIHCElR/8xbWXtuQOVQTQEnSCu7eEX6OwcGAtweCb1Frhzt
5DQ9deX29pom7qkevkNLW7sjoP4NTWorcKCVRzey8nE9FgtIBqoK2306Q+NT8CRI
X4tUFKiExpiew6TSeDNJBRTOWOHHYCZXtBSppdw9FcUpzzTI7SK+cicSuF0XrIXK
VduGOGIrETpj0w1L8NRl9gjFyzKh3oTU3rc736Rdjb+vc9hpM9lrJIzMMXxLLrzk
ObfDuE6/BE89fJeZ3BqZRtfZS1If0ngIzKfZ9SbxKVC9j25fro1Gx9yUQca9R5Ez
UeqcoDbZgh+gaivr5sNI9A/bxTHjSaoVeVUOrfH8rK1yLa5mCTV8PMVnrEaEQWjE
h8KnyQdqCDco0RBqBoOnwjMVizNpXDRkpLYFR8b6vqblvALOEs84aUZjsICpSTQZ
Je15C2LsS9Db52Cazs+Aky1n25M4fSQ0glnEojSfnWgF+fIxA+wZgl26nbhRNy4y
LRhcS7EY4iCKMrB83gRH7GcgskAVZFa49ql+U1o7fSA01E7nUN5few6mDV0kFU77
gGDnfWP/DA8iB8FucpFT9gghhMnPuV3A3geXt4MNc6KRS6lfDMGK16htJqTXlUew
AQydZ/Wp9eE1cEQCW3GcIYyaZ61HDHHvQ+MMqhvPkQymlk3vloRyZN1+cNEAgKHR
CI3B6HS1G69vgArNtpsQltBodiyWJRpXMhNt3iY3nlBm1uBlLLZMMnP8/6HuZU78
0qNsl3P+s+Q2Y/rkbc2+bf1lX9l+l6v4265UNBi7TZDqR2DdyHc28tZHKHMXisRS
Ur7FSqjPO2mrGcbq8TZUTZ2zji2n5H65ZaNSN7UhvxkUciggDGDtjqIFWxSn5Mq9
wuQh7D28RZUYYkERwgYq+ufri2pSLn8wrjKx/m1UmoRcrMefbLltcyMEVc8IVi7N
XCTtdNcN7hchaKwyNGT5WLheLHTwWn3akn7WbxOwgY9QUIUtQaPUbk9aE02OQC+E
uCoukU2lYoPnmOWdl8g6ay+so4oQWDdoc/NSpL21WHHOQwEHS01PVTr6oC7oE8UK
DOcAg3yutaReu5Xk2oXskv1cYjT0T/sIcYJpgiH6PSTykGhVZ0YvuKMIcJAI7t4t
XSRA4F/pmgvaltvplvM3xa6+eQg2lN1qspFC2Juq6bV1ddyI/dBWLBr7fF0yv8TD
Gm9vq2M6mhQVgrneVIIDFNzB92CHAq8Zrz9WJQfHf09OVg1M/CzfGKtf45dLW7pI
FFh8/c/nlDH/QOBm5F/p4lUMEmucN5zHJfoBIX/aT1ytLyeP5kKtZfCAdBcll7lM
MF4J9WBEMswojoyWIy9W1FIpxgb61zIMstr9GBfzvQU20N4sFTUvUgMgWBASaXk1
K0F7rvYlslSO/pSuo0LewXWiUtKIOYm8PGu748wedM7kgvvKA6N5dux/RF+GNtI/
5B5DFiIemvlzzn0Cm2j1AyDG1vj8RkAXkDGo2boIW/iUSNMI8Zkzy7HSh7AJ+BsE
rU9A0szD1WSt67LHBxZs5eKfCLHWHNDEgk8xxNmxra5ZRUCeNTqe8mYOtZiZ8ryq
6RjB8IIGgSO3uInCOSHP/CVqvkt4RzTH+3Gc0h6H0F+w5iUSOsv0beHfbx8VQFLM
kL9zY9xiqWtHCGpLKhkBws8bsvWDm0GhykN4s93StvnUiM1SWQemaWSh96e4cl9v
xgR8fU/SZRzl4sMQx1ksNMJf+WZWPquED8W7ffIlUORk9dLynXFlSywH7w3WURnH
Pfx4BcQqHu4LnkfscyZH0JmY+gpMCSZ0guHTehFGbJrX4LgstEje4wCKwQi1q3VK
AU416UmKiRyEjLzL0Arx0a8Zyb0Wu8LGkYuzzOrlc5xvBZ9+7klViG2AVB5ksIiv
znsIAdsEBENU+pgXT6B3Ykn8s+YTVWmzR2ClL75QBzjNB9WLshLlmb2QluzA5vSH
El6ynwQciY1etFqaOC1YyvxMLNB1jk3QdWQGnbo+oH7MBtIAKu1qFUzQ2mZYP684
h7ChbN+pdR8Lpb/OjILSBUQjiGMKd+mw4e+fqH0JCa6aHYz21AkehEkqY0foI/wp
EZ+7D6ppR3gFBqSOyvrh6Ws2mAexNkPnKm093JQkZR/0kl4wh36gQkcjKj8UJwEH
JsjZk5vpkJ1jnlivFV3DCRi5g8AADkMDwOIF8k/Pmo19VQNLsMeL/getZFultHmE
6VPDTOlbeQnT6pViJk2/zXFeKISkTnvHLz6qn+O1t+8F/pfU0H8W81Dci23yMYEy
XPe4sQuFregIFkkirsTrnBL8L0a8V8OJsOzKpT/j8DcpdSjrgFB+gvtxYjll7ara
+tNk2pSi4+++eQ3646sh1loFLFVQeVX/EUkFyvcELfKr9IWTEw8SmvtY6FhROQSK
r80y8M82NwkAUqw52HBOX/ax45lbwSP3Jjo+J2h7ZTIea5mX2owMfnHBLNsrONZL
loulM7hqc5ftjKRaTbte1wHm2LPLDVyxsD5spohG26xHOXA/r8+9t1TdIMoIM+nO
Jtrp/Nm4YyE8jfN8ZyaoKCJrv0qAxX6DJdaI1tTClnFrj/PB8/aAcLsvUY+q8sms
kTv3VRpMt59TZovXBwA8yy/dZ+amsTtx48S1UjJ9pFC3ciZhhpax6PVg/ShjmJH6
D+36Fuz2IQn4iNo7gu3LcB6m9oD1kTd/10dwYWVGY8AVlHeCkS3dmP6HIlPPuXuL
uO3sw2mTGD9R31/7HKpeqg3vkKYGH5Um0TDE0gsr90QiQuB9l/HXCk+l7EM0LRi/
J8XozBpX6rRt9mehyQz7QHtJRzP5YE9wOWNOJYh96savc4/VXjOKKaANs2c17DBW
i1XKyQnm+JR91WH0bUY9+sDmt4fNwIg+X1cqHBbrPCs4cg5Q/I+sPqhYdptOyX9U
O9to451oOX6hYmnrotElmsP6+1oq7p2S9B5TMhzEnYJdBusGowVfEHJCvDJhFa9D
b3kdKuSMKPfgS143WqpNMfRmQwJ1UXAQ5v+jh57M7taFuVZGrLiSveK9/IRnDcTa
QFB8obs+2bIq7gG4EQoJB8kiEM5a8BZvqdCNgjay/FeyuO87r34ac6X4Td8XRo2U
cYKJ8Q8Qc2LULB7eK+rT4UkjjXlnSMohfeMB81B4WYx4fpMg2Js+VJsCrn1EIggE
RSFNr9UAOGSoc1h/96EUo/qGC2VMUnYDf5QeS59GKiQepEmd5XHUBTm/6+A7O51y
XU6H70guE2bidjH2xypfObSjdpuVdigDjgHAFobfqrJKEKPowsx8SHBH/Bge/qBI
ODCXDS/5pH9Eo+BQShacy2X/cZjvVEp9zNIFtCYLR0QBdyMHLFfXiMHrc9sZER26
cLMaq99BM76vc+f21dQDH71ZH0WZXTMJJqwAwEauAW1I8l4yfGdtY09ktHjn09Lb
2qTgUIJ+CWiKp7sfsYG19NluAfnjY6k6ZmwWhZ4DxlhZ1bNjheq08yUxmAma2JFM
eCdxZDj0c9yto3ooskUmjtiyJy6Uz/KUg8eN/+eOlsjkoWz/JNL0VXCZi0Fy1NWq
gREUHGW4ILr5Fbv3mckBo4AHSlE+Iw11nPYmJ39exf9nkSiAv1BZQGHZFV+EYMmW
++aW/fhPDiOsKY/sTYhlabWq1J1E427c1xbO0bFwZe7OmbAADtL/I5005cB/LHww
x3Sqekw2Nj6JEf6ZlPSn0pvUYWJUhWZNkdJu4Z8dT2RgI99y6tesrT/UZ90OnnxZ
TKFTWNU1yuxdi12Gtp6l80TLOIXZ3QwcioNWxah3X5qMjAy1WXfSqDTP5shqms3Y
Zhj4km72c6HI73XDBgNNnn5lok85RUicang2jv+WP8TpxHYDMt5ehSJ4fVnK84bZ
PHDKpVlrAUYx/JMTeC+LMBSXfvhuSOUclcUawO/Y1W2e8dJOC1geX6uqIqMYoCFm
QdDzn+vmG0OxsW33Tgkffy6cEk22nB6imDyhqjZuEn/vF9NjlPH73UgxQMdGmns/
zHSMECz8pzi++CWUYAPUsyj/hvnA1E1siVLjQSaZD6KwAvlO17LzzLbb2cpTryGR
uTyw67RfyJLnsZh7gI44BSJcP7YLTO+J+3B/qFq41TskViRgfp+LrVpFne938dRx
z63QIZVQHW7ChsP9W/DhBSJhj643TEMpPnpXqapn7/jaGZqQD7kXjRafKBxUcRE8
Axl23I2YKD8dH9eS1lZpeDYfPF2nN0+nXeH+DGxHscGh2DLyhOYkHS0RUCRrMmKL
jw6wxbitpRXQc13myoXKVureLAHNPx3XDS7yK1yM23E0plNQNZztCHeVfDjFHQJP
06XbqJt5+NgqmMNAcjmgJ7df3Fcyc4BKVIJpqTLrflnc9IqtEZNa3b4psqdUcORG
NCWVh7ImFqcwBdsCHaEfkrufynJWmQjQBVU7KcLyZS4qd1OPk48gaswo34gqy1ZV
oNA8/Fq2bhpQ4JNNCjmzDVl4vJAxZPL8S10EKLFJG4CY0RhJcdwEQirZIDKdX7jg
UYdbODjmX1HcUAxCgnzRNPCd14LjQVn/BpIpbgGYAf81KZlh+0SAUAKe4OxbkGjw
zR+ftXZ5z3vxDR9gdxCjWX4GyZpmxgYIhj0btu53o3wizZYs6LXUAPWDeO4xFuk1
kggQoeOmzPG26knGfdk+GDExlZa6Ljh9A/7bDUjOG0ofDt0gBhpTDDt01ETI65sx
5a8H3Ec2Go0AAGX7F/BY7OwOATs/Z4bXsoRplDFit1KzPOAoqnuq5ehraX1/SKvO
uRO4tPNtiUBsMGTgxh8cUBTiQBS2aKdlxSswYPSbKn1gK+1ZA/p9kG4wyi8vESDa
c6JFDXK49zHo/o6U6lt5vWgEng+HM/+pWG+PFvJK1m1v9EnpuEoeQo8Z+T2+zNek
Rw2BGBxB1nssy3IpsQi5HRXjab9TbPf/REXRvTPVwGzFWJNuEbZBi9aw6Ln0W55N
4l3w3e1uWYNeLIMuPC1bot/pI872tibOcdK4KaFHWS9DbzF1mKX0Xtg0cU9JZJGD
GKw1doRFnhHLWMcWNos3op0zQbxXdw33vvTc2rSWDdclRYJsCOmUBxjIgZ47JFIe
SSHO/i8qNe6YPzWvfFUIPH2cdPo52M3JtxfiCSFw1Q1co1yiJtZ9ps4ebWNxYI2S
BnH95A6sbfIAKGQDzhgwT/dh80MbMGmZuAnv3G6Z0NUsQCPczsfXljswkDsmHcsM
CvmK9qxa9BAATxCmee5byi3NEBgdN9tSC2ug9U0q6OvA7I+KM6P+SO48utEKyJ55
kp1dKiUmGfIYeMyuierVCF6xD4+ybHiKBQpsYVj+RUFhNI8fihwWZn1Qccwzo1D9
Y29+31LaBjWYAqzIg5Eg11RyjukXGA3sHWiZKXKnF+wSAJV7YnSIlplpE9WE9aY7
JGeiqm3ElDa7h4E3h/AkFbBQDR/v0kJ1HyqejlKINhdWZCL+l9z/1t8kLpyFrJ9i
1AjprazqQiKnXRD0+tAwNanOC/fxbyg7oqQHlPcfB1CFE3FUlhjhe1pYSOF6QBkU
pL2wfsQIksXE39QVHVqxJ4H5klPS68PmWja4Q13rn/wQrAtg6ouSu7Eno2Pp5sKG
Mem7E/JIzN0sTp7AHdV3yZAgvQJ/ufkhAcavQbK0EHxNvGMAPUGvuss26eS8v9+c
D0GcOl13+rWmx/N0Hy/TfmoFWudom0auN7SbdeJH/A7jgGHhLalELXpx80RPoXgD
3zrXh96yIteJMiz7CzqCD6hjHEhrGZSfsawRxT/SiZXnnNIcSH/cgeZkUdOjX839
ALlWg0xuUkVVTPAmvvZnkPaObK/WAnsTTx4etU8dgfleDmpcSIKpmvKAUv4VxVEt
tkbNZp/iJcNs3cI19Zsn2J/b5C6+pfcEuRMc3JqhOatdhcSi927kMRk6U66H5BNj
8p5hW5CuQPlhTs+XBnJG5NGtQ4wqRTz8sKYAoC8mhs723jLrc0VRL4RE8nlgeGzi
FsN9fmyXUFKn34PeoJ/aqmDMgSOj+nFGTJnAD0DJkZUXUVIiaEpcJ+1iK7p6BnI4
g66cK1Y3dgkRV6v+xVaqhla6luOC0eZxwpCoxOO38Yhb0XxNftBHPTO3GpaEFd6f
vIdtKFJsZInfLhpaSo4GWWMj4rVhxjkMYg6boXDKaldGQ3Aaz02/HzMbxtBTh/ei
CVMmlsugDtNr1x91U6YA1jaMEjUbbcC5cBliWIwzGUcJxesDgl/5IkhtPoH4QD7U
HHYsDk/U55MebIs9b943JtWnlVU4FcRNpYyB6tNgLpNJ1huEx7H6m4NB2EX0RuHR
WDOtIiJntWGfOJS7a5BU+qUmC1rIFyDjC4bUPUQ4+maM7N0nEZ87C0JjDb01UCP5
EQRn7pLE7CdjBpTTQKlTHj6Jdf9iyrqH55hpaQZAsgmEYekNtNeFGfBUs55Kmwr8
i9EVZBWNluUQJGYDe32jB8+PsSCElGSVYAO2tzZDOEQXreipHeEVvYvGW7hf2L6c
sfzQ98V2Qsm0XWL4vUfAygngvr9saJx6W9qjR0ExFgmP50KlkdvL8THmuMWMbFmR
i1OFA5GG4bUwrzsU85g7X/F2pI4m3PCze1JHlLmX8oKynTwvOOmSzyCCkeKrYJZL
aYVEnMdSqrn1dOYZbNWRHfDD2VPrqk6NTRNH6+War41dOs38QUI6OJBTs2EQtbvL
WJqq86RCpEWminIjICeXiqUvpqyXZxWqIc+CGsLS2s+5Xk8ecUydMTjVmoNTNV82
OqK0fJPG/SoGyfrdmsqcUiMydbSYox4K1zmY/ifyLKOxVJXI0CwYub7a6S+SsEXz
nT6IAHpj79CWUCQsY5cCs9x9e3Un7iDoEnz+gPR9mWT8ilx5luxX4lZzAtywOE2Y
CmBA1CIRU/8zfxUnp37Wm2n0VmpGm56E86RXFlcTx5ido9acok99lKVQzqzEqwUr
E4b99qp5ENbKaU/HJCXGx9A7BF2nzX53I2U9lNrFMTZG+ZcjvKWb6BxoQVh/y/SU
212t6FF2bITrLPwJAMrZUKa1Ck46gaZgyjA56vdke9gC++Ge2BEVBO3fJ3sw2YNl
zmzKI+UbRlgpfHe4BxZKK4YHY2iM+GAqI5G/+wPvWRJ/E95JHzeLyRwPWW4R1qXw
C8iba5eooA9Su+tahe6X7rLUe/UTDXu2pSsvHWdgAGFrDPoigUxOMuO7nX/DvOSG
a8JbDGyJbdPsoFbR/vkcaFp1PQaL7WCiDjYzAs8IUJXEpnvxBS78Fhs69LR0j9ar
aj5ek3N5ugU6vfRIaQ46Tb9fZaGkUT0emjFXYMix0PAiNErTzDOtwDt9jpuk3UOT
I54Ipbrrpxi1PyRWu/bBeHca5rLD3/xZh8SjA8MZGNUzQIue/P/W/8YaLvoEXOh4
G9i0djpo+v0Oj3ZpDAH4QhHT/CSWI8jHTq0YJhJf1wbKlPy/DX1886NDQfIEGFAI
zwSJqK+3ts9xo5BwrTdfJwbUdhxnIGl6kOBf7SPGoIZds6LKFunkOE7c+2rPab71
MgkhMYWym/USxQCJujWEe+C5TWSf8xHMQ5aGj3xn8fzIU2bykacDCwHrqGzhumAX
0qQJ4wS4MG3kxVFYeBPt6CWpsY080q9kYQmphieOunO25zjAn1Y6v85TaOnpmbmA
eQwrjEy/T/03BoE21q3JxKJzOdCU98AzRrrHWHQgxQnkyZbKNUwjCK381etVpg9q
J5XVkEZoQfcqDkmBZnGQ893jdUqNmMy9GQApLfOjzI0kgjyDT4tr2PC//mupMtRZ
zz07Ue6QZ9Wdi/q8a1ciZVotlgPdZ9s4xGuLVE9zJcbEdIBLtZ0TvqW8F8ckoctY
eVhKHlfjqdUbwI5B6lkXdzkk5xRPmQm+3wQvFeMseU/2v98sdxYfuS/UC4O0UMpz
vDKjOfC4bVJSnBmraSrees/oPKDc1xTusDW7vBfloFiGUejPrvSYXT4uXBAY3l0x
+0gikgXU1H2b8+MHQPiHrjDYAMwDxqbAHfInsOoSHoh9Ej9wnudOxt4HGdf2r0WC
LIsTqxf1WdYnFZRopBNW4qdle1fq5e/qIsGdXW0dD2/o97s0BPWkALG8p09LNUDX
9hLtPFoEw7tcaKe2Txqq9Go+4CqIU+8vwOCU+aw3zSTzk2y/BxqKbPn88GtgQWK5
8adV1S2GGftxdrJK0oCOppqtVh2ibTcnvq5vw1fFlbN+EJ2BWTn+hr4iQaeoZpkN
+JvNt7dW9jj8ozpZj/BabSNgVk0NRe4CU4aLPKsqPKm8ONwnIEjwYhyXlrDUBlv+
5Ajv9HohWd59pbxBnk3yzBygd6dgxPP6E8132KjjdTuSw75Hkf1uO2G8nGAvD95B
PHbuIW1LLMAfeS6w+nxI7gk+ugZ9ncARuQdCk/DDS0rlXuFNEfCB6AoPpXhduwBI
mA9Ly36zFV6xqi3IFXZgncmJTJOmVJ/7/dBxChN6WEmFA2bMFH7lXQyggkh6lGZu
HzJ8jN4MatG7XbrpQjzoh6NMa53skcx/svL3sDXKnc/imWkvl6bDyFBdY1iimi/s
MDylURe2XNlg746MNszkbPttdsmXLaQi8quWk6nK81IYuGlK8TldxJxcmZVwtlOz
2pKykW6+qKizAxu714D0rtntXyEgCrtcH9s+f3zkVqwzV8+LJfk9TVPvkg2F/pNk
UsPmTGnPJMKdBcReXWZvBb8S8gkjd/zmtf4FD1ezVmSyNq4cqoJjxaYa1598ARq2
/9rfg2JUgv3Nw0PBoCNwoQADdSkchZ+vbdyjSPy2STajaxC8uVW4VK1wVYqnGtoU
rAd0xKwuPHPwlchvMTNSfZTB7EUaQf3KRPOYTmIsdIXH9/j/BKs+8Xpsmzavk/pp
DClhO6K4x9oQo1ejz/yiCzNXH6V1sSArheGTfPlCv6XQ1pGXGLCe+H5vnol6W4UD
kreqJgTnaBRrRIY4l+Yx/FubXuTYYYuCW63VxAbjcaMMgHcLxquzzpSOKvyIRGap
zCtnfPdI40xrn6+3llj6zKFcitE8lLQm7yM7+1GRZIsUY7OHcqdexlC77OUrG23L
06ZPXxeTzKX3OdPhVXZayca+oQKe1YwpM+bX/SwInV2TocuYlo7AGbcghtHh2cLY
ZFCgrQ+NtXpngXJs+IUwFmTHWcoopsqB0VD9cXY8oO5iW/ijZ3R8y4vpt34ovf0z
CWkKHnWpZCzw+y8z7PfkCCoUVeFKKPS49plfmu9lY6v0SrTI2DWBnON12iRlqhNm
qczSXLPiftNXuV3rJnbcE0mryMhrd9GJsXHAowt+VkdhkJ5G1x5OrgQj420vOAmj
EKQbdBD0h8HqrChRixCwja+tQdAVPV/A4e4jOb9SCiR0Kq8Jx49F1YJMIGwibJsw
DMq8d4puq+VQvL05iqL4JUJ7+aobm5/DnxuVxcDI1umwQhFUHqNPPXMlXTULfQki
fz9OW68p3sh0MDe4TMd5aIWhVfW331GJ6XI7RswAFZnex4wJH0OM6V0dyHuhCSXL
nztHo00hXIuKOoabfWTworzqBLVZNngSynh5TExIk6gzlZpCliODr1Y9Ve+NVxB4
zxaIae90GgChCNTy8RD8Ip2ji14XdGNbPSY5zwK+u39kuNDOlQrMCf+LyW4/86SY
pqNjZXCtAMq4HFGfC0TxwNm18KGvKSrCV6rbUqWENAhGb0I3iAjinCyLs7e3lzuO
7qCXPIL212iuxfHGRaEpgNIwmKvnh7+6L+5SVcIosm4jhT1vOeaad0IOOFIu68Zv
Y7nABapQINn8dlJtqO24zUr9fFqaDZhBbnuMq4MMIz9q2MzKJY0FWVWJeVSMB9zK
ijNSl4KMekLv8y12w7XFyta+0G3WnWUpTRozWq3/KJJ6xQCSrMDKHsTBHtMFS7y8
3dVi6UN2akTe2UEKplrUI9kPUzafzvg+OCbgBBqqR6IlDfZl0iazVEs1mc5NYsH0
jr3RFxE15mtQW6PHOk0zILlwEjitrp7AtZwVZSKv6SBrZsYPIO1drirZ0rh3gdFE
uRLCYBysr8EmF+RbxFBFu0YIMt/injKBm3rSMp4/wWeFZP38DVJPvonq2O27Vflo
qses1oiIplH8uq9BLmSGXgjDLnHlsZEpTH7lS2l6DRt956Eb3WlTPuuyUe3pHImB
bnV4O9S92bl0vwT27U3InXv8T7ShUGMfZuovDnSWEo703jYy04fUjB8XBbXmKpLH
jIwJSZk6d/WF/kOkvKsBz4ooe+wcKQhXi6wHkv6OOw8WE3VJTOQDL0ChBKH8e5S8
jhvn083xkiVE0R95YbHv6L1NNcvgcvUqmz2DDUdqzuu+O6YYtvRsW1OGkIOQJde8
2hn9ldWF+TIywWs3w4sKdUNccw4lRj4cBqpIU9DW4FWHQjBwEKdQJwTXxsLogp1K
9C1o6hC0Pxb3Qa3PRzSKVXMJ0wu5b4peZ7W3COJYaA7qw0qzMDOM12RUpJD4dvMH
+nZ2EBrEn4a8ao1Mgynp/TAuQRDTSAnYzB742c3/lZul1TQJvwC44XAy3maBRMFJ
LrpVO8LwPshq9vuCvvOszqy2lX0lO2GGAHSJAit6HxZ9f9OfsnO2SRHM8ytG7rBM
1ZkOkQFxqEMpS4XCKa90ElSyZqisvCLcPG0GCxaMUbvkgpXiQNHZW7uIxGbOfP5l
ta+bFuNqriVFevLIiiVEvVFYcA8oLte1Crut/GZtwXOwmCz8kIP0mmFebfR9UioT
JkclPQ9BqlUn5db9AZgNsjIuDyPVo5e7eQsdlGltL8dVEYcfp7Z4tUSumVwnPG3S
F8fmurivSECgrg3ZhDIwwKz3HcQDeBD4DY6zgMSCMAveYmuNOrgObpna2MfKVClH
vZNTnwa07oC8enHqhGRHFtqZmmt2qbCXPFd4mJ4pMnNNO+qRDrmei7MNpkde/hQY
I633AiKARLrJleFMQxANr5+OBicVh6G4bLyAIlgfAwuQsnq8oVpTvsdvVkihcsz9
VFFA79a1ZHLDh6QNzLRwq+IFUWBjdluDWGQ7uz8NsSD530SP3qC6C04ZrrclTQwl
6ItiIeQIaT1VIxX8eBtIg3GcGh9NlibRIKxNzeTLMxq/EtSCYoly3u5Kqrh2MbMc
dhNZGomPEd1u5QryEQwiE9Wm38/O6Hm8p+j7YH3jQ0KsM2v7c39xs1iQ0aL9iRoM
OnQ0U4mL2EE7M5PNxxUp8C6hEiLsE07NneC00tXhi+RzEprJfa31/UWWZKM/hrAJ
LxPCsJMS4dAo/QzMaGhRkKPyEKDMmq9AxA/M9R8j5c6Ng4W5p/2CNfalZ2Ipok/+
lsYY0LUOxRAHRyhITAUymEeFRiL985cuHuvfY4ejtkN6F6VyGTmGLNumEs1okqf9
BGlRIH9x/a9TOFPerg2dM1DURjGVR+jUmUsEgWM3YibwaBFJ/lVo2QMtFuJjw/Ao
0NHicUpAp5Q4lQhuKkI7nZBHJpWAbKjagbPppgJr8HEG2hhqRc+0YnGX5DqjNAVU
21ktYje6zK1VrvmdgfzRa+qRq+vGVj5U3bjwfuL/kbQ+GKtg1zQ2shZAsLjtADG5
ZJAK9OUyErN1uOVxXhjx1TqJnIWs5kFNEWvxNM9i4flcbkH80Hiz/p35MZweGYlm
o7k9L6negqaW+/sT2wezEKtBNMC1t6o+GAVJKO64XH37ujI+fyA5rlfgoOdkh6JK
U9qdwOQKfImqQEPHS0deZiFD5dNTXQyj7GFXKR/RhwgaqLn7QnS4z3yzBGYt1yHV
tSKqPURFb3+mMYBOQU5dBL2AsN3HnfWKCREXLOSZZF05lFnIsbiErdTHC7gZQx3V
z9hy8mu9pLN92UwPRz+HJP0mCkopRFm9/VWBKpGDqhkrpZfYd1ofwV6zsuTq4sTv
4WxlWFSsaxRkytfOOh5LN+OoTsa3pyKYoWZ5TUk3XSRSd49bXoUVqjoGYjZIXIWy
Ns7NhgWE5XugVtyH7aXjgu+uwA/QAtpw74HX6No7wnhRGPRlSRDMh1CaKPiebcEx
TXejihtQzYs7ctm3B8ziArgKSsozGpKbHHJeDN2ZHFWn+EwYvEAcxY8JZ9C1SAlX
CCneqpwKm89ErnayB1+RRDrgrd/0tsbO2ppLMt1DWkH3QPkaU9zuvKDE2qAGRwjj
hb48kBbfpFnkcfpZPb8/aDh8yLNfs0n/e4n+d81IGrsRN2Xg3+76zZhOdwwbe2ck
rOObWadRLUPcIO3/SslbF6ksGSsiIXeN5SA7LTyINindbk3u1g7zJ8t4yoebCBUg
cGa8mEP7pOgPjjY7/uL94G8J/NADU1NFUP0EI5FQtz5dOk3yP4q9HX4C2LNJz2WO
EAxCPlrgWLnU8PVIDQGe9Qbq0QdmhJmINW9vL0YsX+a4OBofhM0nqavfyYrkmzJe
Bs0NFAP484QJSNBjK8td2447Tpa32vikawuQ6y4stdK+QmF9Dduan60CIjIYl03/
kOAmGkH/JNdzun3S0kIxmbAwPEJrXsh+gKP9naZ+NY/eG7Ml5hc6ue4Z2UjWatMT
dduIERQIsp94uMYdgH0NFV6K59so7PLrx7MT73tpBGMYlQMCkkBZSbpHaIIIo9KK
9npiw751w30oYIE3Q/aqjRY5FOVeoZ5M00AyfVNGlD/zxjpiV15abpwG0tqy5NZi
zxRk46D9LFlBRa41Te4HLGDVcFRpI1UwUWROj7j42nGU50JyloTdfVO7SnMZ4UfK
KVpFUmhymzW7KRupGASY3L8OiHnsr+lH+JheDTCXtBxnsaqKX65ciRv8MCDWdGHC
n12yItbma0PwDOkiMwzTx406newfs+H8mu3fDiij3GteDHhj6QhNFUCX36p6b/13
N3USGZ7WYw0VEZSg3dMHXPD7BVZDWGn2NrmTmVlzadjO0rzF0HeioX8CYD5Y/oqX
7vGxpW0WWg/pqS5JAR+P6Jwv2131mAaVnpX3u3vWePS/SE/V+Szs2n6W4zHqiiDA
1A+9jgsJbbKRLNIyKcRnYLK2FjEmgDVkqnhbEH4ZhGmT+zSBESvMjMFNQXR4qiLR
IlWZaX1ls4LhOnrwSbsp0c5cd4fgVA5+yRjuij2yFQxREfG019gII5NbzJghZK0b
xoiB+n7b1vhStPNgdhIfbwrNUkrSacHaTMRrSUjtN8W1QdtVojWq+gQxwd8wPR4N
Q/HGGuy+yz46drzNrs0tnWkFoPgemHRidul2+0DLZcPXYUxYe/IA+Kg3EuuzWIzy
U1Idv4y5ehfQth9d4JEwRESrsScrZWUOB5crQVo6Q8JXbSUSXxxzg9UALN4boCaV
ZqqZ0ji6dTrzV8aqtPSqjiJkscthgx8N3Q7rZQ4S7bsxC8SIoT47WoVoYb1yC90h
Zv/BcIIRrBydKHALMC59GGmeAS0BdP9c5kvam2dt80TKbU7DEEDmaO70nDQ70lt7
HJ9XuwIOamWb20XDpc2xAWJYERs8QmoizK9a7TPrTIgwTJSKDTRMJf0JgXhsI6aX
WO1K4o0ByVjW2aJi8Ch+7+WOVQdPcCB33dW/uNYjYe06AWf8/ZgerO8D82UIgFma
F1eco3YDnbvMSZT4LfY25x1SbLLxFhKiEQSmadwCbj9Z090hSsitkqCo0YzjZp9m
WiZXebl1ZIGTIb1DSBZKiKzI2MvrhSvje/EihTKCfuG7Pv5Vu74ooR+LPqByFaPP
1/N8JrM43FXLO7BWeQX8ijE0ePZ0oApUGI6ImOqle3A162I3Ly1U0/T+x9OotIPG
RUO9BF3NbDBksbAx/KMXH7+46wlBcAkn4RWtO42YUflq4Cq3h6+O1uSTk7zSj1mq
nevrDDrI6VE84Q66NKl9xU9xsFDVVNBPebrv4RYyjeG9CURDDroAp0Mjt/7k+lXP
fjRXzACytEvViHGRid81BW+I9IabgK2MPNYcj89bCQkFm40YdWibN0xst0Ug8VBz
iqcZ8e1JaMtqwzr5RdaRR5Oi49E6YOJbpwqqw6hswrULtOWGfC8PKyIAjfq+2afO
1rYNTKrqZct/kDwkIIi1TFByI1oaWskoFzJm5P21g6NydCgfnlnl8QHJ7QuffVXf
+OYE5uorSuw1sMM2rhIWB/uNq07eXmVQvK1R6h8L7ZZcVFdMGtaZ9xeBmOKKD6BA
KA/nmxdK9Uf2hFYUFjvbjWbub7cvaEm0xWZZ3XsdmT5SPozwiLbfFAkhwnNFDM2G
1YYoeQWKpIX+1cUnZ8UoIqkeKB7LEYoNoWmM8VWcEpmHSNdOtJoZlRFkNkb37Xjn
SU1XwjZDBfHi8/A3BLH2t/m03SebOkInN0cIum/iJD2RyPNiakyMv410YmwuQDkV
qOj5lnRa75WjPhwcjPxrFY2nQuGYlIQr+beV10l8GekKQtv56P4OQ6mwxD217Uek
oU+P9CeRWVXlIGsbLcSB2ZsoADAWcO+Cnb1DrDIWvn6bJX1voyqwXsMuufPYEvk5
A4VPYGyZG2H92I74XdabSmmjTjV4A7xfRSEC3t3/AeGC82uFBkpzsqBUVSHeR81C
Xkoxnsi7dHmvfn2QkHiTjw/AzlzmtkABWwYlC6YkwEwjF3Xe8dqy4BVbU25ijxy/
w1WUAK29JELWLqwrC9cxabyjvE/nBcy+tPuXRCJedIV3iVH4PtMw8LH5uNM9OoPe
vVY87M+ps89l0REYHJOKWbquIB1fojmrRLg4hZobDG/DvoVpuiopyO3RyvBIXU7Z
BcYS/lQZyXh8lziyC4Q603rANQCcfTsneChD2TYf4mFzZPAf/lISi6X+68G0nUsA
YFItlVke3GyTM7GcBw3pFrIIJIJH2KSkGCaPcBSeSaYNdNaXQ5p8WiPjAmTQCo6E
cAi5iU4ZcMKZfezzPqmsP9KxhgonHYp9LxR5Cl8NgVqc2woCmmFfP44wK3HiH0NH
hiLBFvO4UWI/qLa/KsGB60yMCE4kbgjz5DcQIYeeyKDjoSqhIUBNi8A1RaTWapb1
KMSeRBz1MFbPkLCcYuVhs57KyFcgJ0kFI+XvpElUawhIWksJtT0BjdZCLWeGVeFh
ADT34IZBFkzCDzmutBRKKhKzu7aQhdl+gews1I+va7brt/PdnxzqK4zKpULx7Skt
nmmSn5O+yHk65BNTaZ2N0FbAqVt13IegqJ9GHS/31QQx22CNF+7L06xLgyG2Umwo
XWONw6KDC9vlVRYxD/xWdelRQa73+ldo+wugNfzPUjmRIifuuWc/lGzaQQCIR/1b
6YZB0+IAYt0Me6NvQXstdHW5XdHdQf+H9RZn8AOo7GKjy+7JquKARYO65V6fXDFA
QTyUmhXYtbyrdRzSludHGZQJFaOuepsfy9dhxwox8vM6d4f/of0hqHiVzjIjQVzL
i8banI1nhwyFvWGqvPfUjv2p+oKU3ehZhLK25OOqYFm4FIK41vy/B3Wg8SAv1tTR
vVnokCM+uAi4E+qNtiDo7k6NKXIP7Ls4rygWz8EuOjKMCUR3YgNzKCk900e8iM3I
aF7r4E1rn/NpqzWqd81AymsL4vWW+xOA3CUE4FidV06XklrgcgBzff13zadNNFz8
HGBF0u45Hc901PJLMDEId6EUWX8TndzJDUzkYJWhBeSm8fV70S7dFHw4A0dL9huy
n33oquV93DfN1PjcWwLh0WaPr57aeuN7LPhdumSEUrhkin31p9BFj+GnstJ/vVOD
b1ny4zZBPtCNYMGj7o/nP/29131LIRr0lKTQZ62firb3N28ZGhJ4QETcTqmsT03X
Cot7eIsJIL7D1mzLoX6eyiQW+ADTnzaczc5Tq94wADnQ7gBpHI+DNNeVDnMGSXCh
CO+3YP6Fi+ARQleh118Va1ipag5jaK1v6m5fH2CtRXTXq5x9VXn3YBu3hyUgs/dg
8PAUEtLTB7GA5orvQ9lt5GjJafPleb9haw5bhlJiVK1zOXUWKlEKvTHgYZwucDtd
SzEnPaUF3DwaQHQymB0FbPjHzDyYYVuaYvU9QsqRk88FUd2P0yZrb3ho3M09Q9OX
WQI5h2lmW5/52TzVDvpzcWKrrzN1V+C37bSMgUNoD/+WfsGWIRIqqOD6LlFkJV57
MrEnuk0S5G6QU9ZQdfz9P5R0R50tuWoM/H2B6ukVcD8Ipf7utaYvLB1zN/BHYDi0
1uCw/VWnFuFQ0vv/401ptg==
`pragma protect end_protected
