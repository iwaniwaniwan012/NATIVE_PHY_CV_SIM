`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ocsAhua406tEbFoOWS07sivx6QTXlzfu3fRpvSOU2owDiWzaPXaS0k8y1xvYJ45B
LUu5cJGfN3Mz8b0g/3hoXcIK6Zijm3d8GYVfDlqFRVFqHSBThJAkB+CQEO6efwLm
bkYnmbn6699SdsIqvpunvDBNR+/fo0uPnox0ng6p9lg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 174144)
hlGnQtlrdBhG074CrlnlAWEYhMl2/rOAB2PkIOh2STFL/t2xpS5368SpsIrG6AqN
2WZDFRz4LJosyNqBNTajCWWmTCusNHs8bdIjorQq0J8za3d/83T0RMzU3SgDBYQQ
M78r8ObwO9Kbcaf/GMN2OsPhgxcQiWVVMsxrYkN2v4qe1lY0r3WlvIWD43ifQYhW
OyBfiN0909jqovkALIZDhpZrecpOncW+JcMVff5IXPU/dfswYwocSlHRVEh6zTQZ
Y0mFC8+xiNkU61BG3B15OwCMoftsZnhAZDsKIAiocCbgEsgusdgnNBWCnuoXmUzE
uG6OyiUGXEWhZztktyqwNhGE3vRg7lOaec/NUxiHwmLTm7NFH8S5SHV2UBVzONZz
vtSC4FuOkSjJNbS5sQpnjzS9+AgOH9BriJ8EIB5Z7KiqeLtKg9nPlsZCmE4o2eQA
1m2is5QkBWUb8R54WA3BP26Dy7E6HRf4b76tFhUF/AWRU4wR/ciVkvsIXkbiu0JI
gJtSnL7hc5tGkKdm2tvM6FzwhJplE+zqU3SuQ9zdt6u49s5/p2KtCo+3+GyKQ8/u
bTakRs1ySjZYPfin3qTM77ZbEu9PMce/q6Qj0WEI/FazUJm62dH1VN0pGz1gBMkm
GaFmcUNKSIJX7uhHSFBgGdmXJ2+c5P2N5tkcC/40/QX7ba1VyzuPLpzduynuSvZ8
W8J//3XxRGQXNQHehbEurxmVlBc+IGf7mBangcgzeUlUJuCAlO407S7kRYVsDwS1
znM/Qbu9KvCy8EzlhmfHST9ggW+3hZAr0dH6z9YV1lDIHVtvmf+lnVL2VEHzlCxF
M1lxau538AyQH53syvFJgpmSjQ92yJkJqCwjem2kwtAW38e9Zz/c7pUqqR5B+4Ml
blpR4PJs21o0L63iyqSaJVf8BXCc2wQW4Ibj5+d6NE32iiih+HnNBEYqq5e3n74o
cBlUSnAeZjnAVX03ve2QbGd/ilLxqY8oUQCUf1C8xeRIAKkTgdLNJOvC0/A86XRl
omxzEaeA4/wLL2n0HlPRvlQNPg+0QH8wVWPEbOdByyQ3gyoaJ2wwJndPIg7HCKt5
vpAvh/ad5859i44H2a1FACJWM7nF0xMmfHRwoXzP85R+LiE+I+81Vznml0KUWop7
E2uwELeeqjJkq9svuNgezOUZgx7QPlQnYiBvq+raaPR5EtwaXaSPDoLxx+gKEEol
ujJS6CO0Y928Hq8zgQeSrWxmp6Oou3+zJoXrO9feo8ODjAxcQm0bKspaCFNoseMH
ewMYIfNNXf9i/6Vduhgt6aKMN1Xth3fAzAaNGX2r7/krVXWM5QLqCITq3ry+jL9+
+3JKsRw1ocksELnAVHcXdbNGPdq/oGfY5pdBGneVtyaGD7QN6l04v30AuSM3mq21
dtc8JdPUVXGbLVFL+1tv9crgLSafHEt0q+xlBW/r99lhratDoh4QerseMv6NhyIh
wj69V7khr+inNYidqwQzMYdOwbsnFFKbrylICzoadV8tjojJF1H2EdtA25Zqeb1S
IHGaWKp3wacgWUE2q4EyuLXMIl5tHaYkYaf+6fER7k957CbyYATe6IlFjl9t0mBZ
i2rip+RxTI5sYVR7T3XMJDM5GuIQ+Z+WTFOjYicyGgnxMWPjZTMYVrOWo5ccWb5g
Uj99CUvKy7fcnCBjGNatTSf7Kf4sYvzuF+mDO272cDvBq0n3YqZThMaD+SVA7yAT
+acEEG1lGJF6dFtZzLTkl0IH9n+sMVsn+NE8ObNG36kutP03UAaUlwuSfZggaN8F
X/GwVGCr/7K7vzAPonkJoWWjeeolxAmxsZ6U2BpjkQjv/DGerFMofNmWC3N44fta
FIa4j7nnSHPIxu4NlMIPNQNYdsYu1WsPHdn4YKkIQdIQ4zCIDUWoNEyW3KQbsqVK
uhLZFbIHQepphDhmV29BMTbMzIG9WdAo8ER2NnjBshWI13Qw+2RtD8VKtytYG9QU
UvPJzPlHYBctRdWrSrm6jehgIfQH94NSRfP5RaYpqQwCJ2Ov1QhxUHC0zVoX2U0r
g7Bl2GCfZJfXOhQng2WeB5R0J47nBPCsP4UBqgOmFXF14f3f1MTe9XY5/4fJqv6M
q6UC9UWcpwiMWI2+T1j89VZzyT33GAtJ3+MvVkW4K5OFKVJau6YzG8zi5n1swDoS
WqCdSqyJYdKXJs/hned9EBrWLx7FpEKM25OihturGlLgBhB5pfZSu+eUwf17bR0M
R1bhzJtQnHxkgyQBkiLP3cChRTMIQgjlrmBBRSfgxwF3AEaGFmqQvuThkclBe/xd
ahcUWcPpncjzIo4lm9zAOCR+722eXrh1fgLsstw1RKsYaDXnhAayzhSVMVAwAgFe
LO5w+jI3kE6M4DQzWwqsAP5Uhp28leIdBrCSlnrAKQLwiIvkJirXOPFAbcObz4+z
RXFrfTmMeFnVWcQyHJavUsrdmfCW/rl+gUifwALwGz58Ghm1y2+ef1E8ExgodSlf
kUb5bllmrhRvQ9VHBPoiZlVnBaoQCwp2wgnBkaS296Jyz9F/MF0bcDf3gYC8znjx
RNKmaJDBw26+kDmRWgLGnS2FsReq0Ucc59nNHZjmRM5R+saDrVKViGV9PiaI5BBV
a1KELmfZWRUg3pP+gx1l/7T6DwhqvI2Om7AhwpFpIj73e/uZJtflrPnSIi6CGRUU
RJVps0LVCObima8+IWtZBVhP+k/mQVj8dayZXbcIjcLKiRdsHApwiOBueJve3xQZ
zlWvzTJTePG9veYczQWrgDR7tCi2gZR3JO+fR7n+r4aSHM8d9tfXr8bPcEaa6OSR
kx0N4bccycg+4vuJaH8r7AGdNKE1BTAgoD5K5Ei0Do+WSGvlS+Et0NrW9tVE6nMX
JLGBphoCBSrlFRsUCUEra26mRvKS5K0umKqBzsiJ/LNIiyEYqTBnyKkDLYJKvj+8
xuJknJGhG0dV0+NeNxpgYRsY9sJnvcP7f8HjvaQ8Q5xAedloA+Jx/d4VOx4bjzWn
X9yEZMRp7Hzj78cHTbP2cNPvMkLODbx0GRtHTVrPpeOqbM2NDNDaNgTKjk1DaRiL
xSrV1kTFb5kr1vUqYRb1yytg9w9ljAoYiQ6/aYxQL8dGtmB8bEzH31jutlHz4ys6
sVBXCy+begQ4Qqe96nCZEnF6Kw9LW15FpwmfBCnJbnxYeZ13ZJl67t05yD/HDDZG
zRxkoAkVp5zfD9Wb+tplNrU+9xOE4fwMJojCJOqGVjNYermN8dGhrBmw2XFN0L8K
svGwh8cgjmPCs3Wxcixd6C/9aLBixOsxq1baDiB7x7uCqncTbBIruen9sBmiNNr5
svZ84gCeNnGPqH8Z3GHfmfPv8Enio7J/JcdEYKuyqR5nTUhj7VM1G8VnjzK9rebT
nt1++fu4L3WHZLHwFSK3neuPmFxFcjtgdHRymVKrp6WJR83flHmdiLesVZqTamwl
iQz3xsCaLXKD5f/wsMZuRk8jbUDxXkB63Zz2tf5I3RnlnemwBQMSTUM7pFkKN2mV
vGmrh6BITVzRUJmx3Rguzz/hMUgSnPRoqbqQipowrCHPmcicz3u9QiOUeVpVEKVE
Rapj+faqvZMb0BHXNAcIMtuI55d99p2lCFoK6A2Hi6abbVhsFtn2DaJUbWD6NqqD
XrQeXv8ciAl7vabyObI0jMvoAFvjHWRGG8yJfSGaOAlZaof0CTVmRCMotsRT5JW9
Wdwc67TZYqHaU8o84g641svjRo0o7srklMvyTKbbUaoE5p8M2qsciiALVelLf8bD
rb9SbanPIlKva5VmIMPH21n1GPEqb+Qf+bJNEARaQL4IYKKkhpXi0ZFfY5TMBZZ8
064lIxzi4KcXZdD4YdvoPyJa0mj2H5/aZKs8v3DykgoJb57PwCyzdybKLN6K3gTu
QBhSDC9DbSs1RqoRh6P8eVupglj1BWQ1qtcvjofWh+jttHNqJrb01LedtsgTeCGF
iUayAHO+FGj37ZEi/plWexzQ87oSeTHp31f96LrdTr3UwbkkQnLvxL59qzZx7oNT
adbKwxe5+RBDjVH/vITxkONm+NtF8d3BEOCgBgdywh3tXeYDVE/O0S276xQAzfzN
sTy9CQwuSJSEcEKaPCym2pG2JIv0IJ8Xl4LTAADovLQo3Gsk6vrMgBfI+k4jsnJ1
CLaSGFGymQcEEpEyEVxciufRGxlAYTx7sUxcq+qiQnUHEp2JcIHGEaKjijcZ3qfR
aIHaLaisk0NlCAV21JXdU8aDVl5lxS5HFXhY+dy8s1xtCi6CC4l1cM1izeuwHcZF
/w1Pluv0KdQEcnAG8VBQNF2MlbmHlQy1OgO3Ql2ez1ymimk4m+945T2gOxJ3QAzf
0FAdWSrRJkvNm4CoyyLsH/s+TXWAwlTX2dNGoJ89omqkXQcMdVmv023wbIi+0doW
UV/uMRpalYUjqUkhjDJWmhxFfn0DO7QbgXBEDbTvKLk/HO2DHgNd7bwKHavPYEZ/
e4zR9Gj64/uAKTQuZ5N4QK7NkesjgvihZ9N4OAVfc6D2US9Wsxz+SMBoBpgS67Er
Nljeh06Vbqgmnci5UslJ61wp/qdUSFo7Q3pPh9RnMBQAXFHBbMNDszm4HiD0CB2x
Wnx+CfVXoG2hP4iGioyuTKLvCWAViVgvWpWL5dIS1PeHxhlyp/KOGRuW4TTU4EL0
vu/G4uxupNvaCfxiv4DHdVs1KfqB1WPAFlIu4bE1RbqG5GUNwzejMB/S2lLHBsdV
MqbHkXxTQLG+9+GSsq1Ew8exYpkCsvFDsZ/A7GOY5+i/L+5Pv2A4WxgC4Ay5H62l
D7qMrvjYbFvuAqaqOPKeAnY3T6SF6jF5XQWXWHHWvGza+h/VzXhCTo7+f82vh6W+
HHicGvBoVvxj1PaQmFRXXSdvtghHZNgWei2Rq8oSHK53lJd/SNhmrqdIy5q7bna9
x6/Jd+ISoTAWfMCI2W6hc7VAMN+5/XYKHuWbDVaTsngAmbRC8eRv4pa8E3Wh0TfT
idt4rOxFtqmzG9qdXtRMIL1Cpe4C85U7X9DlzX5RtBvT+m1tRZ8gUQniYuV6sZA5
wsb481wyAcIfEWoE7lPrSX02DF/7ZgZXB6FR7yO0SHmnn3HxSadrJfZwYk/c0fGC
jfsaobh8AybTZnLoEamH8JEllgs9rQzxQJZIs648jpcIxBJVBzMLHn9/CK9r+rO4
h6YkXi2kH7Jn0dfXQPQDzhNDiXXsTgpd3M0C+vClV3KKjpiXbPoh6hgCHjAyVE88
8m3p9i4fBTCybbrWBswMqfmJ5fAxC5xQ4JPGicIfHhK5F6683XOPwjtVv6eua8JE
gey+1qbwjIrXdOMSPq18NZ28jU6Hfza8PWqyFlyah8+n8UUWvW6Wurv0zUeGVbjA
ph8P7EP7wvhvsfYxShVqE394gm6yv2bp7cVl+x9TbnslFgFX5/0EMMH7d/lH7MS9
Wf6grlRLTrJs17wxXvYZHFD14/AlWLBIsacwdsOvuidIo+lduxaoVoMMrFwSWM8A
s/T0QhpGZ+EAdo7prqd+lc6AEeNVvPa3cZLehcApKjFc36gAi6Gw2+dgWXHIdAbz
J3J/RYDocUkUSPa3308f5nDMUIqnnfoZ1OxYD8V1kNi3q4cusmPqht79Up1kLTHU
vQPzxi4Zo4lZhnF74oRh+s74xVXa8YBfdUQF00xvUae4+gENQ6vyjAfdHn0vjV+h
t+t1oPN7uPt6rQLNtQ+Fl0BVDQZqBqpgHzDe0hoC6KnkbiXIKUXdsqwTsH9u0gfT
HeQWGnMcdKybZWEESIkJi8aeegSiGfV2tgOjLURgZ2tWkudGrzApppxkpNWGDjDd
wtrHWsqhS2SOESSAhQJBKuq+Bm/4Uc2US4JRm/P3zIMjys87rawM399uxcIj5fgY
J4fnNwPOhFHyb/d54BpL3Arlp1X/BYFSAQrh+c0wM3ijVZGEf8BjJWll2OGNbp/m
9/s6Ok1ZY9i6ardHAC59sZqVbHxNrbUvXvMwuo8XvOuIlKUR3Zz+ej9+cy6M+Jqw
5OAyz9HA5zASDmowsyA+haDd71zl1MYCyk7cdIldnJcL9O60qxs6qWDrM4lIG7ki
faCal52GbJTJZuwnHcEYOZsw5HE/eTTF+wmir9pHiLP0KZqv9wjxS/0WhdMJ5PfP
4hMUFxzN+Y+Hg+vH3arTSD5+uAoBz/+3/1sFD6puRh3pmGo6spnl7hsxWp0RLk6V
gg9Bc8wOx1L5HsH8P4clQ2Exf6FjgemMvwbmFdlipd484JKgQqDYth7cZsZcMwHW
5JiO1G6iVP90gb5hPqyXmeAWxBN1dSpcfchhyTIEji3bSfoaX6ledFH/MJJbZ6Ke
NELzTUg0tKsOlBkv40vtOIymBori11IlpzDmMs18lGM8nn/KyHhqeN63byJVSpgt
g1qP7wg5el9XX700RjXS+CVz1EZ36bkljjkw97aHYqj+BD5SGYuG7qn0x5PxMUq+
EWW1ukfPkHbc4VnkBBSAN5FQ99GYZYa/tAIV7kkoTQ0hPdQ8GJ4RMlGUS2VgZEed
g58Ad/QJ0TDbl2cQhfyX9SK8sW9eBsiX+Knz1+6ItwR62Fmf28JDsPYGk46dyq+3
t38zzKvwlWDbWvABbPkQaSZp+VHTNeSF0j5l1TjWYSQZVRqLmR7WjaI8UwAMyQ4F
5eH65UuL5sEgN835t1OrcEoRiNlOss9UQhSTuhWrxSmIRRfQpV86JdSl4Fc+p9R2
gdWnn2tOa78UlZYoJg8juF/H79XPHZTEZl/02K71/mIrPD5Q2eLpJ947wZ+Ey1h9
bGNQ41qTbUjRFnNAb8CJJ5vYaJN5zECwKJhhja4DTB8hH7IHJoswurGkFR6SflzB
eEQC8uMIknseMqVNgT1B2Nf4Kd5JWpcw/kyUL99e2FuA7bfyEzseZEFhQGAR3qZE
XQAcVyVR5HdLVT3Cvvy6m7Bl7jEqPnRHU5wULQcT2o14OZuBKtL4hoyw8toKOejR
4Q6Lv0adQaaOrh4nS8HW3C/2r/kDXZ8PXxzQVoebSzWXEjYNVAfCYXCc8cc3YPWG
lsaW7HFyELGMHfGdzv0m/BG0Wgf9HPp3H2O1Sn/YtjzS2/9xAlK/X0IH2T36NiRJ
8GLJnE14dhab7ttJ1pdPJPASpU/W4cHPLZCYyNGgETNhHNBrTTjWb7pxz1fjIQVc
NcUAzpKRndsyaOVIhjZlIz7cejiilINeyl6pVTm3iq/84X0TC2jZ0SFRbufOUOMs
bDULFxKm2t3ejgWo0mKaJWGGvlr+li8qwyp9zJzdRQwOLRAzeTj7YlXPx1lEEn2V
FBTWo6Er1G/7JOlZRecXedutluPYaPBGfczDR4oM1K6r355o48ZFeDdNUtCTfJz6
xCUQw9zmwbcTnUfz48FacN30meJLgmzJKyShMBk9K3mRcro3Y56YCLmOFq94hngV
hX+QGNRT2ZAz8EY44zkAXW8KBHhH1vscrcsD/L+/rXieI5eoUpSAfOhXjWcih4YD
OHvPz8SRxGv16OyytTKCemIAV1wJdnbtcrylSGfX5UazIyz30V1JJuao1tWZthi8
CN1BkkCwCgp3ZaUL/FnjZcALG7OqVkhYe4epFB9tDMIacl8CAqMHd2cZgORRttQX
qE0Vgm0Mq5DwrlToOIRd8Wh4eanPRbyYmljnRKly6tH+8YHqM9bTVeXH1ky3Pf5U
Qqv764cremQaQi8josnWWX2N80zuiapz6KEHvUlPBebrhTC6OysHG3WtiQxQyB44
UvjMD/VLRaJNBVSdmbP/W1Lhd9myhBRQuQ9WJSIBqMJt9QJdhFVeT4aCgTk41zHV
DbNb5nH5TJ4C4PV7y+n7DSyzsC543c3oJHYudQBpVQtqeeihQpOq6W7jZ6WVNZ4k
mMeixtZ2jm+KYih3o2eYiElDyfRJUEo3RqbWjPHbczEO44OHnpSIe/qNVP1F0lVd
jfboKdibWglklPzwD9HmDpoWzxed70efKAnGhMZ9pgFGexoeOGUCfgR8Ay6z2+DV
pMPwc+Re1J7oAOv5yde5tEUvrE/3q4iTh7+q37Q86436DIjyCZEQpTbRj1KTNyF5
+Rh+uafaLzXojj4eQc1LOHRRNC1iQQB4+co/M/gMOXwdhiDqrZ0nV7D8g8+JM206
B8qiL4iBQffhkh1Wzm0zp+YNpNXKzUSFfOkESxWh6UCd+NcqtzsE3hGi2/xvJPY9
m2Up5ZDMi9mNjTUagJMaFz/xuQujEbGClsTlRNWVccXiMIqCspX+Bk3/x1M4j1nm
TghyX/akW3x6Jd+WQuQJDfBFbo6dClrtHj/tt4M3Rb48bUWfYBi/4nr8mc2Jd/3b
0paMBc02ijc6gl2VMuv/ucB2949cjW3+/6Nw1K6HPiLCDTcAMzwQl8lusATP6HXY
ZElQchhTcWLPcUEYc6LglEbN9WJwHENQU5I1lZm/ywbLxDSp/BH01lM4DoVEHlts
snX+ADVdzo1sC3Ko/ZUp/Z5T5ue//gReSY062k9daZ+yCkXl6oQLx8H9jXo8Xcko
odQQhpZxOElOYuKyXGGcaZd4xl2S8MKFrBZth1zndrB6lND0KbSaKqBMy5qIgsYe
cEyWUff8HdXnlFFrkY1j6IM5XQiIVPdVvZkt77QrLiLsX6pdS9Igz53o/mEAT/zr
WDgJ+0mss+yCG4A1G7IA3QapigAyGU43Q6GX77P56EEromN1Uk7bmLiJpaSA0FNp
DW2s0tRbcJ8skZnanXgPavp4wAw2EeqkKuaJcJmkQTgdWRGqOUXq0tBgiyR3CIMO
EVla7xH7yCb1u8aSBNmbcq/QhBNT+uZPoaPSxIh/ODvyt1DFWBKADkZe4lXsu33S
tyFn8FLmG4ZcHQ3zXcqjemtLlkcI9SoPnVZ+OPrOplOFgBmQggVSbnfdxYmQwFbm
T/UcOrouhSDNp8w1/LLSKaSl8Rnsfeh2pfhJMOOu98eDwflSRFOFX35SWyywQW0w
quQHfxJyLEDnWf6rBkKOxlvgXeA2KmmpqWJs1byKCR0JQ+a0IK11Adx8oXpmEDp8
gVT/zaE6f174eyTIQWmb7k1FKFm48EnLgPp9Aeb9F0LA6x6dZLkuwLnDa9iy2KmY
/iZcmbCju2+KWRPVaV8b/b9TDcLFU63WfzaF7AhtzX+GONS3whJ4owhaPdw0yBDp
s3NH8Kwi01E/a/X6h6v775F9v/ANuxb1btSW/NfQJRcrv+ttJpPZgN0APGiCyqen
Jyg8s7qaOwiNRrL/0LbJVMciPUtfjdbDOInoEaVtiF8BLonyXPgumYMvnfq0jDSB
xXyVs4z7m2Iqsxme7lB6S5YtIQoRXKQoJGEoowDhl76Ze4LxgLYTsd+jnBvFXk+Y
7RU2n+kl+OavWgH+vkKEqxPUi9ViTJ3Lks6Dv0ZYGkMOuxfGnTFKfD0dEYuEtxc1
yhP37Rv347lQONzl8aC85qUJSvTTApRYBY7AlDAwc94yx2eKUnPNzC+IeVUQPODV
d2XutrFwRK8GH5/gr2CHFkmNcBbtDAfSUf7QlW5xOoBx6F+2svNQylrnmtzrtvnB
wfbEP0qlnMZtgnDJn5GKGY403y2cYbqsPNayrB6jiiBBvSE6EkUZtcr3c+HEHvGV
w4KGSgwUXiMOmKDxDJsrvNgH97gROdG98qFOTVwl0FjBK7xU722xWCYFjw1+C+AM
WUXCTaPHUH7nCPA2oeQrMtPDXhvHhPunlqsOYk8WOYo9mOUsvZcacXTZhkpuPyne
KofvqrWK1/pN8nihaHNmh+plhX9EHDjpcZmFnjvlxU1GD56W3TDbUpyPJZKYIrTt
DQoVz6Y+xVnCNpbnio6iBXQejQDunsKnV1H7jUXiCDzBNaWTgLtCQJ5PTIkMX5Qu
rgnLy1yYwwyb3NhQR46/0fcmUVdcwNPCwPBLY5rT9Bc9jxIIuv5BOxrEFIEbMQgO
5Vxg8WV3iqSifG5YMYdSQhGzyJeBWvDTmze0CkSAgg/Us68FxfrUNiaDsokmjNvp
yLa98wumkRqHN6GlSfwTiKHzFTDKHLvawWmw32kle6uciL8N9lE0FBfQ5RbRBiTe
Qj+XFGv6YkfGFCj9DlR8EZLHDjW0K31s1Em8pK/+5BUeQCXgskQqrcFs6XLOJyQh
PhL+JbuCdeQM6Ifx33sVL3LGy87kZ9Zq8XfQdutZ0GfscLQyxUIugq7F4LjhiU8a
601rpex5zwo/xhc6S4C2hTlPny2qd8Vtom2fXkkBGilNOTAFLEtce1KCpv0ntqJk
z4hAOpqlpI8ZsVuChHQ8d3NVXJf/TTJDgiwBI0J1YAkYoRoePJj60e3gaA8TRjpE
Zt//jZMegU2T3p8u3FJYuM1jWr2ScFQd2zdSthgNmKwsEKWh54lolcccWpnGFqMd
fKHUpaPIAaybi6s58x2vqRbU0oWBdyRmswQNLEu6nBGgOf77Zw33rBGDC3pxN+xD
mxUeK+Q2YKIeBU2BnbjQFm2wjnqeqFggO4nOLdMXkz0R+VZPtDS+j/AI7+YnbdGZ
YUTmL8qLYc9I0zMTzyOaMctujfYEIoYT8ecZBYOF4DvKDnstmRnJHxWTBcS9e9ne
2J/3BdfmnKv//LnhL3j5y4+y4bq/9y56XBOlMoQN3FgLb1+UK6opUdImX4CRCd/o
wP87NwerNkuKqTEOldRUp45nRHbNZQeZO3V8lUl5NqM/rRclQLGBX3gziBhODXQN
O57lCntOTSHwaDHV5hZbGscA6mq29GSKXQPqFIcGfJKH7pu12sDnNVEa6JedoqaA
YUDigS8MCB56QQXQ1YCUDheC2K6qiod4YRnFa2wMmJDf3zGFnP0cPWEHiLFypKTg
QwyxqaNsOi3Nh+UcHJW4rUKYqzJ609R6xsG2GcalMydVne1XA+1kWcyiAVet1+EB
9ev/ET2QQ1UzRnv99ErUb4/DIc6pBZoqzEoziJAx7FXroRKbFzSyUQvS6iDwFPUr
nsxcxZ/MDDJsq1IWR6NcC/s9MbnZ4UImfWs3tLcGrF27JNn6YKXryY4/gETRUmc6
Gkqrsi9eOFOpr5B8zCTy32Tm3Dmsmj0JwNpXDTcOnJdiekAGh559RbRRg6aB/JQW
yP7N2djOc4SC7I9TSifJbmxMJPA+LKDkV1WKBQ0tphWjArmbNwPXgfnwFOi7GFIz
VVpRI2mqYJvMmYyFUEDRwPKGbY2Tc6v5dSAFxxgx9a8KIdJrPUtH0OEf5d/kG9td
HDE/+3AfGE92fVwlf7sUNEyas4vnGomGI0ElbxiTiReui1j4Vm92soW/pW4HfqT2
Ke0Slmn11OY1/K99drIwa5fdqQhg63a4dcxxxAtEyWG431ErYN2VSfmYwLJ6WdvV
EpA1anK6fSSDXjc1cIUqs6/rmZ2nFpVqcgoKykP590PX5mDsQn7Vvu06KOrXNh2L
W2mhwYakYyZGUXrlKYw6osmutTnlNVwXpa+fhoFvcBMBnbYiAlAJQEwTwF8DCK8B
OpQ3LrioZ5j8xe+OhxGO8lmwET0LcXuLdDS2+eBQaHiBFy6UCLmkcxAiy7LI2dHG
BPJL5U73cW+2j9N2LeoaaOzu/qBntO7jGy8fA0Z6b4PkZ5rcKjGdEE0FHxbEHZhx
oqfCboWXoFwz4v6EcI7rJq2HML3XKS49IsdfXbV9OzW8wmkjfPh8f4OprMMywTZ3
6WSJD3MJ+uNgz0657i+3FKVlujL7Nk1L7S4U/diweD30OwDj9d/YA127IRIm9ku+
EiZ9S+ftV3wJOFx6K5w0WFS00tzwhGkMZZgmVsnR+Gjeg7TKog7RUJpvi+I7sfc2
jv9zcotkV+g0zwXxFu3zWhNJJFJ+Un3NtnEPZ7lvxjB+URn1SQYvKB4cFfRcl6lC
JulRupbAHIc1ERme5mumN0B+7jIK/kZpQiE5NmOPvvLe6W6lVyB1EpmFfb6p2dEL
Rz6IkDbkL0+7n8qGASpOZmnWP2eDhC6jlWayGO/U8UJAyDOanOnxaQli18R1qYRI
I0oyePYynEEaSfV1J7WhmsT5sy+OwQt7DCU/aKOQfF8HKskjzZHq/TOJGrQnKUji
a0x55MD+RFeY0iXQ7PN5j6cz+NhfkNcIwr4iUupvsYRiocRDAszC4JTmKcUPn04J
5U8st2e7JsUrembeUfgzGyshBMUV/NiEiUXKUKUU7zpmSGfbgrAsJJOYgY7QHlRI
+wzaqtCMT8C5o+Bb2pystM+Fwa0Pxwv8zfBhuO2qfur7zt7bbdplk8QWkZmTsqC6
tR95kdo2jwnvvs+Nu/Q0U4FzxOLW6AKkyOEMq9bsUdx7aJfBAG0na3bwUJjmpnBb
c686be0kZX6i/RzJDgDfJqvvWfAdFbrS8t8lLqkHjtYtpOUz67KHfzSJCip3hyPC
RkZADuhFcOLkgpTBVY48deoDIGs+A6JwnhTCk90LGBRFShR57bzMqQjP8Dn6Hgg1
Tc48C/eo10SwuouvEFqb/zC2hDdTX3cKQgIxulxT0MCs9OPw/zmteot/HbWxQJqY
j/nxPZhlkNOINV8TI4rpNPPxXDNLxwPvcRSbxCb69+HxnwCPgO0onpFfIJzMLMbB
+6/CrQyHBs62S27EJ4rk/+69v8nk3mBnlCaytUwtgU8Yy/ItFosb86mKomw/MwNq
5+3F20BkY+HX5V4Yckfn8Rtucj8CBIc3Hi1TrcYDX2lKW3EVOAY7OJe2zIpuDxce
hhJes7lo3YVABl/DVbL9gBIs9BRrNT5L/7elKQ2a1JchneZ9vydZKfxL9quDT7UT
Y6fttw8VNcH5VNeVXx3+rNXJDAuqBcdAEVC0gp3RGyFbJyJiU4PwUp9fnb3OuNun
wynJ3bvEEVL3lI3J5AtjmLSPHXdvVY8uPX9Zvt5LuU2AqA67YSseYR9hQR64Du9S
W0yCuf+vykz36lxapvF1Kci8hIBdeE+eoav/KNm1epsDirMTlM3wV/7vbVTyjVZb
HK4nH4sib5G7xI0VOxFa82iDX3HDoefrcTtaoXDPps2iS8nxj0+05k6uUb+hGnsS
es4CP5TkwJ5ULB2yycjLTFNm0FVGE5MVcVmPcGuv5JrvGZtks5wIc0NqugQBIq9u
/UXVYLSGYv+BGOPSWy4sETYNuUM5l2vMDVTmINYZkw9/lPHqYeNTZBfeiezo3oEC
2Kpoo2vQLircXi1FDZI0BxwRU++RPvb3OH33EY/xYrsTSSMaYwhblvM9QzEKcBfp
5T8WGMoucTnndTFbgiUHRoNiucQBQB8rxTDoRHf8AjfBpENRw96hXtHOepr4twYD
d8Gag2cqaX56VMeNWXHfE5nbAWg7jpVCo0EAlhPeAcLMJ4cK5LodlJ+RmxJs2Gpn
dVKvDFYFdkU9YqRbTguIAKM0iPy4fAdNd665IWqmrP9DfbKQVUqhWcitJcTziS9K
MC+6tvQkPTUQv5bpyL9ismd+gN+CwinhMgkrDQt7pFa8UurIFGKt2a8bhrzf0lTn
ihcyjDQX77hMoke2/MTJcg1GyKkahGxFXU1jX+yXfHtdSjzMtrkblN5UQjzPLNWj
RUPZiZWwq6hkGMVg3qT/78EgEu/WDJWXAD3C/GPdD+DV4qqzgEE7StlO2oB6iz2x
+xfBZyKaGuhUaET4epkKvwE4OKFkH7xiFCvNSEC6rZKfwEGEpAjsjQCULnbMBy44
E1IK21vdravPkTM+szhCRAlGPQIDb1fgdtUzv7vV+M3HhnMj7QpdhKWDtJLj6jdX
DXAb304rbNZ/F4dl4iQKxyx1BPjr1bqSUEu345TKJDAnDio9LzZWzvHG6A68AMwS
/Ozm9VaC/xWmpojr+cwUT2sNQFKjgT1mG/olHA56mDO0hKzVN1QjqnaEnSLRDnDU
Q8B+W4abJRCJnbCwxZOxqCWEmVCb/wkACeCWpUyF9cOUmZOwBhzTIJrMF1ZZpQI2
7J2Yo94gcI0erGQLS7ihHw04VSzr6UASOsKkkRHImUWXziLrQiQc8oayTETjARbf
kcMOdH7JqhHpHDqPjcEvtW4vMiwUHuQWCCcFBJhtzfW2JHluJsf8SN9xROFjfX/E
VpHb7o05Q2k5lkqi5vZkJ61bETBe6FIEEemfLkDh5D1jZCdkuxcKfb8rQN33uc/1
WMGLglFKzfduHes1qr+87LW0mP4wMTpbhDD2xgKiydMn4dDJHmEdxuUaXuLMUOvj
z+GO94DV6JTEdhe3Lp2kpieRmAdnyvjUucz4ptHgn5RiWkI4N3QKkqJnjQq+zatV
hK1RYm4Ym7yMgr0ihlMphoxsXRhzu8fWPdObgg7TY9pzGt8wFu1T4GCIPh1isURu
qIcThBULLD5eNL5vCUp0Ak7s0aM9d6KMqkoC81IXwG9iJmgw7p8qGXm21ftrp5WV
6EZd+Zwhx1Z4JoHFCmoopfZky9AA7Q1+nPcoXP+Y3GX4ikbrGNv3YsxYuHxd9Vb4
WuU4kMEof5OvOf/0HPMtr4nI1JwY7Aj1yU/A9y3WUUVRV7vsoMTx4G3hlzeZqm1F
dUVx+CErTsUPEky34QB0FTwtKJrzWVADJJVqdu/lG14cLciUnudyFJcf8Hqgsjq5
qJ/cCeeE7hCXlWWRYtB/6IBF7KjW2KawBHK3ju+ocQWZffBRuuRhgFqMTcrwrwj2
SqkIh0FDOVT9mDDW7Y5Z/aAFk4EiNLJlN5RtYgtoY6kncDISeGFRmNDwkfTvSLQJ
MMELErByygeNtg6QPtR7it/2fh9HcBbnKKPk15vC3wMVhRyIz4UDSZaR2h+w0vB2
SafTdO4g23yp9stZjufvAtEuKoXQRHPVAR3e9o+4z7xfOOj0wagKBzrEtWwLIitB
G7DAJ5fc8hnUO6P4SkkAP28PgIV/jxf9hiFV40MtcSFsv2HuBzhhKfYKqEXU5lC4
s5m8KUPQgT5w/7YjsieeAAF1/g8sLyRqgCeru7vppJBfTXQfNGtCySw62t9xD+38
ShVyEkXFWJzo4NUh5C3c+U3fVifB64Sv/lDaNIfC5jFWE2+BHLozpnFrR960wMa7
SGlpKrY78/Vn6ECVC0xnyhmQvlq6t4wBmOUNM6odxGhyjP0rxzIcFI/RmolmhiQX
Br8iDIf6WQcJIepbFDdeXJE6q831ueo5ofdW4mthut6mxgUl0gyrW8v/w/Nic7AU
2bN6UUXxKUr5iOfMt5MLiP4jnufU7AY7tDERkFpavML+dzZdp7QqDqkVDgszfJ3S
uBEE4o2KJ0Re2VfAoeUYRi9AadrhrReubcm47aW81rVQ0R1disVUgMbBufTAG820
FwzxRlzYSP7fRss2QmAf1728ZuPMNIVMFuwWlnmb67BSzrLyQvK8cLIHlih/ZGv3
bNXregwN4FOQMxuOJKOMsdITq5DDAdv5EDCj3Lkqff4rXy8Vuw9bJioBlEwDVFgY
EttY1NJI0UZimIxlKiJF0KHJX4Aw+cNYQ6M6+KBlcCnvrLsOOQQYN+o+FSIiQVJY
pP03hD7gKPM64KimgANV0TpZWd1WQURy3bVjdXaef0vKBbanZK8vlVzjIe6EOECa
G0l+OQ3lA0+q5iUQ/8mYPgIZLu8PjBkhmWN3iptv5D+9sy2amsch77C10wcH0bHn
8gN5qO52qoe1EbRQinlZBmoABjueHtXQlrcRGdy/1cZTprJPA5BMK7SCbiz6yOj6
ovrJXwkcsj8QRENK4MCkTtN1/2nvkIp/3AbxtHiJ5HOZ29Z5JKGawaXQohHjMpKd
6/bTmYvGW1QNdm9UcpyCUGrIZvkyLQDaZdX93L1gwlHei9SAH1ANYYKOczHt3LJV
yMjqx9IP4UFbpbAs79rpWxwz7VBNhd/X7LfvZM/SWqmSyCM+TRUPu4pi4YeCh9vi
FTl1Xb6bn9c6y/STpRDoveEC/egeFtyJ70oF/8UFWkIYUtOtV0XZcOpK0nqm0tzO
jnNXC1OEU34ZXURQhGDNMxlkpL4r2mNeMna+I1Tys68TZ8ywKPHSt6l479bVDYAt
C0UG0MjqGyeA2iMdCpCWDB5Q+MFUnE4osHifF/Kfyp1VOGgx9y8JVPuhm/aqHRmr
uORQxP65lRI7ds1AnSuvnbG3/z5mXOJSBj/EdDUbrmXgW7LNKwsUW/0HxPmUGpYF
275kituy40aWU0jj9IpCzwAsIDfRyzdYKl6LrgrrCm4+A0yuw40xtXUzCexH62aZ
RB2RCCI4yrUFwM/NV5/M5VW4rw+14QHQTSoQdH4DCnE8/+sOMQTujAWmWZAdgbON
UJRZVsBNq6Jue7OzQWb9oX/HLCRsnJUQo2VC5HtzM3JCA3cinDFm7LrS76Madla1
nSNr6vy4g9JmqZCrMGX3ebolNUhd0d7xmn1gHplhR6UOuVcznw657NGgQNU3A+Q/
5lWLrk72QoDo6t/mopqOBIgqjw5nOsB3uk17CNrVfbfzjRI60oCCigkRBSRH+mPw
5UjwTFIWbyIREDFLEgIMO428WSFllEPgpPw6V3uPs3CJF5Yz8fnesUNi9h5EXrnA
eqr3T1pu+9YtbpQ9WXkYr2t8YTaVrTqsySY8nPBS7tXnBe7RdDYED+bHtvu4x9X9
O5q1iBWnl/0+S8mWDJD41+dA0TNdAe2fpCeMYckhS19MEncCes9ednMFpLjnPCP9
rTVgzog4h6cTJ9WYcP+DMN5ko70OuTyrZLOdARtpwiLyCP53ZqNFxGztn4OF8SVs
9Q2OuFKoKC1pCWA4l4TSZGf2o207YWA82yflmORZES61XkVsLyKxXgygo4UH75rd
cx9L6spYO1mn/8AHiZ2dsLJENqxSVkK+U8kn/1UZeIwlGfzwAzVZ0cnvq8zSrRQe
pznWGR3+oGqAaVbL59vU0hQrfkd+8RhFvk84R+2r6JU2haOmsSmUwryDFV2pk8vU
5MVBZpb9eb4lMbKgzHb745hWame0eseT8yOhexqvD7HkTlFp0ELthP/wpKAvJqJz
lsZXV9i09JXga4PjpK5e8ZShpW9SB+mFzwd/nVfb2LLt3/70frkr3eHqpkWuwitY
Uhq74ubi4aabrTAMmGi1EcJzTGNb0ihQw6jzHRa0PSNIw09yxr4DlbiZmygAHrAU
vcjFJrPCqQGhp+dvHurkV0D+uHbM5mt8mXb6iEWDjNvBV3xHXLnL8VX0CUjk76P3
hi0AZxttrDmIp0ka6c22Fkl4BuWxI+JUVSUJcVsLQNJMe5J6rEE1ugD54gz2OkGf
hsiNDdCFXuVZVBjhwOVJLfYXmp51WYg/NmXEsal3pYjZAfHiGQYzgJUuy/zRwlbB
jd7XfZIPCCX6YMdsYdDg8XoURCtnaKUPguWehqJU351QsibJr94/8qwpA5ruL8be
0mpitEZ7teABMr5pz8L/3wxMHEpbS9cpRKKOvtJwfh89bYOqLiqURcZdF4O6/xDg
rAJVK9HShYfS7lygHEj6KQHOM7eT3bp1G0SttmwnOw5i5qrkQqr8xA89vgH9WxBq
7MwSMBW2lByWDMOZbIpnNnFx+XubPaIsl5Z3F8rRfBsvQ/lPKvF+UWMgNblaCmDH
fOZOLsieq2YVLeFMOqLySLuNDIE36W3B0IqIAbAoa9Mjyr5/VTA/40PYvZVOOut4
ru7whGtsp9x9/BPOGaFMqdDweTzF5l5DnLkTrmVfKXQzL78GzyAfEzKji6ska12f
dhk51k1PgYeQr+5aXq0G8hB6i6ju1o2OwgfdCRedsY8wtrbK3p3a7s3wPn7609hy
40WuIahFN7U6FXTfQVIRWMi5pahuGjB3gCvTlyFFlT215NXoP8/u87LgPdJCSPlJ
GSOLYqqObwKKoCXTuTpQ70phvsSzHiRtikXdMr5V9tQGnPQ+JtXbJkiWdfo3COG6
H/0eWnPwTapyRU6LkBl1djcSUOow5m0Wok6nBOHxPaM8gmgaAVaUKwW5zIXEGuB5
oaV1UVtYeyyW5wahwDXwuLtXOiovua4BD1Rcqt0vmzFxA844vSQKo3j3ZWO8Nnrq
JKbjRZlUevLYUm1z+xJI469hENVWoY2vnseKakXd6Rkj2j7R3JnYO+eUQeY9mY8x
jT7N9GBeOG3UWEP+WixZr8A3qHaTvnhnfj4WqI4ycsGWFpWntTtc+kncIj2gWtxn
BLmyLRTza7rQ3xC3DXO+nZHmsm8NpWuwDnf8TBBMWRY71BHsXb1ddaygebkkWlFJ
KwqdtyNLrATatsoS6voLS8/w1UUyT3LecMkVdwDn9ug/OFoMEWGAeNt6sHDjzEIl
qxyJi9QUViULcY4e4ubcmsiQZgKyuj7z8aYhpxtV1t0dVn2DAXIdQ3rVwCQl8gRW
j9akFqRR84RENrILiNIubLJFFJPfFHNecmhtHmEAFIBlK6Efnb7hJ+qZowZkGH2J
CRRTO+uAHu+TAt9f6OdnOz8zSm4LOtDRp4/+2YnbhfuPtUVempO1KJjNraWGGDXg
6NCCjrjTu9cg1/U/hpX7rzGfopENb6U8086J8wJ9D9UCl673Df0vNzBSuIOsE5ix
U8PQoCGH8sQ2K03pE1LDCCNwxfGaXKkCCOv2Jm/R6SBvhMvtVAzAxCwIQVTQkHNc
OIFIXXe/UTAFqYvN+kU7noStlJ6qYyCGgrWSl7KHASIWBd1bio2hPvvcIES1CNOP
mbz2YeCbR4TLGEUfeH2S3VPne+7n49FF7DrQsvsswmJZmp1VTieZLTykoSTZBDkE
YFRrN8jgYTJjnh1LeqwX27NqOduoeLxGsCcrvCNm5ukQZgeMFkuFSLeimnWfZ1y/
4dDcVtbSpOSnUH9RXSOxddFTT/+ULOuHfmH+WCqwGp7XgoyQQPuR0En0okcft4ay
YUPy1tox/ZChnbww8Caa7rD2KO9jzKG9HiXRwQ5w3ELr6wdOVnzSB+znAWsheAGj
0JoLcDkiaCPjNZpiAdwIGBhhwPVmDe7D/Si86Y7zuMYow/yBEhJh+ncE7eQwys9F
2JNk/NuBLF2cnizSUG80KTN/Zs5URvEceYaCGxbfEV3HEnkKBS7KqbWZFM99jYBG
Rf9rj/DkStfaaBScUnkwFytpqLlfRoYtTbQk41ToRhX5c17NCCmbGK1T8maRUeC0
T9JMemQ3wQIXZHJVRUzv1hdC8xP6R1cGenpQtMTxvoYKXJnMrGkTwAo6G7eiJ/N/
/njaFW1BCkDvamJ3dGzPcoiMsEw3q4HtXQ5bAkCSaxe8+kOLSsZcdv9PKhQsH7Jv
483/JlXp6wPqobx+EpBbhNp60QOZWYYte7kIlPKsRxWQcQ8sVOhZQXPD6l6NwBZX
J9lfidkWq1oEM0HSProyVY8ixWPp/TJpXRV9uE8FdN80gMFEjDn7/untJgFGEn63
DmzLv02Imk7rvgaDYe8NOtjzheKia4QlQ/jWFMAwaWkM5BK4d+5Q3iyrQok+goOM
thHgxsWFhUVZTzxa1f5C2Dr6TS97qGGtRtPW1ZKa4uEycFsX47mM6jVEd4eOjeKJ
ZEhMaO1rNf1uAtD716hxVqco7I3x+4NftXO071qpgxLpSttE8dSohzWHEr/39MZH
sLbsoS1EW1eoGZAUmK8nlvVhYnu5ZoJRMEKQtZV0zxrD3swaWAcwlF7QLdTx5IeX
1kOo708qXJ3E+KKHAY6eLLki/Sz2y2rYyAj+hA0wvfYLX9y21xpD0E+7wkEUaaZn
zOJkd1DnTInhxl8o8nsbo2KAHelNl36mTYLIhrygJrQ5LpKEomqmNv5ztUFmXAUX
MmKVRI7+7e2oRvQq3MRM/tlJbUJpaMyd/IBfC9YAGtM7+0LHzl1KDrz5I9BIIdr2
SCPUc+prsqNYf5N3Wz0lwt/mtfuzP2XDcnt2xNkT/Hy/ZbyGqIQ8Hl2fTyYlG/DP
UuDwJfyGYKv0StVvEKWbpDucauUaSZqztijvQTzeLMKxFpkyzEgrkEkG+0Ez/MVo
U5aBIe0uy9OV1Bp3FKTHVzhgHaDEtSp4lkGNSMYIwbYnFNG/GZIx/6aYRKgpWWt/
mDqIE93vMnts4OyxEGOXPoTso0iJrj8WxBB2MUfXdWhC3B/ZkloELoJ+PmTqjp0u
k73+MqBHihf0/GPargf2kclvTySinKsV3k1jDgDKGCqaaq+Mq/Gor1PGHoPwT+9L
r9JiJXSU1j4Jxs8EPvE1BgfNuC83sejx21fZ0X+owANOMMv5Wu2Y5d/DBp36HXYg
zPUUCOedKrdHcsiGcPGPRBAzGYwqqCvizsx/2wvOOMPEhi8zKuM0EgD5z6QOVfgM
BgSgzmwq8rb4NIuoOh+rSRYW6CP9OOurtC0i3qC7C+eDXxny2DBUJmvLGi/rYFcn
RZuosH/M4hzTLotHCqawPsAabd7wQ5DXh1kWeTUk9acN84dW5H3UKfLu61klYWBt
xAPrA4JVBsJaVDJ/NSgqUV9EjfyT5IJWQ2jmhyBEEsVw3bRLqW+th2kTKOTrFkwM
5ISQsU9pNKa+Qoqhl9iWsi2K05iXS6ZlDHr8DYLbVWF06zXzUxVnZcus7hpk+OaS
PG2QFhPhQnOZlEOh8Rn/J3smBhFQ42jgXRWwMPH5e2N4fEfJL0ORDYuuUQVixrNW
pUb1dpUjAkTVgVMPQOUfA1wCydExe9mv7DvKWHNXgFAhZFr9gwVvCechpNtVH+Ya
pzQe4leeiv1zYZ1a8/UboNLDWlKQFhzh7J4HLFjK6ip/6oYYu+MA0Nc1afkkcLea
MXMcUnvkE8B1ikuYbQvlthkvxKhGSASlnDBg3tPnHO7a8hRahVRWcCezo+txB5LX
mpzpKDnvXVEf2oSK3frLR6V/XWWAdYHY8ng2wvgmyNdl7QbyJMtVIDBT1R9rAvqK
jNg7QRFq4aCCTcXTRUtAYijmnl0QjFMdJArwZOJ42UrMznWc9oD78WCk4r2+KphC
GUu3nxSmNfiyMnz88Ffj5mGG4pcBpS7Dgh57LSC74MwPE5RvMopTE30c5OpNU0wx
3TpwBHQCspoVaKyIDF10FuObLM19X5dm7+p+wwGsc5DLcQ48Ql+PWlD+b7pnIF3P
9uQw6g8+aFgvJ3S1Y2E5OypSldAmmuWdL8EHSXvO7r9f3nSRDHOGGcbzFds0Ff0f
29Tkbnd1T+xbGj/9oJp99bbmdhIAEUx5l4K+6G4nbySw5W4E8NyD8Tt5YcfHS2RN
o2gX3gKqJjwx/Vjv19MtTsXuWWeBqIMNRdXMUZCX8CvBub18yYgSNtdVhyuelopp
ygNXH87My+V3diiyaWrGfZKoAJ2KMuwrWFRKIMw4xIlEhFfKUFq43nEmUq5zidmP
DHSG33xwyYmdvX66A+9eKsgrEa8yoZp7C/YCU2I6mRLoz27nbvzJ4Hg3WCExKUxA
S4Pgn4rydk6GEunhdFUXwlEIRQeZS/6R5fGe7g3u01Ba/b234Xh5WGXS1KtdPsFo
Fj0sm1o767qv4vVmE5nQBvNJwLQjKbjMbOCuXajzLq0vZvDlD/Lh85+mldG4UnZ+
+vbtqqgGGo+vH7VLnwYc0LZhnvt66xzlzAZ7aT/4EbLtoBcm7kRujaaWYhfeQ4NF
f3wG90nnVrodqMwiQR+jjhIh5u+w/1+lQQki3sRIVNybl4enRHIaQ4ZHG7ptw1dU
FWsLM2BrXNd974lloj96/fbUa690c9r8fZtrBpMgKl/CvpcFcp/hGCHte6T82Qfq
bTWcNB/6AbRCs7GxD7HHt1k3qjiyhxQfw7GVtPrUSw74t6CSMr1isWAmWtSb+X9R
Hw6xZJJ00IYVE8IAadPnNbabOgaJmmHHvcdjQI/TY4Wfa8TFMjPxzN4HrW4cxqbI
JTEqkAJKIG1EZI2MBKbR59YplJj6fsppS4aYk3qZItwKHpkHAMYc4G4hzlY1I3CN
mV2fT0Y19p60HUF4WEJVNbE1sFkIDywmldl4mdkFcZzH2h7NEvO1GlDhIgLbffOh
M+wEWRCLqeflsmst72mO0xC12vf+NBPQ1taiXXjJs1QNL64yXL7m2cFLKok/ViLE
IPJXjyQp7vj52nM0h3S+2JEgLRsOB12RODOI6ka76Y1C7tbzfs0SvjQaztmv0ke6
k7hhzzpYIfUJRopMLD3ZeJGUGEcXJtGvrn9ZP4CNC7RDe8hlUgMBZ8EFzxsF7b46
cBzm1FXlU4JRtyUO0eyh3G9OcjgUjsEgnVVhrDLwA80xcG43A6hZ0SS6anr3kmTO
oDWPKdlMAJODJAxOcSxzFEe9P/2gem3OblLiLlsLkIQqdWootnLX+kK3ql3nez/K
m502gXGsbdg/zQWbDeESaRB6NTL54gROGRmoW0SMO278GrJsL/WIZNFJ9DzOuR5v
KwPMXphs62eYBtYxW37xp3QsufISa76OxEewz89sqc/UNUHMpRyaW1QgYFM7J1wb
3EWWPMgPyJxaPnya0r88si2oZxztSZHrw1s9YS5+uRWY+efNtizwtU0elfS49hi0
ReFXj5dhUvv4kapTKZQPd5qwICMFOoS9CDsBczyn1s3epfisOzVIen3G+wudC3QQ
/7Rznk3qESAvxjlAPM0J5j+Lz2zM/NQUiH9aI4Yd2GSlS4n/KOhqoL+0TRksGN6a
tHYg+ArnBg+Y0C/QFZJb7mu4rxfY5UUOxd+WhL0STBmoKVcnXTt2z4ZbGrKSsFXh
ND+i1IoBjhLxOnEn4Zfw5P+AlIKtSAuCDnaeyAmgBi+vGE7gJnDqnbgH3jjmx0Le
FKxwIgqtxnvRTSTucljGrybfHJvwCqNcBdvIyWKqeZt6Otn5+F4bIWj05MLUHnRI
Znzjp/wQXKhGad9C8eG2Obr6dvIJR43Zuxmq4PC8/YxRv1VedgTpENc+pTLbJgLa
7PhizqMe/69655aV2J4TVTgCUBTjZrWtE1Tb2SVgj1nZCQXcaMjZIvMoUwCG5n/n
3mziW1YwBTZnzh6UiFRxZsXYKPOjSQUGyfgdB3g854nH97FBjXQ57MTKc4Nek1B4
CeLTvM4/R07hNNiukpP9ElpmnDclaOf+kIkJMtI4H/wtFHmkx7eRFF87C/BrxEwc
0hvSbC2SsrAex5RbXXSIoNEMH6HGgXF5Ton/IVwBfk4VQAYBkFWcMV5dCFL5CQRw
MErYBAPhhSCw6FBlx2atNQs7Ko0QenM0ipISo7CmcRsHdp0UvM36kOZXLwm2XXrv
bh/h02uvXp3XWioaoFJX+1WOGml6G4TsHpwkUgs27HKW3nyDCrE07t403klwOUT3
rxGwGThcS6Nvvhk/vkTf67j9HpEqCpt7R3tD2Pt1VXXON7QOh4lYk8hS4aJC7SEQ
YsmPJvstF6QXJw2B3DmDW0tmUVKzA14/pXjE36QkA3HqSYUFQJMCHcAHbwpzaf+p
Jqk0zCkJew0WLxLWQbCjO9b2jQkJeU9R7QvVxYPXNvJL4xzUVhYIOYyaffpipQwn
XDan7D0DRT5PLaOzBj2ZpuxT6BViPLrr4LBId41fbmZ98gmb3Srt8oQdSSs4Jphv
oykkYTdEwGlbfHXgNkN/g0sixa09LNz97HsYg2ij6Zfb6+xpLyTQ10yble3yE10Q
DUu/OmE49bnyGICvQlzyE3zMo0zVxtmlT2kVONho2RrC40FKA6q+eSRq2rm3yXVy
ZCret7k9VWvpqFh2pJkn/EklHJ70uVLcd9J5EEgr+LipGIak3j6nyst2jz7Es2Hk
Jfw5DlOCGKMWN80ll/kZJYPxiy87H56ur83mc1gMj46SziDIrrRomy2WFiJJg5k0
OQ++iFqOtyS59cw4Evqu8GFyoQl557cy/uWKbUB3cUG1H0E7XSA0wAo8xRwWa+zG
l0fddmMF8IGmKh5jcUTayFoacdd5eTDlpB/7y6+pPTd75iw73kIn1iFCHYpkSWXM
fE+WXRph0W0ifiIiieW9DFrQWNrQOb1TDxTfecHS40RpKD+HngwZF+C13YnMqz7n
hOh7SR9ZcNj9JPiOEl1lIt/XbO6Jz0TPWt4rUBkA4F14hxzW4MFrLFxNymHbPUWa
ZcUGpcfd92GtOKd3VY+o3J9V0v21VGD0+pgDn3rJXK72TYLjInoITP+U7ByMjIkE
tsmMW7qkrEohgk899OY28nb3bHcyKcIqwi3NpY680rstHWzSbKmRW4FXhbM17e80
4iDlkft8hkAWTamA9ogE3v7yxlso+jlqj9I694hxzGrknZR0s7+udQnnDs4VINFG
JlvVrsIM3wa6eiFicJFOg4lNL7RvX5lcvSS1vIT24UOMDFbokIXEfqPa/bpWqOSs
GEY2FXuHpOIqydsoMKOC5fKgZwRICgIbcjhPYAqswcz4ewL+pITeuSQo4X1IXLxi
8si6of9pJHLzaX8vCLYBKnRf1jgUMvC71kAHX5rC8SXiyr5K2xaEpZkNmlH1VmPw
YEjU9IGSU23ogXK5eHw6NWBu4KxqQz70XkAc5TxQZdIumMoYUVwbT2GYo9vwkYVa
INkfZ6hPDfIV8UBAQ/GZudHdsb/9MszIW6rzkAM28cbbj22NrHNERgpxpxUQ1ZRq
7huP1eEZjqtzNwbg0/Wmb2b7et55MitZ6RXemGpoMPemPvdeMjsP7v/UQllEEz28
MViidlBxljW2KhU6qne6k8oc3BtocvogVzCmEKzzastaXzJgFc5Ckl6RFN/giSFc
1hP7m88skfuPUqI1S3LjuDSmlLFN6IWggCx1j6Ajq4mwIqIz3L+Hx5prV8eHLr8z
k9yYkCRnKClbwUnPxRFZZMyrIiHHS17stCWzhbZwoAKQMstosfzppuqyOf+4Z2fQ
+W6a5IQWaAW7LlNalfWOa+kLtiIsQBh8SNAvmOWl6YkKYAwWUgr12MUYDkjz63Yl
KcsNYdRumkcKgkSivVCDnGZO+8zb2CI/CT6ZK38rxIHR9Z1vgIhOU5apcwzpaQZL
BYyyquNs+gQ9V+0w83Ze25g+M5mc9LmCg5P2P3e/rASyR418tPPDgVoDtPxxnYRQ
1vw3j/yqLRdOCzYT5HzQ9L3ZsAPvzHCF/oG6m7bndk1zribjIInMHaBQpWsfZJCH
AK2K6uOSJRRth+b3dEqn3n17K6ToqkapXW8xMiGPKbCsVS0kcn67aAclfBA3mmr+
02bLJUCDkCEtoRtq/U+W59Wvgxmnozjj8VXB/GtEhG+gFm2bTHjwBasmNIdj8zgf
wIcWWNB3TnqWr4jrVRZ5HIe7ldd0nIcAfhoQPxYNO7lG93JHL+nhKaRMgYn5AyIF
hgidqvJ0UCGDkg17VkNpmgqWur6PiV/1wqn4CDFHmxFsy36SpKwnte41tfj6PhJe
gaO4N5yFsMb/w5hzY+j7a9YdY6anbOmlf4WrIlZmxyMO1Ruq7DK21DeJrZtvGZac
m4LPmMH73XD7fh7tbVvEDY95vNVY17BkHufheBlRwfeQGdU84gEqIxzTRKH0+Oxy
07YwN0A5FCOFpdx/aE1PNXXZfgvgFksK9lLrqNqATkqDl8xDaTcjNFzm5vCMo5ea
66mobjQokUh7i1EcDG5BqZDt3gEkBfVltDZsIWQPXkNf+9c+32IWq05j4ESG+DYp
jLxjErUa5irAeFh2L+amH4VKryQBhq6gBBx1EUwQ44Fa9rwvmXFGqMwRmN+2rcN2
6OfKuZqlbKrd+6kILmzs4iLv0H60JXlJTBUi9jZv97K094O5DLjdgXnZ+rTdKpgp
C3/tdzVvIah5ywdL77/eBKEdc0JbUEqd1ghqZ57axvfSYnuX6r7WWmXcY5Z+fFmA
90hgicUb6qmUiruga0CjV3jGNS9tBeG2M2DOW09IaCsLhaI+3Zk3wZk7WhM51hdk
pl4V4PfE/jeZ1AjJT4vZKyrGTrPSoYElutsQ6KeMSjhjNgaTG7Pw2jbnXgSrbXVd
1gVuMuB2uiVp+TEL6BfjJIOIS2D+B1+ICFeUWo5BQRLf9HBrHD2nxi0NQP3oJwns
hKWnKCEPPsWG/cTMKfcZ5uDef8AyIf+qjayM1XocKqQKvSdWvxmLiwz/TrBwFKh3
R6YFeaalh6WR07BbRS5P2ctSihxb4lUg9UHne7T57+pcpW4j4C37I73Ajj13B6jN
UT8kWAFJ0NtnQXBQbaW4RAoPSVf5RB9zDtIAn4dlvDr56rr/lnRRLCLANWu4686Q
w/VvJ5rILjELgQlW6H4qBCm1w0bzhCSIgNtjpZKPva+/SYuKD0GNArF7/WFiNVmE
b4NJyrod3yAhbG+nREHH0VYgJGfEIWQjnlP+jxVjiD1SqQioNgoQFCPwdJ4CTq1y
v4LngVgFlKUr+j8pjC7H3OIxscv7nfwg9ySBKL9uakXw2w4SWThwJFl2th5OiAue
0QnmPBhG907YPkrBv+VNpeslfkDVSFqSATPfuDFULO1mpaizTx9ElPuq4XtQliGA
KsEL+8Xfmaov1UV+JFyziTFypGj8D3CpkEz0c5/0L1P4yPaFz8hOBf6EWxbKe+be
k1b29VatdRInrJEsZ0Ppgu/SsARy08CN8fshXqTdj2V5yyBSygKvuD4PGHSeg361
xYnmt/sqUMIzF8jDDDQJZAWpptpisq7EgNYKhQ7tKKfpMcS+2qP/0d5s97+4pGPX
fi6MK21+szsqd2ihf1KnciiqxK0WDx1HGB0GLKLhoe9yf3Cr2c+8d1Sp5S8iSRbI
xzPblXIogp4GOMYlWZGmUzq7rXPDTDeHbRxdquATCi2XRik/AdmZOUIG3ssnJD4h
9rqyjp0PLDKDdbk981qjmoT1CYFGqsFFXDiK2ccKGp3hUEtN3bILVeHjQJn3kOJr
x65jEWOmYAgkdTRsz/rGB9mDfBBIV1Hn6QyimZrKHSZfAmOVQHgwfiBId9eLr5Nn
lk611aJgDO5cmoFaqW5I8f162eeQ/k08y/ekF3hoMFH1g6IQQiUWopJo6nPJSJNr
tRaqD4Lg5lgwxshulur1aE1rSLR5+RBrvTtKi9FyiDCX4A6gAHJBGX6t+RFqszqs
ttCL+escYVS/lhtfHwyxe3Kvn3jekrNtmk22O27LA6wBxfpRgX3cvyzqjp0sLV6v
FsYSVWybQEV1beOc51ZnnUSUvN42SFq3RIeUUx0olL3ad6CQDaPD9n7fah4NxbgE
ykyn8ni8h1fSAWpWe7bUYEuCJz7EEOVff2rdcvh2xd+AMiVz3mGInst7HRRS2NdS
AmG2C6LJQmhw1lLB+ZEXGdDIqpzkjU1idR0xaJViC18v8eptjr75hY2v0I2ZSG6h
iL9sP30eh5OwejlYSK+eU3eXYo4l4wOtxxhFPP2MTkULJIHwKhJrEeGjwoq68t2Q
X4l75+NK3eKMgiXTosw4YqVt4uzGNwpT4bcO82hODlaOxGpJOWOz/VMoUxyGLMkd
9kI8e/YicI8sZJrOGWFDJB4kELoP/rqlvPsnHp4otZP4LOWglp6ylUV2rjV9hXSR
wpbNj57E7WXsisBDwdLVZteT+eLBuLJRyN7Bx8EH2EJ0lLW0j0REf51UGSeJfADa
4LUALJT6yBu+q0iYkzTPE/x3gGBLVXCNb77RWMN3MLf1AYn6MScsHvYXp74RIoEw
K9AWvNK5UaL7UaNJ3/8V0axjyQon9MJOYhf05bBZ+xoCbIwEzloqaAg8bbFnp9UB
GUIqW1CXIqy1oGtHhvJKSRWuJM1H7RNHcXUGX+hlX3jEJXngqHGjHjLEsExQHDAZ
aNNDlK5UyS8YfW9pjmFWrjsstN2Zvd8N/OoRCM68Om8fZCu3huH2kgMn29sSDrsB
0U5PA6E3+XvYuS+JBU7+c4wtUdnlXXTL7Sp6NTNOi0Wgl2rK3ed3f0KWeFF4eEs7
d1pEyN8neupQDyMdmuqoHYYm5y50n1pAEehGBGj05e8VE/ZbZrH91wvN4efEndUT
oJY7c/Z05NeKElLpAkMFLucmKR8RZ0swn7TqmBXvl9rNt02oRHFYY6nez1DoGygF
gYnS0ujfK5vkGSpdVX0/9JLke6XjdFEknKyUSjoQ/6CqwIPj8tOSXpQBXYH+neUH
f+w4EjcHE0JxyimcCD/D1+6cYuRM2HRph9qmP1pb5u18TxFhH+03tiAerUnqLsR2
U1UF2+g7/9mHGm+xddxf87gqp07IbCeakknDCCr7lVUofOSV8d/RCGOKE6Zf+0Q4
U8nZVxlNg4D2pCU7VKruixEKAzbRfMJ03GKPlQ2epY1RwKc6jyU5yYxsQUHW2AEH
5/u3vstyfRSSFtEsbeYY6pUbv3XnU7ztGQNWAuEt6YIXzTE4Uhm5tWQdYuAiGqeN
b42MQltZL/K3rb5o/hSc2OtcxvjhYSIt0VT/FHz2bRjQ5FO4h6Yx7jLRt00Whzld
VSxElyXh0Pr83AZceVLRNpbzbdzQI/JjTG1w5EMoRedSD+rmUMJMbon337CYKhVd
rTDHN8jVgNBMF0nQpuYVXzxMR/4ZbQlQYyRedT5a6BG061no2zEP0uUfzm6+n2mH
qDLxKPTN7e82mOdSnetwPnU8fVpjOABb0jlX1MlUSOFJZc8NQoTz9ByXfW16I3T1
ZX6V5rG7lxbpxlUc2nT5Ua1wO893nlp9tZBdezMJEi1a7bKl32OeZWzRUmcHtBS9
nPQ1KRRvv/GpitFbGjGNsu6CCKPxxwgFgHQm7VE522XkycYaTcK7jNf4kukSK/G+
H+D3Zkg653xulSj0KbwOCFde9KQqxl/zBFJIh7ab4+1vaSYkISA9azKkhpv8Sg63
HcYBggt3hJtigtx5xWDfQHcaOu6PAPV9s5zSCK/tcqp232PAowFa++nX1CrBp3xc
1fM2A5M7dcBx5g73a5NnySUkoykgGJ1JmYTnBAtE07rc5JfTpt1HyHmVVoUNU7fr
SKZGtUpoCDYurXFSrN+T09rWYc5FIqYEp+eJQ+FP1uJ6fnlLAe8mTL5i2q/e48PL
01WVOgn+jj520cIsyXToEqPkWcMJ7VQkFOhcDvcsqWbJ9QDQL3uFhDGxydG8tGQ0
G1bqSkEgfp7a0t27PkdTxakaaxz4YoR7FkjIMskDBpmtrmm32onQC+i5uPsNEUtt
yaGSlL6Ht0LAXrWVgtnX2nA4xneaf613TOuSN4n3uxnkZo9Xg00dE0guMApmkwY6
WUpRoq4KZxD3e4wKAtUh0O0ldbwGrUYkj0+0TPTa4mWSiZMFB4cpynTBfKadnYPM
hgIP8hqLZL7IlySQJlSi6WUADtIhKCq+TjltmcoYfjyHgnsTghPNxs5mkWxBavhd
pcuaArXo3ei2HHW4w7baBOblUOgx09EzWc6Sgk7mh7/W1bxAzMxUPeq0DyVexaaM
aS0uqUCqOpHNoeRqWqp7mi5kucTYOj43LPbMptcvtXFlhZARPt/F5AXL9s/5vDU4
1lMkiQo5CpyhDhu98s4CYvCBW6T6WL8wK4Fe7DkreIDQpNcnM+pnYshzr8t2ZDxk
NdRBuSxwwScX1Act0dWOTsLXru0ZHyOxfUHLODbhs0lq/9YGr8QGFr3DR0trKR82
82bF7ok5uRxpGyY26WsY/C0JC6sIznbtH8iXdSbOPtCTLs8d89UcsVL2Jy+0k8ww
OsAzvRROz9vfaIhGZ8w8duYIg+tSS5o0M/3X0qBidHK0mXCOQuS3p2TDoPBHa3Ag
9GtFQatsZjqMsZB67iLWjWrmb5go4Hk0K/w9gNlNiZECKtgrZmea7z00iW+kje/k
b/i+kjyxMGi+CmDCaws30X8MiF7Vii6QH6iDKxQN0wrq74pUmZw991WVOf/3X8Zp
wNN8WJ2FlTprWsX/ieO67Gb2ljcDpqXlpN6ECYIWJOF1IqWLND3n1Y0FbePH1qmO
te/7cnAN+vHgiesD7cM8ppA0xS1bE//9qwgibjDl+6NVlx+HQNBmR1levGG6M82b
C3aZEXLVNkAx18dIiwknq0jqPujyQhxyZ1SIoJ18zQHHm40Evs7jv9PuCmGN1HfF
ZA1pNjXFUcMhD/QicXqJU4M0ya2HUYgqMcirm4oNDrUbHPU1UTAr+UiTfl5Dat5X
oQ7buLOqoqQI/o1903QzNVfCAFEHpW2reijT9Su30x3dVSGXtz9I9eN137/J6WcR
MLNIj0rfH1/dsrUFxYTTq0byUjWqkZe5zzG8ozjopJDAZ2rF/aLG6KVcLooOLUIr
ieCXjY7344MHuiSQ5acVrvQiFn3QRyKtA2iTU/l8mivI74np4zT4vTwWzMzwW0Tw
HVGfK2F1M34qt9ZKDwgE6Kaw9j/IouCMGmpNkc0Dhb2bJX49iTtj2nayUmUu0XeM
yA83NVh9++vAFLm5XZNvQbEgipuk32tWs/n9swHZKYY+bbOI7j3tAo/oPybdIOla
RgO/S4b0qr7iUHQyozYss+1J/nzTJPAv0nE9mSFM1Q6mf++LRSn5WqRF4zgq9nME
8v2p4UIw8rx9S5f/5WLWds6Bl0DrkMsJ0t7mkzeZdBblYFJrdsz5iwN+EISjONqP
2GDnkVLdPRbpv8//wjz7524xhxS22/cDsyBZ4m6lShQ+SAKvC/lxq6nUwSqtt8jK
wOoQGFeG/IF7f5YuZKU6915LO+KZRlqFVMrlYdDmDIRi0Dtv8goYLrH/p/YCOQOW
9yoS597lxGSSb+0bNr6KGouYG138FN3WNamJDa3uFd/VGuoLecfzoVjfbXoq1JQO
jAqVlel3hWTYlUmrfSnZoGx8L8MyVYbWoAzssn2nHZ2o/1kb188beiRyHFhMC+xd
Mta9aniOUA41no4kzrTB8JH9mus7CgJgoH2p1brwu54DlpdmBhxziyVvZwa17Vol
ej/0KQqI5sUGfLtbf77+qiQQ0bpPsDdQGd+WIkzzDEsnEhzRNqYzFdRazrxBFIrn
NaUkY/kpH/DwaiEtne09J37DK52WZfFALPhD7bPWzPdBtQYCh2iG9fJxRkNwGjry
zkCg9nMRdIGXDL6mDaZ5+86YBgSBr7lunTSWgTJPqtLeVTGSl+rSd5pPOaOiUInd
3oJykLNCt+oVgyRrsbSK4ErKFs/JZWDMcAUydMGXueJLCTM/hMdSGeJJeP5kqUFb
zF2UvZ1zY3h+pXgl/I6vZ1pq5xLG3hZxNTFFaNdH25pfDZuQk16CMzhh1O9ZOG3c
g4K5c1Gk4W9bBdYotoGu98t9xfCVAaFH6eVTLNRIARbybp4R+3QnID0//vLPPtPj
TPlv/xwY08VSe89qaU6bsjl8P4WoY23vKHw41nrlQHl3hkFQIpcqNjgbTBlohzIP
9Eki7W5z8ERgtbpH8ufR2h6H/2Db/h86xbTveKjSQGjDiCDtno8+dNQim3EenHFy
wziRaYT2SGeDWyXEievme6sKQzzDBHu1xIiwLoETeZAijRU7xCDDeK3fIkm/Jl3m
48u5QVwfyNZplbirPMFMK7HYXVgTD3mOIlPLDiSDxy6ge/7TFzn3IK+JSORBS1LU
zKx2g7pKm7484xmqCuoKUa+W0Fj72FFjQ7sEQb/RoEquMRSATUyR2dDpzghq0clv
ypRLsS+IbwmcAMSyvw36QqyeXSshrUwedUYn7+KPaVgwioI+P0TjMyP+rRtbwuf6
6Q1mfqRiDvpMYjYBEZTvTj3299buv4E3I+Cen6l1z44/Vq4RIGPkBOYWtXAG3Dq/
HUOfHU2jgIkBfV7xI3uGr04WVFTXKxBZWN6o46PSzhRvrepP0mGKy0ye+9lWmPUf
AZmwa7WPyhbjCYGAkol5f4UwLWCeWS7B2xaCnv/S8WCLYpxfTokoJuZd4lbYimGW
iaOldNeEWEH3sN7tB7mRcJGhJWaxuzkbRCunv+MH2LKEqm69mWOF4QWIb+bqyBnm
kbVQ7YAUSWh4G9bHIxjn01gmrgmIN6CFISGTf7A7GzTxQd7KR2ligczX0GY/YG7d
9Kx7xci6LaWFF9IoinpQFH1TeeabhsFx/TkmSN3q7toxCZwRQly5+mV2Q6Nm1wHt
JKLpgLBlM1PWaRZlQjsEORFTMJxTCLoJV2XUcif2qEaXxIfbT+2q76JdsfReHAJQ
6zj0Hz1m6Jl7q7sHvJrnbatze6AX1Kb3VofMYByXV2Mz0gYL1q4g1vFexz6Ezcl6
PTkHnvAi0O802wt2O32eMNPfp5RemL14af6aCgNW+QE8cuLzJPvWFwyDjVhX/eP8
PmwNu/Mz8V/SQFzMhLBLuLlKhVyPwt+iCMuyKbeS5qDA+Do03vleDOicnhDEvCF7
sEhNNMQO/zU4JUumsm9KuZUm2AI+d6LYjnsCpmc35rEAJ13zyvquBIzQTBojLAHv
1IQESK4QPA4a3im1e5k77EXM5V00oVYiP85BjpTA2UT6jMgjsYSOcSZhgLjekENB
UJ3Q0ZuZpUMoqJcGVKS0lWw0f6rqFP78EegCsWnAngGd91CAyvKPkfLosHkiDO0l
6B9As5aG4wV61cQjey0KQvCNP/PpEG0Egxg6w9rM283r5Xmmc0WHv7333/+Jm11P
eUMFGqKBP7AvvL3aLpo/QpMJ0X+409SQPqzzvryCBmiqOFBDlQqUCNrHYfkI4ezt
NaojYgiXxDiJ5IjwR2lNcfybW01A+BqKW4suI0Abx2Dp4XpTpkB2AqlIdD350YEZ
ZxwuPdbmoVynzFP9rKoergw+Hv64F/JQzNv4SxbmoOoQCopUCqAl55Z1Nn0igvGm
nIBR7qzf1sPeF6CRrSWXYAAlOvGFJ/yGHHnQjM0qnvKPVPOwu2ZKBJoIhBrbWoOe
jaqgWKJliEAfobH+nzcJKXoCOWCu/QGJraJIRGdBicam/U5ab8k3ClDms/uPUmHF
rQslpvI5e/r8yv3lnEtsHvgCRdkmyAZf64IshUPfoXclZJpehByPko2CrTp4F+Xx
SXcfki1waaq7jAOggVpNQ0ISbTWarJNVWoZIGO86rhZ715yC0KTrwmZkuFI+ANGC
7FsxtWWBb7m67PRfHOZvT87CJR8qAomSR44AnHuaLW+AOmv5QYNxhHgFeohp/gpl
kzDT03VXCHgUiXI1nBT2sbAO4nN5VnQxxMaBO4D0zoM/rHNytVIxW+HnL5n5sESm
RrM8Hfj4myECQXhoGpeL5t8meH8ogP8g+jpo9+u2kzR2/Pr4bGqutrlqGfWFDw4E
C9TycNcsjGKSgnuiMKOUujmpeRJIOWXlmXECHavsCbraE5iHzS2xMaHxvjKsRQFZ
qjXNjM5CJDjqBkhBF/YOoTioYKzACvcvaZtjqBzoEKEhm6ZT4enokvs+cHeneaNW
vNe1f64n5wLOZhYhRlwjD9xmEYelEWd82tfXDFC+5m/xFkvKwMsGeSNBgpCIhNHL
5bhqTnKK2LL+cMG8+Ip3eg/wD7L4Wela8PLl8Fma7/ahG9qfE3S32anYNP8R1cM9
9WDgODv7UmU1wX8wb+W6ZFePljLfLj5lYM+s3lHVLL/dL9ytplR3v581g6z6x3Lm
GIm+aufKVD7AwZqXERJUbfCeniRbXc8fze7jkbC2pqDaTSJLWj0vo9f0Za8geyuo
xdJ0Tmc17qGAzCgBZEE3WwEu4cxMLix1Z7mlj5vgoDxuYSv14ukRHzAksOeRjVXe
Kzrj2vzqxOoAR61jexozflvYHsZQi+RGBtoQBMOenVSgdaNsDItow+37yTY/6Pcz
O93pL7Fe8OJ0HrTvPmHRlUikDUpCjdlixBXWBPgrNyO0a+t8a116NoOt5G5WF1RU
9SADaovz9cNBiZqEIRNCl4LkbakkJh8lcWQ6eIy859/SnAF8dDuLq8D0NBPqY8aZ
nns4SV253aZMvWgDebcUg61IPavISjXkAN8r4I4zpukopGVlX9hS1Q3NlrqsnzUB
LTWo35cDV3BHjh4CDRuQwblb/1lffurPOdy8mkxwlBxtL8MnTjmn3YZ25FX4BB9h
fjO4ReqzIpQX8Br7mWOZSa+77hI1qmPD96eSqEY2hkcq8NRHEtEhdj1vA73w6J35
KgwJfU3Yf92lbUwav+iup/oULpRLItPrilb5iO/+BbEfRIg0wJl3BGtWdScRwB4+
22bWjer2A6Dtn6EQjeRDnP+WvSfrjkYTF8t+q2AFFrQkZB4bZ5FO2c1wNW7qNIEj
6u5C3+zwJS8xjtm/5TQi6+maSTe4lntXizUfnza6dNAJ01PEwXIuTO41MS6ITs10
4/N3mPkdCbauuSAruFihBnENqVeDZFqGsMfhXbAC11uEU6Fo1ff9TpKhRfW8mcV4
uCKoI9vd8oOedyTHBtSk47yAFygjK2Rc8kEQP5fZjpOU1cBFiW1ipwIku1L2+sAD
/s7kGIwxbY7J45ClCfRHuCQaFaoA6JXigmPG/jscUljNYcvvQn25kIejk7+urR/S
d+9vk2fhs1CUnAsrnrxXmMVkEZ32lMtcIVhAM2brE4CN2CAm55CGj2LWBeCPBdPe
ToTmhcf3OYLPHMG93zg2bXDDfZbr82driL5CJvjWZRrYAGdAquRj27m/KMa23NEN
3sBjzn+vixHMnhVs7/ep0rpcEseELKBimngUONBI3ApBNzg357mjmOScR9LNyDkp
rk7AcyCaz6epS5rbJkJxl5TnZLeOQ24MdMlgRYnj1rFNmiH7VAHyEbMC9L7Ftv2M
L4Wq1d/p3gmwFXw/LXFzBF8l2LPMBNmDBouRnm97lYQaf9LRw/9/YtygKuw25fd/
YINa3ixTLq3V4Xkn/ts1Vg6MVSEzKdnVnssK5yQJK9ijKAq4nhnJuH5bTAzlfgFL
91muHhcRINibGR/Pw9LZcDpPeJL2T0g4dj3/4N9pjfr2zfbxZHe3fgd0BFr4Tdio
tZ9xILM24NIiwq1AuJzL6GdIOShMLzlwtUWNKZAFmXX+HiSDahv8wV9+i4uPbI3c
cFK7U8MWHTpGMSq3lgZUnjRAxSr6cOStMLNeEMlQRSBiZRkIDFdfFyyT2jVmhQfH
vhZoxoo0BYtQtNzXn9X4fuDrHpT4KS0Wckxy8fK1SRwtKoMQ7ISLLapzO7xESdOH
jQHSXocPBVQ+5FK/n31rEVZ934d8O1N7XtyluZNSsniKgjvAQm5dL3ZWo/+wCV3n
pIuSOe/Pj5oXjo+rVofpmkV06rCkJv/Xg1Umk4AIKW74+ziMfIfX4US6rxO2UpPP
und7qbmpyRXHi2dChn4bcT1qCUj5d/kjN8GiQqzED9QHY8jtnWmyGfNbHZya7ix/
sI8ppsRD9+LOjnOFP+SDuuJO5kv9gx+Fla66ZM5mMi0Aj1BihVtDjsiLXuXFIrQl
eEm71HL01yZrm+MjdHDIzNSSWh4vHoNDrcrqYVfuTULJBIoxhKzYDXphwLDtC0ir
Ve7Sr6Jvvz1WMBgmHrKbCFkVa9jUANQF6LFayTUYDao5+aWtJqRT26uiVTM3/gKT
q0437Y9yItnM2FkqreuSFH+rIfIP8uenKKOFajUHEfCpdBeau6yLeuZJFc50ucr6
kSjqWgEf1JQR3wxTxghmE2RWlAtsfqCj5yhOTvNG1HanXHDdHGXCMLc8mlUYcs6w
oqqafzydjL5ib6VHQhWlppGX5Jyj+2vYRha8pk1uU1Jb8xZFY/3MsouYTeukuSb4
Cl9Slq4fAfq7H4s4n//GM60hKlhlvSq9eU4Opj/rRzMFebsf6woLyZWuGqS0QPrS
npF7f6xV2rI+EASZV4qfJCoBifwnNhzoaNMuUBGqbV86gOoAEVYeySahtMfDsKpn
ji28Z6Br9CefaaXTVSqX6T/XBIDIsitW8i6pkrGrCZijlXJLMMU8O/H8nZSiUz4r
V83yi6E+5EPY0+KyVv0wdD3FGl6tsWm6s1ALEqvYdPEMZwvyO1l4EsU684TNKhXs
gqdNgPBFbuG9L1qWVhr/QUshGriK+QpZykPXciF5AHldqmQr1XKKY1SuaUh2gyK4
QFuypWHrTQwDxNtSJA2WGhiquitmksb32dLwfFmkcKluJR1mpF/4nt3b1LGKuBy5
1ZoXJpqH5VMB4lZVO6UIC7qINyPXrxoZoVtzKw2KtMfie8lJWJhojYlFOAmxglTW
flu/ZszdqDPxTBDAeYnf5hFy3UbJ4d/l8z7Ij79jz+VsCzFQDeqqJeu6CmEYBzEA
uy+b0lly7jkG9xO/usDbRbJMFl3BDxV8T7XW2GlqKkVxZ7tnzXidSSlIMQs8wO+F
CrgOdZJDwr10WGXVt6rd13Ff5zPHyaCZ2npIS+Xdt57DS+W9MqXoxdrmSOpWooUn
8Cg3WppG2By5C+u3tgVMHB4kNnRRu+wpYK1k32WycoLEUrCKZW4hN+0OKH+G518C
SIenqqNgAy2bS1mkQDOxJBxO355q+igm5o8BbW64dVVwaWMeME6YovuTgLE7tJOM
N1wMNzblePF6jVNy+0wZ5ISho7iuf+sirisXi/mMtQraO2Eqed3HCTZl92ue54DB
v8YY4WZ3bspYxm/9TxY1C+BAuopTUlyZYAVSkv93mkAk90kwhsB+kpwwfvjqv+Lz
qKH48m1dyGfqW3vTQKMIv/BEtgdXXuirf4QBYCdCszFsflUn9Ad0UrFgMivl60+D
zyJJ2AxV0EVwgO89zlu5es4i6gVG8xE9TWAK0L645bjqYj1jzlmJjxtytciBX9e4
8bgp7sE3hEGgM6ZIGQDnxiLS/Hliei08o4hn+VvtoqrbK9WiBtJzDug+GqHSw/AY
ug6K38Pncxqn/eun2PMSSDNGWbTEzdLneS2jxnAF8BqPsPflpSz1flIe4WiMDZLB
SGIMo7PF/GWSp1XbKzSDYXxncSDHSnvZDktNMjsM1CnbAvZtzf6X6iJ6DhPj252Q
ozbA0xWrt0+voUhKgm2Q0lXRWbCmb3AcYqCIyaXlCy7+vuZsBZRBILB+jPZ2zB+Q
sQs8TrM7/z4KBs7lTuNCgpb9IeCvOTMHtMSgH7Hlh0/5dhfllcRYgJZhwRK0B6vp
Cqi4BvL9GDgwHGQF6Md1txDcQ8wEoZcBMeI/Rn+9EpKIuzJiVcf/uQnVPk6i/uag
O8mjffi2g0z4sNyhodOnn7oTftQGOljWb4V8DeOrTXK2grMTIv/dzO2XwfI2ejcd
Yey3o9lvpeud5a9dFJI2X+fzBDIXcuaVE01wu+ciflpdkx4y/UUtXhTnwCBo+Eli
HasHS8o25GIUBz0gOQaz/8SCv60EeOHXw+/rJjSTnfNAszjUPPP90fJkGq4gSj4U
K1mgzY+VhTcpGQvFxcPd5kIXo9vpu7yPHtcs2ZLPKDBXnU9H6P1vnfCYaONqxCOt
MiQ8uf4QnumbBnY/v5T50blmnU7qEOVNS5AQCKguQZRKHR8mn5+GBfjchRKBkBfv
GZZEV1D9cbi5/h9gNVrcQYtXUTp3EKT5RIVs6QpgZvtVobliSvPvu28J/wStmEWC
z0ZqlkLvYfqgV6RB5WPuNeept1CSB5DveQpqirwDuUvOUzxKpy1GM33XzfMt0dof
wCuVGKUeg/yRbZ8u7pV0TTccfwcogKFq7TpqVYonJecQAUj+LLUDgoiTRzVfwYgv
dh5ebMTw0L8OqyXjpOnAi4ZoQK5V57Ze4lMuk9kaNi2V/3Xzu8hZKFesup9uiSz+
bSoSzPNZkzwC+GoyqoVD/xr/3yzFBBVsUHGC1KRYhZgN0x4M2sKOYnT3g9p14D53
rPB3dm8hMY1os79IfwgijuYQb87+AJsxNzYFTFSjN/kjxarg/IWA7FIW2nS0hQGF
+rLbs9nNeYwgFYCcYNqtjcLh3zI7lgidj+V7eJJN1SLYQJqSTmjg/J/GmLt0Rnhx
AiaSzf3vu0BWGM2HXDT98+iOmoNRnp+ALrKXcNpTJEQrdILQqdYFpdpqKcosy/Ky
cCKWGxJKY8aLMRRE0t8p6IyZ0OoXhLbTLa2OwukiXo9ymbC/LXxpgneiCHOJZj4J
SgHGH22hw36dD/WG9eZ9XWv1oaQSqlJDbNiaW83hVz3XXazLWkcUYcZB91MCW5L5
EYy55TsZWA8GpONbwJJoNPnUoH1Q3lMjaeEll1sTHPHiaT47Fooz0AMOQqaLtYSc
TY1o4XtWiNEXjlvdvjKH/kA11hjOQoEBvPrOA32FwA83gjhAEoR6FbYATdxiCgRJ
6QSQI/mqqjudjoscwpM/QQYiPG0g4vWg9rQRyzojwsMhFpt1DQSZbngVTyZvsH/L
sqEzaQTLM9FLZvz6h6zPvj9ZkJVK1QsXun7U/97ZjZB4AZRNEUQHOB4R9iLgEQUg
yqCdxb084QBBZZGx5yWO4aGyhtCTjq0zFwMiMLX+FN6nJ2bUb4PSYjVAEv2yxGcp
MsAlUzTQ+667fOKzDWj+HZvv41JjJmFQ/9UFt9QXLrgRNSL/pALa+JtXsn+YFT15
NwmHNOed6REZNUmqtE2hzpQ5gxQwfDmAqLuALZctMr8c7iojZ30dlu2ct5W/vUB5
mhwz+cgzHGm+uph88rLvB7f6pExyPIH6/Zeov8x85OB/mdZkfmVby2yt6+7uNV5T
tBzJD/0kzS72ZswZg/ZiFmQNIvD3CE2WU2q6Rk5Z0GIdAUcvJU8O88A0BfokwNbn
X+PlrLLBjHc9+Y0nTkx7mV61CNpr1w825HlzQYM5LU0vEBTPSv9db9PhM1lW0t6w
wgVZZYiGZWJClrd6bx9NEHh1tCVqMCH8ghGzevhtpb1TQPRbud6208skeZ6n+NUd
ajVmq4uUWYJXpUf5dN9k2WOHCV3/ban/o68dvYD4bw/bfHhEYCiP02NZra/00U1C
K+EztrRPRhWvPZprdR4JodNADFh6KhE8nmkZjaxEjsXhFTFo5vG+ixdGY+13pdw8
CK1weeZcSUJNq9eFhzl+BoayUph5oL61w9x3FjMeAOO8kgEUCYcNHaHJwgdnn2kb
nKOjBy/z7AjVT9wLSjsKnBXWe4EX+VktLPX8GiU++sxd86bX+eXbaLpcwSR4xStM
f2nkP5AK1eGs917UcyfJH0wxLd2tzZV+jHayVPzWRl4kDazb5Rt9NK8VyL19mLnx
boXaULlHJbvklAvjc1+YfwnAWmyqJeIw1osmsz6d7ZXQOlv4g4BKXa6de5uOOyN4
IFMUMwGnPJet6bQPwHcuKHD7XMnt79/EI2FozNSwMnRfaSJ0tVdQUk+mdjjWnFSj
kTx0BOLoE66DikNSvafKv1uhrDuer0M5KNoQSKnpSFhLRXCDCPsGnfkhAHxS/7+g
seSro0MtWeU+yJBhZj3ppbuMe26mhKCil+6UIcesRtLdFrpd5bVjDME1jFKAQfiC
5qgJ3lvyYkuWEL9MhIuUC7VVDyqqyOUT0cZEiUkVWVQ3DJhFUoFhld09fM7nuRtW
EDp2HHfKsav4zAYwl7pAYgZsIoRiwaJanIo7V4JIkrgbmoPI6oj+WMVm1NQFxTsZ
Oyi5kwek2oNPb3ufn5j5xCFA7zWvmekJVK50QmgUC5pzBVvH1AUiFVeB7IwppXhy
RqMQ11bsG6mA9HdKnuFBNEPNQ3JG4gkbBFvjcmoiUAuwtrp0sBeAnGIuOQ2EapVy
8WfdscM0LmLJN9oZJludNEi1QAYzyahCyJqduzYgVGOYqJ9SPMTGPe3Y+ilyHnoh
RonW54wECGJExzcDd39qbId+5Nk4e+s8qs0bhPsGMRsBHaiLo+1xc/cqZV42quyG
RQENLXai7t9Q2c19CUuAaX50ZhHGiuybJsacZSS7xeX62ltlc8mYCJYWBv2Crxe7
c69QnJLLJwr8V3bLYXkY3UBgO4jJUFSQcEzal3+/CZ5CF+xctvinJ/InmR1U1qsp
5H3Dk5JBESSJ+fLuABCg7IwYg+Hju01jYean87iwIwIkb3YLpxtvZbItSR/FA9YW
lNuY+Zcbyf4VApVJriym/CUQ0G0grMey8Sjal0wo79kW1YKaxmI7HOnvXbDvjjwv
ceVqkMMW6OmtwCt1mhd7QdSE9ZrE6rviCOeKjujS9Toq5zNJGqujJSCJB6l840gb
IXA394POpS1NKcyvR9jR1xgnKs90saujNyAYfM1Wiw71rjhcVdVm0/5v50ibW+UK
aHOcCusxQ+bNhH1FAtSgCySCvp3j4rli+oxzTBvP4m/gaQ5iYI/HY3Kv8ZGKumgd
hKvU2t31Nek87m4NMrEVTP0sBM8rlasTlKwUVLUq3qI4Hxrikl6MYEjSVj+g321V
WgN0DtqXUCMgeID0Yolrjqx6R+Ik0IwztMWYR9vZGqxfVC3Vo6rvPqcfWjHXfLK0
WQnWcAwu7/GzCOKVmdICMihu8kG/myJxTwsUy49Qv2gywxj7YtTe4Sn/9mhazqc8
+KYLUhsbJtA6gACkFV6vaA3qet8o7pkoM124FQ56CRV/w6dipj6qj1x2Wh7InFG2
5TGb2YYfy3Jk/yi/LFJGrX+JwoYwFZ2a5JO4u65Of5Xr+PVS38o4eILP/SDqwhM5
oEWYIAVebRxOQ/hycuO3Ac4a/0FkFF/yovWcxa8nJG4qPIznc/FnsouHdjQ3APUP
knScbLgDAQTXNdUTC0HLj3KUp9WU3LykBAQwgIk8NZY7v+XXzcJjm391jkBNL6pi
FL8I1fSQo6BuP34dVNpejfQBVteNL0e3J608YQYYARi8lL/dL6wpFc7XBSIycPxg
mSe2Y4EvKpmJn3QuD2BDS5wgBp76MhHRVmQuDi8whhck/faI0oxnp0izMkJMCXT5
qAVEdoH/FDMVKL6Nr/Sqoid+x6e8gA9vyGAnIZcH6wAil/YR/jwjKDz5YYjsmzkP
LcBBMFNMV4kSdVTET11DRI7Ra8kVs99DyzWrnvNW18/PCxI83hRz5j5MPD9uLqJf
apUCDGW3SZXPDjJAMBMe+gqhkPGpPw/ics0fn/W4259m77eIZbMhNsoPz//FV5/d
KuYOhenh3xc5FYkV8+FQXyBiEAsZ0svE39jEiSZTjCvH993gmpn7RPimYlDdMOgS
zlhFUAHFs48IIeQ6n2MLWFaTAmTvdAJgrkFVKAEhersTnVLzIb/IJ0XJvyQAOn8O
r2c3yIQvjeQ9A7nhyj+rL44GhO7kpL61cgDjpoarzjaPc/KUxXXk3RSnmoYwPttV
dgDanKWgMFQ0EksdvVoDi21NndUYHyLxligSkr5aMbUFFdtBkpj0yNiuaGfX8CVJ
JHlnJDwsPKezs5DjQk/9chXNGOfvMz6KnN49YfhLBg6mt4GyetMDk55ON9h+wplu
VwLtDkM7wDz7U8cE0JCmrXRX2b8ctqWP6CHvx/IelvFCb9BN/CtpLPvgztGHF1o8
fL1lCTLfyv/3LXQIYUNgjZxn5I+4B2u06p9vzuf2VZZOJEPLyNjzHsOKjzz55ldQ
mehvzU0hWjeGPEn2yynHXe05jpNh5bokiYueh5F4621XJ1qT4AQBPu5FgZbf03It
HiYJmuSeCupAJBVeWeiq8RujZCtS0pREplq8tHxI6spMmPaTBuaKAN2f12GP2Gv2
pZHrAs+jEnTwVMSPiCNyNQ97VWBudC+pjJNxgoql10qRQHLX/bGoaH3C3XNljVYb
53f8LdoCXRx2NkfDTJtA7D4QU4DroQv/FA3niBGZZOPScc81AjT2T2L/LEDaDpMc
pN+SBBUpjt14rdITzZgs+Id43f4duSnFXGJUIdIV+ZyXdXhEuzKriP1MKNxs+fNW
QZOnjwe3y+MynmU9hcAw10DWuX0VfgRisJJ5EOIhOcydq2LWbhgnHPxJNNaAYrBn
i87zQk3hNmwkiC9a657bJX7p9DZOI25PCltMefxyTAOy3WDcWAiPgRSMtQpRTuzc
OQj66+hoLN2rbIduAhmqH9VmW64SWmQbbUS621R7PGH63zSWqePzBDsMrYFP0CCB
3cpWkN7PrqVFs5DCTav5wz1rYfrAezPgSRJpFXPkkTxwyxHGbaKJTaS76Ov9lMTR
+BtJ1/wKUV9LEk65ZxjJ2UqhDv0UnAwgOyOruPP2L+n2SNBriadt+eG0FA3iB/eB
A4mlhodcxz0Cjarc9sVD+h0jUEd0tcx64fxeMzgSg4hS2q2WzOIIiyuVkDmoBbe8
3KYEcksvsgrD80BZZrO+SEaKtZsrFaZrewwxYcjO7piVx9/hqExNDWXwarF6d5ky
tXDpyCjl3I973d5P5b6JGM+jiwNTvpiC10mADf0CWq3hiKAysECD8MLRNV0Ti9S3
Yzw4hjXKJqIfw1hLQ+oO5uOUGv4dZjERCUWxjDsYnDWXPkLIutI6PXgIfyyq5WjC
sokaQ5V1UH6WF4is/xqayIbFaszcOe1DVz/sCCzd3A+EaWYlHVV/FqGSdREKCWMG
Kp+E+gPj2mmHAIsP8+XMT8gh8sihpFgWLE0PYJvuOkiIW7xxrXWIyCEUefVz9XgZ
+FpyJ/IJcWjAzi8Zcx00vixo3xZ3h0/DqU7zBC5RiXJ4s9fsA2yUfLQFnDy69ZMj
4/KttQ4MKfhG1s3IFYHkHiNXzHAJb07uoeGgAqZ84O8EyubbvIcn8NFCxWfjD1GT
o8Cg4OtnM1RgUjk3DrvtO3To24HXpfkKgTXcPJHqi2lqPuVqjoAYUgnY4KmngGZq
Ybzm2pkaBdgU5c816tk8y93PJMPABvt095tM5BitJl+tW0EmjhfTe4NyDATEAMiu
dI9ah2cv7qWijfMfwO7US2tCFBxtCNPie0A4551YvoJOJB9bHV+ZQBfSFn4G710Z
d7L+6PVG9WDNXCL1crPAWmf0suepoPA+0nlqeZXLNUTud0pKA3G0CJi24sSncQsA
iLXJB0Ct3exteiiOjRKTcNzSaQy8sGVUcFKXEMQjmdLattywp1mt+SpIi/w4fB3z
0guq0BQ9SmtMb3GcX9Hw+zvAbziE4d1g5X3m2J3wFfMeU3vGIC3chhuiMu9Axyzh
/CcOtPVpdsQQlfWMuB2X8+t60T4vbTfUWZYaYsMniqk7aKCr75RlIjfcJ4M+gxzx
l/D8LA+vGNDKOJpFTKcK+4+dARNvfAQCxDdd11twzoQz7fbD5p/o8JiS2VYhRqq5
lN96b5BrV7jUN0g6FkB3iH5+j9Qh3igVGWYamCzW/tsQIzXXTpGkPS1vQPAa1rg0
Kit9QInfG9B+1UAKT5/2qi5850c0GuqXFfp9Odpa+R7eYGYvnG1aBa7OcMJwwxv+
C28dK38QMzgTia7mjJkA6FsICW3q2dT7juNxDOHhIbecTeO/ms5HU84OwNgnRJsu
4H5sM7miriETTPre2SmxA+74MEv4E+n40qulWnbkY/oPEJNvg2KAbE6Os0jnTWLq
9vWBtawWkgzx7PAg3OGX1aYx/vw2+6SbgkwzluG55vGlRfQPzwqc7PdnWrXTmMqf
OlJC5t1PEy5IKvc2B5Mj3cJtVEek39J3FiQBflnqwKBW6p6w6jMtrglspTVfJSSv
ObW/p4UhI2r0QQFHhpaEUk1vL1V1kGA7zjsqejGvae1B6K2O2X3eYkR0KjvFY0ub
pghiYLRA19xJugqNTIjY+RafjiaBVB0aPZlrxx16N8F0vZlJwghpn5TVv6Zo8Zx5
QBggccsVpIMKD5m2L5ck+FLMMqe388IFj/ZOugmaKKuS51I4BO2mlzHulkTl9DHI
SunSgk7t9RJcHF4/PVopxu9pOjZ4KTvFOe4zWBcugkff9xn4Abt3XDOam+1Vhafc
zJk0mH8da+/eFm50+52PXa/OaTkTQxjDVGtK9yF/dusx+L2XWf3UnYOKamGm3Jv3
ucm47qbVhX99CqYOj/E4bcLXIztfPaRZbeK9vFPuAnbF0qQAHDMDUSfyeLwujAgk
q9YFkUqTPGFx3mmUGuMSrU1ewU3LDxyE0hw4OBOl3o4SGrE+WGB7sWvGyoeufetM
dP1ZZzv37w6jeWCAzPuacD1c+RCrmqap5sZJr2eWVtBisYbRqLjkdrKLHtmuKmwF
Dju5iPy6AzX6IvVJPfaz7fPYYh1EbYfjeCXtPgJFEQTeDwKe+LARQTuqyVHfBeMF
qXScQnK+zHp0DvSBPJA66LxiuyO/lFUTg2fvPNs2O/VH9q1BNIow9n0aCSOPDua+
lU6bsdAu92XEhS1ASCdgTd5CpQEFY9rlicvfZapy801JHbkFv3iz2jdw8WJ1j95n
jqMCqzqEsqWcbb19+IPx11/sB9jNzWL50Ztw0EAcYHxZXoVaPsU75CjmKtGvrEXt
MnD6WQbhf3CDiwxBYfo72FVt7vl2h8py9UpoYOV5LupqNDgt8WpddDWGEGjzf4IP
SSt/eci0Q1MW90IFyZBZVDRLWDLhFTuPvxPheMCP/RiOmcq56H537DM9X4UDSDW2
9f2aku+LGphlNx0r+M5+2NIM0Noqz1Ka/N+VJPwiumO/iZt/LayZFuu2DBnG24p/
j6zImWg82x5Z02S9Zy5VWVmX6sPFoVxjtyGf5eZlDan0HhQyudgtVZxOyQB/51My
nAzdW+YYlbBKUYLQOsq/DIeE0NyPtYL179MtxW9G0cS54oKHl6zv9SQcAQQW7pC4
QHlO3s39AHXbun+DMtZN9Rt5ygqNBPihgOBaeH+0lRibGq61Qart6lYv6FzwF+Ff
d3fVaL1aq/12Q9rUIXanklygt0Ol3bzahDzC1hYtFbmd9hqe1eB5Jpq9KP5uVUam
3rucrrSR0dzcUkpPtnlvE69yT3Rrbugf0z16wcbxjh3l53tKIHl2pOhSLgOK1Y5B
ZcFpVMY0CMmCuDdDHLMQcV1/vaaW6uxN7k3WYPPfyYL1vth0tDszT5pfCerkFxUE
r90eABOx0LuJvol1Ao4f3geotiPTKHPhy30RD5yYWha4BBL8HkMDTmBYPPEXvKZz
4VB9548nIuS8EfdGZPuBbEnvAqVjTVL/S+0V/qFtwKq9DwzP7Lyz9cHdQCMiTQQH
BsWLY3Ll3rem9jmW921oeBLT0Zd1nTfp1z4WEamLpI+Ap+P/NJz/X3ThBFOD0RrU
BdwRq1UZCYv/r4Yt3TtzrePpb1tvPIF6S7lxqJO/AmhyuOVAeTQrqoMppMQJG3YJ
De6s/qPx29BnMASbnuIGjPn6cNnYra9yPrcjRSxnge1jMuicRQt4TsVyDb3XDjk1
JKnLsCV+4ulwfGqN4Eva4QBAkflTImQCTczgv8TS0Iho959/+1HIXiyrJfKzW2mR
Tfq1B3IEwlxDlJomBQAl8okZx859reY1w472CDMq0XaeRL1HGQ1J/xiIghihWL8Q
LiJhqSE7nWxWQSgwFRHRumaYGCk24rtMJPmzKOm7k/73nD90Bv68Lp0JAAtLIJxJ
K2dq7jaMhOUn5lFU6qeYscnk+Ds7GRevuuZcZIq6+nf4xTqZPmDvfNVPqQNalW/F
NbnGGIN21u2J4SI8/WnhVr3ZYUSTxTpBIH47OXmsT+7XsmbdmAm7cfBft6lcf4/v
0jgqIvxhOpLD3QXE+bLwPDVLfpuvyf3FfxRBp+7uS8gAKsObRs3iUqtEF91BhTs5
OJKfPnNNaqV/kzYjqYKVhWjTQbLTgFM0iL122hZm7YOxAW5eObQQ2j/lzxjpBTyc
xpohbjdfSOcdR5bXN6BWZxtp7CJKiinRPEi1OuMyHsvEgm9jAjx8hYCc+0WNKLKd
eIwZOFMpa4ABt5kOdOEhrUCWVDMTrLgndzyXJ6FUG5zFvKHNOCr/RX341QR69UjU
HWFc9er6cbjPRwQGJzGLQ+hIgzDZ9rCn9KPYNPJUlWKYSp4xcUFb7BH1mG0Jcn95
jsz46wBSPLnp6x4zwubVOk68JPKukd83P7BdDDRuwBvu5sMQqxJuc8jA3xfGETeC
a6qTdy2WE51WT2jS6SlWnK7GMoaB3yDRg5TY4Xz12Ma6YcQCglv0GVtunsrOVzFH
Z/1xBqfCYuezoeYF/xVu0QdS6FHe7iA3OjeUKLjnZavhsjPpNi6UTFUf7uOZYtHs
BbM/P/Mkv4yIClvTcHOUjkj2L/qRujVp3cETVVDKp6Ehd1SQ5ftDGgXH2udauZ0v
XTYFXr+FuFQgbPIEUNiWA4EmZM3eVyQR2PK1/2jeLVIlCEeZIwASZaEnJ8b+9fc7
S43rz8mIkCORoV9v1cAxVNxtPeACHI+uK5UfExFBPVzwGAXU5kNpnHAyzdLa0uSa
9pBNPN8oUfXIFLhM6UtSB22CNMzUn+H3IjdFLUsnGBczBeurk+Dh2Imawy1YYzSs
2AvSFFIn5atnK2qWVaV34GV/ZzYvWaQZHk5DU/aiPReSBGAOpbvNUyX4kGqjkMpc
Br/GGoV7gCT1YtgMj/wODQiZzKxyugdWuD1oCV+xDXxF+8C2BZabcBE6636rZOMF
tjP5HPGnzhYoKTdHA6r54K/YrtIGbK32R8Y2wqizQBI6p18LvV8Gmj6/HckcACVB
1YQT/R82ZFmvgyoGYqUYJiEEBo5pF29qMMBh7RNIi2w6Vcx8EO8EasW16Us51YN6
eHzih2fqePghTrc55d2gIMDBs7oUbooU4oYE/jYCE5zlGy7XoTfCRarLIn4yH2iZ
6oYvxcLHpTOh1n8g407uC1h9tpR92/2yuSzOZVdGoMmhOEb+PYGutItzsA7QYK8C
SsRoJ8CeLlzKCse0VzKVA9J+fQSsj/RUfWIXA9IcZaZm2K5Wfcrhzsx0C9HC/WoZ
1nF2r5bVkp3Dyua9fUdxqcH26GPu8z34Phug+xpI+MByZd/byPSZKT3784YYUvO2
1r0C4nS+rnu28CkhqLtHf2vPcl43F7vIkqIe0OYh+7DvohTtGumQ+zLZSM8BSn6I
IsU8UmiefF4ads9D8mt7b4o0/7Ux9feHKxMTNu60j0+5MrOjHs9AprvlJGd2GEdy
K9v1lDC6hRxC2P1HnivQFEY8JXvZHjJlM61mOQUU44lnqXxPlQZsRtn/cQiMS8E4
kcyGWkMfLIPMJEZL5Yrmg4PQz75ewWsRgIpk4l8EjqBj2LdRNsA0l3E+4BrDtapw
0RMOOmxbz5X/AUDCovIY9VSQ36RhRIhEnbpSKVse9BWMzCKe9lfvR09rgiqwWcRc
+dsFpU6CbbKTZRS7FoM5F0mCyaUPFSZ92ooLVrihZ2U7x3jxDQPNQ8TNS2hi5xKT
n5oyZXsU+0+ldBe/QkRYqZ8E/QrKALttuU7y7yWwTBdk5pgMN+uPimmzUhf6Mnj4
2QhEItt/mJASjiSV/xd5Jm6VoLMFncEeBFUjzmVQqfIPzJn9WWk651arGeGTMN9g
NP83X1/VLSXW4BmW+WQeY1YOAQSN+woylKM6JpkG32xLgNsk5YjiidTt02Wx8KzF
UAltX3xEAsVzyWMqZxVGk60j+z0FXPyycj97dLbllRvS02auZLeUvq5FouiJ9V0n
YQKGFXuXWxgcsD9eXH96MVOSQxmt+CBEfyiOzDafFFTVOt+3oaccU697gWiX17Xr
82FYvVHKEuCUjmHBb0DMuhrfeMyZUt6HnWMIz2iX68cxH4GC+faWHFtM9mF9DnXF
Eu/I8HXYMQOjrGHsmk1N7zhEL+zvRQGz49czitxZwOtT5Xfy/lRZKCjAuNQhd50T
naHpKBzaIgRX602M9gdvpEPzVC03Q4TZb6reXlPeIwJJwYXi0P3iF4yRU+NKAZEN
80kPCSpe273UjZruyLmYeaNM8ftYP/EW7yriGBlcZJeIoEIifqqEnfb/Z3ijThZa
NEVeluaIW3p94AS10O3BIP6DTrhTPKslJVhzTG+vncO0Jt1LnxE3FDH9FEs+Zsgw
/8SLNa+io29rg9w5G5BAo3NuuQOItbV0IR0yBwKdErR8uI259+AeTtOLdu8t6sL3
U5mnCAoR52NSA3J9ZvBEUAi835nGERDXKsrtR+xzDnCIQ3vSZd3d2e8s5pEIPvE5
yJJE0U2fFjwLB90w9HAWvK8WhXvaxx3QiGTXRLASVSHx9Dl7NfedDwQupPn+oe5H
jE4RnMW5lUv0ta/8Hmo2Qs80X1ekjUsv192LCsHVH+bHAeM+xhKxalxOicsugy3a
LbW0YeavJl4DoX72GKZTPOQzhXMBQ6x//CPP+8nCTti2Q7FzUHKwTEKBhPg4CeqQ
594ppfuFuCBTUkWP6qeOjtkK8n2ZXDyaCi9eFbpDY6FgFi7ktj/f7aa8CY3aKB4s
9Sp2J+sJEPCrmd05EJy3w8bgMGiKR08m2RP8Tj7+t64uB47P8Hx+cu7g54Fgdbyt
UwDW7TeKscxxhT/MKZo8rTf8+vnE91id++TX97lFKsxFHSInc3aVydQ3N28f0qm3
NGcaX0gMTYFqnmESc3XJ+1acnCD7C4Vz7TtLq9ahDpF6JMOdX4j9TFPv6A7+JkFf
aPwnpXP5DNyJM/h1sPL5qxyHZu6X5GE1Wp56K6mC3thX4tLKjTiccmyY01vhTLBW
rj7n/lD9zLriBLRQSf7x/dNGr5JMSJOscD6DYYOVVfoaHrPj3ezI8NoFO3/U11i1
Q8nCEuqxcm5VS55jmcjx3wDjv5xc7Jvt3IozFE2MF3XQGJi8z00yJugQQweNGQoT
k2ezSqAbXxJIzzRFaEKd/fjijd4wcgnb0wIBEnEVWfOz471720xAuO0HSQIqKoJM
e2KYbe6uuoI40U5qwfAyrPffKEFbo+POtdBY9I54kye1vpHTQ39tG23c5FM9ms4r
hsmYpMLYxt+7yD1nxwCY7dFLUh4qnfm/aYJdbLtqAmDXd02QBQsi7PHQZgx86Y+L
FByU390vxVJyknj4FmE5+tDj8H00qmsG3EDGlgCM+7E3J8jsb1UGnIkzA3uH8kWu
OeuKn1QA2JLZqsSUUzBXVSZsYiSNjWHWkqGNOSlgdCjzwB278x+3amjq3rztkXiS
Mi8nshNB6ikPZVBR6DH5mhTe7Nsk8DYDTKKz89xswhDsFRNkUwIQKf1P3kbl9pvI
9pCSkS5QFLZ3zw1XWMJgO8RprPWnX6+02IxJNoFzyIEDYUVBAOH1apzO1zXemIr/
VjR9AbdTrrICKVvDW54D9yqhIb32yZmI3we5p71VER7OXAwG1bEs7lqgurEN6fSc
Cnd058/1SoaMwtu7xA0aodgrC0fGO7Dsgk/WA0hdokbG3zmLMJxSuGSQ9FgsCiKC
+i8IfknHVvM72GH4YKWtvKxFvWa1GgqhPBURQLqQXV3iGi8pTVsyQlMFb0Aled72
FHH25QQcE1fG5DLJSuF2toNNnGbjvbym7uGFfq1sX1jNJAZ14TfcIaVtGbmkXhPF
L4MFDhx9dy+0yo3B6xG7WB3if0nVW+AZRJ3MbvU7M4varZ51q4oBrevKODk0GuoJ
y6A+4FFX34P8oW06ctipR/r2rnopO9rq0sQK/cQpoaxr8Y1Ha1tcwXkAMHcbbeQy
uBLl2VlKHvWsjMwf86AVHKkdtv9tAJd81Cj5aBHd1ngtFNqUmR6qrKyS/4YW68wb
V73tYuqJjMOnrSujtC1H74kxwpVE7uTRy+bEO82uQiBfH4gLuj2ROqtlKmkgvfe9
8fhs98ax7ujc3KUn4BcjUX/oUT2ZVFGbUIeXd26gDxjgm3EzwkOGVoChz53mrisZ
Iq7bIP827v1N6SWKuq9IF4wpxtDUBbg6awPPuL8MXtz8OrhKXvNxeQmUv5vXagQk
REh06EcR+/mHkgBsiHVsOIxOyfiwNtudpgskME41NF5ITmcl61XT2RZxVfeY7to+
XeXPF3eBaDsmc2WVHk8eo8NFsHX4dHRvD7Prt9pHZ1L/2CmBwb8yfKxa3k9ddSjW
5GSaT38Ip5IhEgjFcheaaqa4NGzlhOEVbuNFwSILZidFNhoq5D4tsQbtt4ZB3uQb
xLnxK2hRQqs0GZB7Vs7yD3v3nZz+W6O+F52knOkvN4LwhSFfA91/Jcfl4t7KxFwf
Tt/1yENUNXgqr6Anz1cV3TG2epDRNBbDFtN07c2ahQhfvZ+UHfkv7RlDPKpZVvaG
EybllYe8xziw5y+o9Bwkb2yuUxNL706CEn/UKtn0jisdvaQl0Pg9r0y8/SahqCiK
WoIKB5l8kVLf9G7glcLpqJYPrn7fHQ0eWhHlPcvj++ZW2vt9L0ZD5WdDAWtALV5/
YHS0NyE8gV7Gd2JPtpb/JpezsVJcnz179penX4IboW22U6yHAEuac+ghxt/zZ+wz
4OlvugxKmTxl/NWYoKXKFP1hF2mcRqj13illEDgjF4ejppHoq2U1V/f6zH/fbSAH
UiOBKj6+4UbUFSsKSSl0Mh8oUoKIXedNvn6tbB4Fn74rlB4ak+3g2RCkcfaGMYra
PQm86exWIiACD70cpnEJqKGZtqL4F7/7eOP1kkANuoeE1HLlk/LMUkr07CZaCStC
HQwN24kpgJcDTtrlyiS1QMJb3vryonCTSa8/aRy4W6TWCwsBBGXUruVeGUNhBcws
idjaFEDy72WLK9dxALjqeYOSd6HLApzuBqUEs2Sf8AXfqqYIPD4ITEyHHoLTihAQ
8fS7mVmjPH/lDn+zuXmTCAYbkNNW5I9Oy052XQInj5S3g6TYsoXAA+qCGzhOyyLx
88d+NTfrSinV54sCjmYt4GoQAFBR4Y4392ba346cszsLuLNMy+TAXPOFw0r0G+p2
M8JEHfcN06LPb23RjnwNYcZmO6JyZBMRvO1oLYgdCTGJRZUKjYytrSe4/zUyVeUU
IrF+GAc13CdnbbzoQSP2tMp0SYIV+FjI9gNsgc5l78UdLOdGgmstlxnEqpAEp5lF
kfZBodg+5FUlrUGtygoJbLb5QpG/T8QXE16gV2k/lozpApaftZEv85yJqcy0SZOx
AE1L4RhzYtADH/xT/uPTp+yitrVueO3mN+POateEPc253lL/b629H3VU8F4ajkXs
HVH2fsHzrx0iP1l7STQjbT5P+cyW7jD899sDDrxrXorZz3AKPk1fzNby++s2uDos
hxT7t7ruy4INc5aNkStDx++jaCmdWOHqpVys9o6ZQlrFhNWJTnL56mj1iHgT2VIX
cnWxPwM2uhKavrgItW9SBVH7++kEmMaqJ3bCH3L5Qo/x0KQALdvCA0naQbXfX1RF
sBa+PjBbUB2TzHwbBQdEvF4Ft+YXi6+SEguKRvyylW9jKPMVH+lw537allMNJ227
ikUtDwCmpeNZJUsr2k0cyFseYXQzSedIz0Fnvk+FaDodh3TUGCNmpvxvioMdnu5G
2A3HmLfoO8zhPgTNP44VC6GTBPADp/7t7nbkJH2DSNlPAIehfZow1/+KfEr/yVNb
q0ye5UzQ4ECkdKD0DXCivruCsrfM5zudS7WvpsT8p+5mnc7VkkllbUhOQhtMbUpT
PhbTPyo4VWJTsFJOExL3RCMN9mNDKcerXJNV8ug1c+9gTNnbOZuQCm3yHv6eIWHf
cI3mdJfQDr6vbvflsbm6BZSva4ZlfZTpg5kzyc2dSNNSQpNxcgQm+i4UCva5Jk/j
eYbF4qU/kRuvRDzgz/e6/4RTN7X8wJevmzeNiWU0wW9D3CPa+VqG/ozgIpBiOxzM
NwjwoPlV4mKafHdRa7M6wg7dPRlW38xunL1n5IsIYIIHzRG8/xqaRWtjDolaxFbU
ds7TkuXbU0jhYo88EY41mAjwFYrXY93cZrDtuL6b6ZiDENVI7x8xLTvNzsNzj+Bb
r3lbZihsVGeSKDRDSNSJJfSCEaOFvmkfPw/wSwsqy56AdPnn+zYuaSZ8MoNP/NUQ
nydOTa0e4z2UyOr1O/FqeGrKijVtaLzjQPdfkgRyRvZsUOUagFlKODRpSXYalw/i
ikXKF9cfZVkZuIHTfQDqEhTD8NaVCHTYoCCIXFPgKfdJ1Hm3qYJN3KE0yGe8vXh9
m58uOi+5eoZLm576ur2xoFKnNvqF/QxeE04NvkrN6Pl+vMTjp4eUMxDcKGW2p17K
J3YuZ/UnIgSRt2MLBJ5bXx4Z1OSl/A/m7vW68eyk05qr6kUWxxnygZXnaW7LG0PH
Xs5OmwD6jtzV81BFkIGIG7L8SvfRnx6v7gN+L8K3wSmuDwtx+69KFBgD51TV4a6o
3xlwloXKkoWBOVkf+VsD6gPcjCzRwU4bgH+WopmPbgSACMNUUaTI9MvuAk5Ohzdn
hmZfE4Z0eCa6vt49lINnfQH5nPi0w9p7ETYAwPnZnf6GghibPu0bwfWjQ3MNIX0v
NzgUVn79RPlqoP2OYV0tnJWsnZry3lpllAFUWqtLrJNh4T2p5OxN9rRRvFzy/T0Q
OQ0GCBktqc8/uayc2B5PT66A8oQ7Kc/HZ5rgR3Etf6l1FxsA8Rnu1VTl06fQqqO1
pGUzRKBJpqvd3+YGiRibCsYKy5BQnfJyebGpNAKKjIHidapOhJQTJTm5xEy0aBca
5t2lNrWLIvRlErsskDvaK4eAN4WzzlhWVwgFcIci2p/l8lhEi0wM0RpTR/rdNH0V
4OO3+Dn4vXkR2gFWUwoIqlkMq3iSGfwfzxNTm6oDsq1477r5icfIS6Or0dSxz//j
3230tGHvhpdc5urdMjTBnRvLh6yeQPLqfLqfuTjqNuXDxfWP7Ta+2WP4msayJZJY
172LtXt3gRW9Paxv4CClZQwounuePX1mcoZXxnr6evag1o/xyAke477xkWWSZl52
aiqorWgPs8Su7vXk7BcLxebts4D6ia6I0FYFsZ3I0juA47U5Or+JSuFzB+Jac1fQ
jKDaD/3tMC7KyRqyMG3lZl6WbK5+sILhpR17gWpluCXe+bSaOE87h1zpM3APaZEb
M461L/+2tACVFQdLIIQVKjfNWifc37r5ReLDN01cWfGgEOwg1eW8ECgQT2R91Zgq
/2E8GbJ7Cul7GvMM4xuYJ7oqiysws1gTvkdMiHXmUzLaqei4WqFext1A/qKMg/IT
ZQWdnctTWViZqeFw+KQxai9msLL99SRuDy731vjc6W47An98rGcLXz562r3PkcaZ
hpzUVY6aR6gXrHnwtuntpyjAq75NsYhmsW0/NdyKdlSIdbe0pPOQc81VTSts/r8I
3/Z8aatRUbbKk2Cii9QLNp7NASk1eq5jCiJTfIOd7FiK8P2vLXQ5M5nXeL8njfES
3CqSrr6NuYb3PL++xnjMmNNN9XX+kKIMFHDXOKbXop25gYCwYKL+WABE9vwUSK57
iWOnds6hdrcGjSeMPf7P5AQQBWxg8LEc8kwPBpKAAbhzlX6zXYsE89A4Y5IRVzT4
YD32kloaByO87KvLZUUkWy/jTzODx5Ntf39fsBqJy5I3lJf79R5DtZb3WRbuxmty
iomeFaBBTJdVAB1sA6zjg3Ed5Qbj/fbaGU1ei0RhoBzfRfX5uJ5rNsUA37AuO9Bw
KcEb8FcnVkFb5iDfxj7iT/ZtZvvPpU87Tt/Ht/i9ioeR/yYCr4HqTdQf4n9vVHvi
Jq04PyBAHiDLJeQ9R4C3BK6+yJyqBAaOQ4zU6svYSjQcM4Xc6byBNogKUJGOpx+X
MauwJbftPZnElTTNe3Tcpg6sOzsy1bQHMYpDimeCZ8qYNgNg6rB5G9owNh0ouE89
mrnY2M6Rrm8qvgLrXLiW9Scldl8Z1lCUNJC3BgY0Dypqc8db7kGyFGTpAxrObUnZ
40LJVa4/gm24IFT5ZZ961gUsSCdzr4rOzQ+ZDa1cnlbWlaQnSuUaPnFOeWVDb4BY
U04mt5inwRAsxN8IPJnxs/QkVQDVwhFYMYVm1VTBv/5/ttK65PhnzBNEyC9OUpcy
FnF9CR8xVQpCsCaVT/p19Y4Te/Bgz3G0KoAaPScnhe46+GzS3ik9GVauUQmSsYpw
0Sf4uescnYBj/lmh78nw2oXUB6toZ5u0cTavEz/D1wqj5C82MTvrKNXbThOTbiem
ZqRf6Jg2W2aip9NYD6epKNnqWknEmve9re9Yu+rfdlpRec/tl3TUNaBjJd0WGnMG
Bg0I8+QzDYqNYBXkaSb91MYQA6rzmLIrQgAdpzrJMeNTDP4onQTXdYEIbhimlJaE
Ex5xrtLiUC1H7nReKqSHBJkFBjudNKxEwYV4NB8gO5RF+b+d6nim09pJFomLZYWW
uOHLSv7dZVCM7ju97MNjJifPIwZu0bFAVB2t8zHspFSTYccGphgIBsNuc3WflzR+
3rEEudgHy7OCCOOdxbWd/oLBsPlBmMTwNhLUMF+zmwusuk+IV5noskNzbjctBDD0
otny5+ONOZok5YrVDwM6D4UVuFFbf12ca2PV8qJANq23dNmC8a16+QaEeW724ApM
aq93rUm7eBSFD3mUVXA37YBaCHIjC3rld/uS+sF1hWOlFenUHDlkHNJndsQiJwKy
EswU68CNFnBZ28tAXyAbLISPa43lds1548LFm5ztgZbxXcFWu5KOuXnTjGMFoXCV
KZX1Cwn1dr/cM0hYgVxv1u+tC8EGmY2kzIP1OfUqi/yyFfPc9C8DQR/JX2DP/pMA
bo4Wbu3itgMs8iUUsKtfd03clm5vlcfLXqbYLX8sVLKYFTs9DlNeIgsZGkrEnoev
QQ8Fk1txzKNZCxbcsMLGzmbIngKn+7TIg1r7DNx19tt2hIn0SkwPXkoasMEmOHX8
wtxgZp2OnrRbzNQIA3owFNC6A0O/16nrUY+tnWo1iWrH53rmbVhiS2z0cWisioom
T/TGtqIAa+d1zgE6T0wllCTRHVm+chWCwHgAmga+alsULEKgJ80onBts/qQr8HmS
UvAjkgqe5L5dzn2noDgZ2ZYXnwwZUNpkmjAeQ/ac+3YySAkok+WCawZ3+kYHdY4A
HHaGMBdBkOwZ73afLNzKFXGp58mXf7Hq6FIgPlnEG4pa4z0ZWnlhUbJNeXFxPRb5
vPLCtwRSffd6QLnH8ourMnDkxDzp7GJmYczjuO40tZeDu+i+VH+7D3Vlp2sDoHmt
jv8WSxV5cuQ9PgPFtlYF19Mc1aXrsfwH7qv+Fy0mp/GHDPZjiJh+K3fLnIDmZj5W
MefPEVkrryOZFMOfOwyq9LqHEuTwPLHzqTeGER8qkc2zSTs2/BweVAoPksk9aqNI
fDfTAwVcUnVBRMmhKGNul9K2oOr80y0MiCIcbFpTbsbisKNZpzwQQRFh93VAnJ2w
RjJk3N2/VXvtoONaHf7wV0O4pTJLOSJ+c+IMOfL9AmJyIX5qSb+EXglt2fZU182M
BZJAtFxxIOtoxN4Mcbu5BJrITRUAnIgv+KSaZbHItybGe/jZrAxUi1JxKbfTtQJH
FTD9nnu6kYBKVPT6wEuSujkF/VKyQjjH2Yb0e2VKndfhINZDHBQNsQXzSeJqlYY2
05Mz7rdC9TEDXizI1CBJDCyn78nLlyzlaohD6P5xvmMWVikeCb/9YKWpetQnHaFY
fFQwXFlN+THJPwPwiO0GStxxRug8e6TnUnMRjL0yCxchcmezQBEk6TQSt0UHvJX7
r0RUiuUoc2R76hRneIfrqBrh8QipGkA4ZvACqpfAYEJ1QWlF/WEGNM+6d5mQdTRh
xZjICb+FDiRzmkze13CiKiv2LDAn9vzbXbMsHCtrcRLHk4HOv+B0C3s7x/WS66+D
U64zbUbaJcp7UnbGgf1oOWvXiJ7GuIkk8DU1x3rN0GYwQZm2vHPA1Su3jG96Ri81
wqAiJA0bd9F8IelaEzLwHygqFHsIG4FIw0yyFo+jWzRZd9ElkNLh9y1g0ennmK85
HrTQlCX7eNikPh6Q9YV2cSbUOR10D1cv3KknzCmHL0vBHt9tvdw4ySNolYgtFwjz
iTlmzl+D9zZi3ucGhglKYO3nGRXl3bxlSXz8rmkOSJHpT3+azW7spLC/SUIch6xP
94+R9EBjZd/7GCCK1/rKZ5H2YBn1424WzefUql6/gtD5+ZF0nqP/IT+00cJuwZK1
tB52LKJa0esUYxK7Vwq9nuTcWV5pktR36nwYc1tgq47iPsNUBsGtoK96xZbp5nRs
FEkSRRryfXfuP0zDhj92kE5mnuPHD+A4y0TiMCOWSkc1wOzdSd4jjHX1dDOq3Vpl
OmyR6t7voxlMTLNtkjZ4IEvjSPfEsm2WKjawEztx0swuJhQ/kq6VPdRimr6wXfTr
pCY3KwwYbsqIQxTN++JdlEDsh7KtDWiYiyesyRGq4ouXylQuIyuyQkqYxynpCqqO
PDxxtdD0PpygYqT0g2SduztJvphYFCyyec5n2Xe4rBhiQ1w8TES4Tr6rUpJrnCBY
jiEQUt9HQlGERfnxmmtbuVB6rTnYn2Cyif4XFWlnjocr3TkGtL6rr7EKRjDcXTbB
SDLKAuOUB5Xp/MjOmsSEN3F0syx5yjlTRO+wCAqRuq7ovNonS4B7zWUyOtoSuVS5
eKPibZ8DEnTBAtoCXwNvHoiLSPovr+hoyL9p+SjIxh022xnq4C3NPqBbwRGffH0Q
2tGnnZgy5xitDD7Wyqv8D5HCqblJkTitAjnOCIBeBAHv6WXbDFd4eEb5ia2aMBP+
Qm5nkhIteOiGm9v32ErKnhV8KL/lgDw0IQ6CUtRcRFNuuRZSYlJ21oCeSpW7+6ad
WE3v9KgcF16wwp7fbz+21zBRnI9ISod/zSzHZxRHicI7EeIzTlJbp1kCHcclTeJA
zpUYXqj/uqsyYV2Dvih+ix+C0gQcjLX6DG4Ua/c7BPWhyJTvi3sgdax7W7+CfDor
qIbYWtaOoz2VNmE4Y3lAUVVlSedqcWvn8qgHnMntAUPhGLVpUPxEEGLy7E3X/hJt
cJyYFAvyEmYP+JXPmXz7nUG4MqHziMYI7BTnVTsUFUFuZSWzdO1zwuwluyW4q4MR
jvp/TFx/VkLVmnCId240H4FkTowzP3Kr8NX6SQYPI5U2UrDXMXxs8lOgVdM5WZNd
3QrXai6NIbzw8azPP7X80aKZpu2zJQG4E5AZJmtADZZk2/Mwdom73k3IsRI4+svu
HeGw74WS2v8XPpoGgZlNJWdLJ7NDBq9wHZPsjQjOs31585UU3dbUbJnX0F7MeZvp
TctMeW9Hrwmt+N6I/+WcMck5fuOJN42yuvKk6yZdO+d910hx/ptO2bJJMY3AucsC
DNHOOOD2Lgn+UGxQjQUwgZ4JDzERDmuvMsUg+eInxvkoVUBg/Cs3M2wnvdgntJA4
efSBr1R80Fv78sb0uYzEKOYEqQDArP4DJrLbGi2o4YAo3C07q2oX0ZO+WDXXdcP5
fXKlimpndfSXqrW1bJYhhH0LTgfeyYBf1EqXH8e8nH4a+gUjh8EjWc3XDLBuyTcg
5SgC3YsxLNXSbafM550TpVTL+s6GY5qHxbv5HEcvwhQQ50SfLxwNlJ27XFVrOKPM
cqjm430ZR/AanJ7n49Mw+RW0cIsS6ROlxZBSYNb5B41bp+xxDpAS1jhEabedJdR1
bzBI6UIr9Uq0KBoGvZb1LO31ddXLHqkwtQwC7V/wa6iydfLLiSyGTIirN2POIyPN
4Wxkx6F87ESq1ZsLLq3LlDT9VRIPoyzcmuIfLmCZ1w18eeXDgewepfx13nV6Zf4R
MoADqRsim3zze91RI6Psoh0CiVVFCfPEyUDV8jPmi/WlJLBRbvv2Ba9LK9h/A7gx
nvFlibYC0YHOmUAV3pUtMfLgWzvcoigLNgbcAiFac2iZ+DKRuGGJOEs4sHYd9T74
2GzgRBfdGYdISX0MV1CDGn95S3sx72BoSw2oo6SjBE/mLXHK+YGOo2TZVjbNpH3i
pnpEyYKLFTnbkpGUSvA0Nqh4B/+kiIdA9HrSgI1f4JEE4Qw+j+6kI2aZuFnBwGbD
7L8qP7Ne5uJKSLcHihbZqMUVUc/td6CqY1LPPrR08HK4axnrNFjo8T1ivLAjuLUa
kvgU+Thft75nuTeCVp/j8uz7BIUR94rQSqVp0iFY/ji7L4+8zfvc3s5E99rh3p01
3ton1iGBM3u/4piVIwhe/AlFofnly0969gJBpzkvNh5qTDBJJYOS0otp5hNCufeq
JgYHj693vyogFt7Uwpq8QyJAaCAzwt2gtPeAVPH8Ahst1HGfoLWb1mP+h8lU6XC7
psw0+N0jFEjPu9AuWh/Wu1EyAbKwVUtO4uObovklaH7UoU13cUjJhnSdQwLc8E6U
stT804zwmicqZFgerey2uE3wFSCr7WMFSOvLG2BjTiySDVcUW/qif/MNzt2kDXtt
+1avGv615tYpbrYHcaaIcvbedlrGQ54QjUuB6yDhsJRcbKzO6jViivlmsLLld8tl
OYpLKAo5QxTPKI8C2mc6V7iobegkaYA7kPYVv1tlqYCDVClU3L9olKJzxwC76ff7
q1qdPuNNwKCZ6viCnc0lMN3uO8QvPOST2kF4hHLnPcCamlO7qauEIfXC1/6HCObE
ymnwfhSJ7ftwCrVPYrDTYMpM1qy5nncpIPXu6xFrQWtrIh+ML/oV4a2qzGekeOpL
I2WmDlQc4w0ybYFA937Zt3VnPtgEatvwJaLuKyX9F04xhCqvpSpC4fuZnP03wwYH
mcLzH7xoHrlD4kDEJfVyib+wiQrVVXl1gDlaNQ+1UWAuOaHLc9VneBSTEynmyjXR
4ixnnUR6HAHOcatpApib3+BMUUxNlckE7xb1W7Jso3tJ3aiRr/HcUu9/YPH6XDm2
n3jW/oHMNbNQ6bf9R/Ph+L4TvZ12Z7O5hvDBneKBXnoVe3dDvOEOfv+g3x3EPCHH
Dc4YHb26i0YHya8U60Niex1CT/eJRBQcesLOIPZFEVm3+IW64S7EktI4s4jVHFDD
LRGGPy7GfpMUPzI0ry7D794ifcEIMbvt0bdBcl+LTiBLK+R/T4jxNNuUz3vZ2N1A
VG0Zz6MMD7bGNWzGuXPLxw5xQWJCmWFCba5Y2Pj3nxLiCHOJKWfCLoowBLj8wAeo
OqBGR1iMTrE7ojjV0AY7QYHcI1yZlDekTPMU+4RfkiivaqhaBxaAsOEwMKvNFntQ
GMlYV37WN7O11OwWbHk1PPSLbes/mCIj/XtPnyAmQ4QqiQATFyLr0NiLEjH9cBnR
LCzmzbBzqsw9BnIzBEX1xR60wUDI0BeDWMnuDkvORAdBRdcVE2LFovXvmaLUg6lQ
Lg6gQ479XC1tzFY9SClQ0i92tfkvy3Qm3cbE/RDsOTLmemt9ESnOB1vBdydwBYu+
DS4MflVL/IKdaLtwVYnsv3X7JyNDNS8rTs1Gemxhi/2egXScDz4T3xpcoxOw1hKU
rVhsuG8gYj/0ua9rgOwHT3pPD2droZ5isdL02wEjx8yVsaxTbddCz3eKfbOeHx8b
lhTVcXkH/a/L1tUyCSfsxivJm14IrRerHP/jiseoDZhG1QiDJgrg1a9OCCWKXCdA
l5ZRdzVVThobiEV9nl3BCT9yZHgEa5cT+zY1RGEqi6h1MkUmhfeamMyYo7YtB8jy
yhXUkbAMdkjR5N0OQZuhia84brtoXU2NBe/7xneobKCoDI+moVyWvepuYKPbrV6O
5FJdE2DRV9HLJcuuN4awrrsEb7Kk+83zN/taP308y2Zi1S1y6NKNV5gBb2GriLID
rMGWRdtLnIrc30pJR+Gu5mjjFvoTpe/Y/CoSEdbxKj0H2f2qtoA/73r16uev6DF3
wNlPpczFBSAbmrnx2IrE43AjQLLB3mDixVMqYLo2elIiwVUYAkzk7pHKPdLXbd+h
v1K/zgKTwUddYDVR0lQyieYouWeFAYEb31mTkwY/GeeHlh+kz0nq799fVCxBmrWd
0/+ixdYSnkZTIziGF4XhIpMrkChe2+Q/wNx+e1T6kFQSkfTD4mpANK0683b4eOgD
3KHShOtrrq1eIypCgLcZfuMEROc2qWuXolEPQrVQrIZMkY3CMrp1k7wtMUeKTLc4
1SfAXvKNUr0jmgcg9VmjCiGkcMynXl0OkIL475fN1mckxZqPhCRxqhDVY0jOz1hr
4/f4u/nk8gQSMtvU8OjF8r57BM8yse0ott1XqAA8x5Kk6MV1oZtMJVnQBSUouxxd
bPCvO0Henl6eeF1N0lzcU18ROA9zZ8cOW28fYU0l0kRTjwKaXL3WrE15Ioyglwnh
ehXy79dWpsdSQ2Cfy/X3qzvNLgbNOfmPC9oCKWmhqMkvDC2hFz/5HFrkk5e/A5mG
0tAs2mzoQvdmIol1d+GGp09Ha24lp+E08F1I23eRC7zbSEXS+qZrlZa1ML1runEQ
GQhGaJ/GSpy6Dr+ReztK1eWBcIJ9Iwd3OG4WhLO/nHZDQ59mlOaNt5F9uGXP75ds
FCTxzCxrR/a+hP87DvLEaWAZzLSXzNrBRnP/7KFFaXz7TM+9Wn2R0tMgnfMviWU+
tbGc8rPMd2V4Wz4JpXuS1Dukwz9ijI5FhEyUjRcsfoilvfvzhrQxeQrMmtOILtwY
bKt4DkbPoDvgR142dpg9EUZ4DPwlzGZlqfNCyo58b0ycTZGrNiRTYXadNVMJrVEa
2T4mCJoNoWEOECKbz+1EIfmKhjFq3Q3SOOporq/yMKhgGObsy6RpSZSAMU4XpFiW
xgRWi8vZdjtyet9wYRllZ8mwcm03XCGAUxpUh2JVKX9zgqoHxejqhg4dWV59p2v3
yyJJXmIrWr3sNVPLTjQQIrEcLPnofkMpvWA8U9WieH0j5fitjXw3hTCltEWIozAE
xQdPsZlrJf6r2ZitgHtTM2zQj9fxNZVTKiHFl9bmMsliJAfUeVe4CfW7L7nT5LAk
aWEHuUd90GhXW3L2KqR2mPZUm8k/jyAlQeK6itMJ+JTJ92aQG6DyJrcK8FgxJMml
rBNuxhwpyb9iI7Ov5uhQg6oZ6gaAmKu++6FWEQvgT1Kt0YZiRGQiTQwr+YK/yGtu
h+H8wtQdYcrqWi5rEb/Vfwar2876MmNzn+JBHREvBwI4yiU+/sOLHi7wt/lYjMkR
CKaoDxyjl7iLhBSBGdco+9bXwx0laV7I0h0sDA9gyXow5iXgqQ8YpnR8+9lcLjU8
Gf6cD8clMU+qToEV9m99gF6CHDBITwNMSaNQBIyqqI3Jl/x+1X07Vs7u9E/kuwEl
pv19OI89gB07oWfaOBkqrKyI4/iMifpB8GniEqR0Bop1Y+7TCVi+bXyErESvx7bG
DU2XTXWTLASaWs6ku0BTO6qqa7slTkLxkA5ZweeRxOKB2EgAseIRff0lKJl8ycS8
c7I6XR2sf1L/mVz+qcuOJZ+adf+JK+TvhQ0pxe+Eg4bjhCbKc/wIPcrP41EYfRSj
//Ta6770z655h0dmwNqFEhObErMoANSD07sQfNHAmuSSy+tfVYNCWR+1FroLDhPk
81ZETJyl5g55lXUleUcjMao+AxBrovF4yZ7gkK24Rr7NvudJ2tXBOmuPhZW30pEO
yW2fDg8NzgDVf2NnXbbijbDgeEeWXQAHKAb8fKV8QoX7f7umIl7YMrCvB7Ec+i2z
TEgs3LkSTHyYYYgZNR3nflMpj+AOi6GzsD94XrbxLvzsVOmFFz/sKHtCv9efV4NZ
mAXI7dR37+vloOKziB6u7vq8T7YiqKz9K7IT9tdkZuthf9Vwv5Z3EmtVdE5X7K4o
p12IBjeRaFvrD8SRQalkLxs8qTKCpc8ihEsm4Za/gsv6N57RA0tOohRer+dKZ2eD
6PGXHG67Rko46rkMadUcjGEb3Xy0V/3lJLKdueA7NoNBSt2shbMLaDzrN/8ow0p8
mnzT2aRRwTHyX4W4oqYOElOo3JbEEOJ9fKJcqilzFbdpA66QWjF89brjisnKkZC2
lQpvYpkN20jk2UfZB3kCHs4u2DwNNSJKuB8CLNctGPNK+hGO2QEswDoylE+pbnn+
9itKWctVLHwJh23huvBGMwOST2T3+mGpwY0HzCqy3sdzz2iMB77MTc7AV5um+zw0
Hff5Qq2DSDIEz4c6Xe5RGu+eklbS+S/kZwuWdugsyKtZuDvOB7d9wW/eUBVpj8jb
J5KK2enqvzB21gozKCmqFLOaOFJO/zkH0XWXqqpNf+9wqOY8WvMH3ejqOAbjTT9o
CdVYKEKZDpIj6w33jx+bNrBAlQH6ej7vNBA4NklAQqk2Qci3HfC/HprHvyaWr9Le
NxCQPpk0VY+q4iILipyfZmZDhhffNGNzRpv7SU90y43sdoPX8uIimQ+rUlxBVGrC
ZmcXPmTCcp0qjkWXTWrVYXxsTagdckd/983Fr6n2diBZ/B3zI9jeL1R50ovs8N4z
hQORn2EBibqJadyMsr9JJ6L+ERI7JFsb3jom2q2je8NAPvVOf43nnhWTZ2qBVnio
/CIyW+NkgSCw2q4qfVUfwU/wKECo8/UA61zMslWjEEXnJ7bzvtD6yS5Eq5bViGNh
Gq316POcZ+sfd8uikMSBWk7gTe7SsLaxJLxlW2+2tolgTeF4paryRoFt8CRZDgV7
dxnpsf81lKkJSr4aYSv497fzciqUGHbWS+nyzbeeNcR2IIba7ZjZ2z6+JwWUlYDd
2TRdXscw1xyyYHXXo0dtanDgh7K6ePV3N+lsYzZ5QaLn49V+WKHDZUgHq5T3PbWk
37Cm1mFD3Dkvdpp2JQbzii/ZiQTMige3AmkbuLTHN7BN3oqdaQPlAXR2qBc/gUEi
xt8HszX35GRKwrLjYdB6pxjhOMeTI6oPE8mrVOId5LxMW7O8It5DMoy8T3MAERRs
hougzGkhMXbM5asW2Ouhrs+HlV8pDcNz9VwB+YG8WXdidzSZng6bicoAwuvNJXsf
wYmQfAALHZ9rmFSuToWai+Cq1vQSXtMDYPBF/ciEh9wwC986e9F1OBmTqSmsy0V2
Qr6X33J8wLrGdX/loYT3ppEwE6iCBf8SCAkLtIaJK5dNcA8av5MRcjUbvhNrEOw4
glJMGN0FF9sP1wGWj5Scb4ofirzdTE8nWGQFRLcqOQRW44n/s3XB17OxBRPi55gK
kje2yqCwD25/MDiRkbvfj5Xqz5xpXIg5pZ711SgiCrkF3NycipJjXWV8ax+Fe7hd
D65lWTPPKYADfE/x2nQaUMedHNZQf9xny1gn895ln+F3kmYq4HK6wukIeGztCGxL
TeZswN2d7LrjuFjyDCTTB0krZktJAAGjv/Tfg0/xXCDWbyClwQNyLSQVQo3yoRpV
0KKvX7BogFOGSrOvyJyf2f6js8CKbvAtSlVkUOyHJsBeZc7Y8xEKRzYSGnPPfiya
IHFAInJQSqc3tohRE1tGiLlfl9WAU7VGq+8EMbYPJh0t4XlJwE7Dq0KsfXcUppVV
W+lA3rs93WiBUbzpHstS4R912Al9Er5Ne4U2St/iGiLv6QjXv7wScKO8WGV0UMQf
lG2epG9dQHbPQScLR9YVWFQsxcFW1kzCsSeVBlDq/1IU60mUo7S8m+ks/psGhD8+
gYhWjefPyYHKfDcFeF1iAlTTCAwNjpi+cf/BPK1xugqqaiQz7kOryJQGfUTXAdjF
KVMbsNnlXsGLgRncBVCYU7xpyFomJTK4nSciPj+BGqd4Zj33chVvdpRyJDagbJ+M
MdfYioCgG2h7j0C0U5wWeRmQDtoV17pdnzTdhvmjcKdtM/7iJiy+K51VA4vcNk+B
hazvX44xk+OvwvFln1NKuOGQ0IdgiQF7ymsFNw0Kd6CXx2zXSbVq5clZpi4DMIdo
gOZzsG1+lC3OvQEXELkjPnWJPzUzF7erqUHMr+5OpcLfCiUYfk372tz/k4NV30Dp
zZf5nqlvEygiJEv2gitDqdXOszt1/bJKNIIwR2XGyBw773hBQ54HM+qZ3fP4HaR5
SEZq5pa4v1G/fBabsd47DifUA031wxaXG55qQ9aqOeMb2YGXUjG8ol9M5UMEZCCu
LO3IrgfISvy+FPQ0L54v0W1+dLoVLSzR3K+pqmB6VI892dkNl/n2tdMvwBnWLaM8
Lu5AV3UrK8M8wqzTqp+ZJgJCClAdOlenAb9MWmURzZf3/lGE4kgB+Cu7Vl5YL7im
GKQQlUseZSUgOriwGnKasvbSZ6r4L8Q/sQKq7PS9WEvGsK9DFFhU3mE3atBfXmJ9
eDVMkB8fvfPXQ4tIBNkJwg6ocyRj/bM8aLMwpk/0jqNMPyf7B7zd/rUMpcK/4uKB
whwG86ZvL2I8UZ4KAN1eri2IZqBhI0tmvGo2dYzhRN00OrSDuohzzN0Cy6hEdXdn
reAX0HdWuS5c+s3VzhAC0KZZvpd/u0L1ek52cSj1FQw1w+pCYE5ZqvF3/N1dKnOA
wxxYhjjcu3ivBsT98f7b9NzQgcbNGikzhg04ORPJJLt3l2jqW6fsGFcIxOMLmrBM
LB++lMjRRY5Tc0Mwv9EbqSrhEHQQOKl5PzkRWcKmvmYR8eKFKTbkTc8T8U4cxycZ
lvSqYXX+ozMTsF9yS9e0AjMpvn2La+jNe8ZyGiSAqVb/OED7+KiKiTImp6fQvhpc
nH/YuORXbI4P3RSWP2CyI2TJdgOBEUMU/4FLMC/GBP4/ylSNcyysnypKehzp0pMn
Ma+ypTXCIBl2uooEhobcEr+HP1q1KpkKG7LE6W4XwOJJMDNbgU5lOEt6ICkwy0QR
yJLVUJTG5FL9fxEXz7o1Tea2kAtGIwAEEiHQTo7UumV0opiriCwy/IKSI2av1kXL
dmxzx4ebTmKx2VsRsT9sy3qiHWTik37Z7L6P56juLNszxVtRZFENYKGkCr1wq5PU
9UjhMpZ5w2BYtgCjrBIa8/OcbZ8JlyTaW4JzjUHpqU2gkVtVinkvlDB0965L8GWn
6Sa9eNS2J6hXWyitL4g9D40Uh806QMPBot0NsUuvBMYs0lpud0tkFTxL3M8bLW3U
jOwOBv6vtu/9sZA6j2DaAFizq/QZp7/ACqjzsdUEsZezh27IMa+CrAhWwIpF3hOv
5+yWxP/M66vvGPYlTAmWfP+uMGX8C5diyxkI3J8cBybk5pS8a7Mx4POQKjk0UWtA
2/76g+ld9GXf0oW9olC11FN2sJKFUa52Rj0VOYZVDa44ZERDvmQ6jTZnMjRBPK8z
7pPt1Sxi0IjmieRu4pS6OcJAyH8mA3QNNmTGE2ET/Ix72tkny3XrL1HwmqIMTS84
H2zfT7mMOiFQlEp4N9UeDvj03kMPet/jS1AwkO7lxieXL4i4JgNfSbsDslD9UQKF
nBZY46q0sx2qjzQNBP18oheowFCwt10gHoRbNiomJgD0dobz5P2uvIDae4wJ0gqE
o/3nweJJaGS6AK+BxJZj+FZWjZTmfyXWfU2ae0TjHaDMaW+eC4X11UWv39dLN/wG
m6e229S810I7YBUWASScSYen5Jteh5VwnBL4GRMHowW2lCwguDub2wFwwynTaV9q
5xcuw3yQgeUtO1Cd9TFvWNDN6ZKg/WzwEnY3sI/OJ4OwsOnWmNjGmssAGmyZPDzQ
jPW8US8evX8DmUsqPOfdyynnOoQxOQ6blp877rm8h5N1PAwkytHdON3xWW4P4LkI
ht39lJEHHLZjGz07EhrsLuVJRt+52vvZ9DhE559SEGin73wz6njS+RHnGvFCw5hi
csSCrPxvHrQZY/PXr3xT5SW5E5FnWtyibvOIUBbQHQX+GtTaQTSM5GdAL+wiivHO
km04ft6BKAyjezjke9OZVOjXDtgCr+iEk9tF/zAcyECmC8f3K2WiXzMygON/DnaZ
ZHL016LE8rcGTk5pqL55WqMgwGPzEMdQ2bWFJ0YA9ur2poEcwihQeLGKHmdGfNq1
GXfATHW2YA/J+b8gqbIaif+nYxU3J1Ni8EqitUQQ0bh//1A62r8CGI3hCxt/hjqL
GttN4UXC/IC5pBzmkA15j8AL7D8ZMjhdM/Ka/IWyHLG+0+gkYC9psTG6ctd+ueXr
V2pNO/f8c9Wu18RMdLfTDwRL6MmLHkBimF9OEmd/AJObh0WWv7uMeakK4MptoQyK
G7btma75P6GwAbUNp+EMShUqMIwk3A3cUcaBNmyQAYoxcgg1sNhMVkOGGCzbpLWQ
g32Skpn2LuOehJW80om+fOy3wUU28YmEDseU0kQlhjcAlHgQ2so2B5ZPoL9SGpfD
hVLt67XcjCZBvXczO1WXeNZzMzPyMMphDlF/FWCVHv78Oi4SWKU8OR+ZSBN8kTD0
fTLCPlAKWH/Ac3Nae1IP6SwGo+5f3cogErz446ryrE+Hp6p/a8nKcWX0fZGSkRog
JjyHSitqnRq3vxKffEbshqh7luVpzD5Tw0n1sYvh5tX07K3JJNF4XCnF5c99yTcd
qDf57xcZKrlKybkMDb/4jx4RyM3IotGE5XhgFoTdqtwMRK0cljzoUaQztZHs84QY
IcF25aaOLnru9W2Qbfh7MeYtY+V3Q3dhwIJAWGT/Yc4e0JdIOyM8CO/bbNUhz5jo
VsDfuL8zxKBxf1J93fnw/lH4IPl3WeNr8sxKIXsIhXTGhvKDiclE5Wj4Dk3t2Qah
fPGHber4bLykpZaNNTVyddvsH6u4EzZKseWUeQFONUvzmekY1221fNFkrqTPiuPv
0cGgDGHtldhuta3hYHycSPTNu0qY4rSv+78b/zjZ2IwCFJhU2Kp0WoO+4k9KbDSj
4QB+99kEHGWX7tc8z/D8qqxfWxs2CM+S2ziWxBp2SkB7Yn14wmXL6wikZhMim/v8
vp4XilWlcUZSyk8+FtYCUeN9V62G9NHj7XCA+RPNkvNaawumDN8dOIpMvEq+rFsS
uk3/k1Ng/b20a0JtvkkbCia1AMszOnRtUYiPVflnIZEnFqx15BB2uyq4ZmAKh3oi
nZvgZA/HIfhpqnrUYROFzvRK/JFWzS9mTofGnAWOmssljhtv8aUCj7Mvy902gGLZ
rOkM3UYJt1FN5Yq7ZqZRNT2Md9ipc2pD+4dUhBoQh/cSE5SOmmgDfAcKzK/1GVrI
a+XuWmXOXO/92J12cMIJnIsMWq2OxtNsRVwm8VYBlkOjCS2l/2zF1hTIDXbpnSXS
KN8z0MYFErncZtVNpXQZozZXl56nhvPMynDVfIIyXf5L2BoT2Mk1FRxLYF4zTix0
L0WhwHcJLuPi8ZKJTYxFNWJlC3pB19ZZ+7sNHoMlUDXzm3n/Tp2QQ+f7vtP+EkOD
xJg+RNncW/hQ2thNm1GdxEpz5ewH7PEEdvOVHKt9LSfnphypOQyTMruTpbNKUgde
QWX5ZqoLe4ooYKpJ+Z20OifByAVKrU17NvqZQvO8XAP5DRaLJuOz9ZxhmKMyqBac
tY2KczmGQ9qoso7Sq14JZUOdHgfpnnxiBjC48oBbDQDIIywNvgmMXTfI4YuQ1ll9
YuGF9BHZ11zPncpUn0dKmrcvVWdwNVFBv/EYfTb26MVcSiOlOkA9/K9+R4xKZyVd
5Bn060VzsCOhWHDEoZ5f7IPV6zOvdpyVpqt1hSQJCOv/yL8fNu/lgDvej3l7cv8j
MG3opbABhKiIiPZ6zB/u7oSPXXy1YSG2k/B8Dy+C+VAqPZOLakcBu13LtO0ClZDD
dEU0Q16nQW02j2yw/vUz/mHkgzCWO65meZk43ux0HlxbdTIsyRm9GHI0R6zOWgFt
BPUVjeeoxF0hur/W2qT/IymaGrgnwrvdu7hRQF0WxQWRqQFQWIpPtwjTJ6IdWmyI
sDUzmmZIBB81tW/cKYl66rPYwkUTxtHfv0vn0DON3cu01ZbqcajvKvE0Hivp3Ane
8P/EqfylVeyEYsR+JLF2LMD5S3aLTdEHQOuhZjrDmade/+0nTlM+zw9mRluzG6wU
1lZa9NTwBTYxh8iuYQ1OEc/aZUbGY7qx+H7oNasRYmfcxnqjTWwaArA4ja2lT8m6
/pdA8/+4HMlA+aAsucRuS1c/hKwWqp8aHHqZOspwEaVtSN5NYvgy81poLio1M2Bk
LzroIU5MCVI0RQTFqDNu38lpCugA2j5bPNqMvDYR8lCJ+234YttH5z5apXY88n0c
rp1BsDN57+c7a2ojmWFA7lWMfr6MWDAoWQj+gyQ6jpjOpNyn+lRAFDdkymrzDjVd
+5a17z0zrf91ffaVrrJfCPBRIMZJeKWc3Ycft6A18+ONGyIrVlUHqRIojMat7Xo+
4MXDjLKKbdIe2FQNSUx0CJQIBGRNcFlFCPQt0Qqlo1FZKiv9xlfxlEmuwU5LN8SU
OgddWFV+tjMrW/5N+27TNSYNXGDWwC8KShgCUoFoJdO3Msl4USMwneUkWFZUSVo3
0enVAtLt2hAKRyf85TQ86CwpoXKf9j4f+k/tjIT0aHH5dYF2nEPQefa4nXSFjefr
cWCZFY1FbNLhLltZGWnqYW76mspksW3JodNhSa11W3/6aDk4C+IuF5T1rx34AJ5q
Ds/5qsCChJZfAgAusDZqi0f/KEDo+AtOnt6EhKdT9Rz4ATgFEboMLQIJHZXARbZG
tkTRCtBzceC/6XRkJ9V3mZYjrLA5u2gy4NNvlm+Xp8TPYx697ooM4IEwQ+JNmayb
hqzQ94JMSq2bWbAt47uSbSAg/kyHH2tNDx6KjXDipO+rUuPphUTslsBaOWxR8JzP
BbnHHmMNCH0apnCaa9/TS2KDPtW2lSLavdNModMI0/oWqoDM71z7ljFbu2Mg7Ak3
cuSVVd7AHN9k750CEYr45OUyVSplle1Fy44XzMsJVQcNS+f9UzpI5PE6zE06xRYj
E/7EQ4f/KwfNBw0Ifu9trsk4cC7XxROeCZw1IomsX606W4fXbYfJ137xjjSM+Mb8
PsxvXp4RjNszXUSA6sXatYrkqdChjaOdtQXsSh5PQ88WKxEHimv4VHxL8PiZVaJH
lbqRNzHqYYZ9VxciLSPwZV2ZKAdpFeSS6zIHHO7sWBS60qF5y06xTIpKM4tHt0qy
M1uiVUBi9/XvbhM2OzZys9XjURaEVnrzuGCmVlf9WG/CKVgzMZjmc+bJHO0PB1Fq
f6vvxdh8xYJu4fPPo0nBs4uozSrZRC/Moqk6rbhbZSS/JHL/glUGq8OkYTLMbfnD
LQfz+FVNkUuNd0svLOYfCCU1ben6xaCKkae/pcpQqZSahJMPV9iM6B2abj080L8+
c/Q1KYwB6KEox3MJlZA+ZWizJpp4ShE25z6G2ZokLpgIwjxROynLVPjwoEj7nCIU
9w3ovWBnQ9jauC7XwdLf49FH9Qmfd0IN2DudyZJ4vlw6dYI/p6UB1NSFWbTW2SLA
Ef4odmB10/bhJXc5pHqgLVxCQauYlpACe0FoICKMGqk8gyoT392s1Lu8bNixnzY0
04wUYe9twosFsZYPDeyNu3wzRn8+1GAZurh6WG1brx/JO2DcG+lMAauJMMGBKCjI
eXwGlSDoX9XFgJ4ggNJGaBZD000Ry9negHFmW46rF1Q5qtaA2Wh5h6FAw6oQtgu6
GJBTXC7KGndwTCnU8UE4mtgDfFevEnUD+8e7KraNuxKmgr2KR23q/zBt87qyRIEI
aYwwNbn7esZlRf20w/+XS/rdRvq2Kkr+V+l0O9O7uv4TQJuvejUji4nUqTgShIJN
mXpJtWcUHUkEqYiDcAVQADnTZza0kCnJZxvdImfSeyO3Bao/F7p6X3r2HNxD3elz
WWGbjwSZmTF8NBPnlesAZgre10k4x7w4WCccLyij5MI4Bqo5ifm01oJmCKtjun4L
okgJz/j7ba2bqewXw0fC6j4hsb1G/uDwBFiR7jce2q2S1jMppwciN77X/2CMJiaP
iE8Xzlndd2K0hx52cLSkc9oeHwiXyP/9XNWiObLUghxprWHTzPYD7Wy0I21YFYnJ
JNuMsz1MI5zm/EGqFczR1lX9Snt6Uta82oCBReZE/vEWyNAmaO99H+YDZCuR6yNs
WhFWKZ7bZ8WAvvI31oNlw/shFSL1DZsHRRNe5M69EcCFGoVt/TDN+SlFmZ9E0L6j
fvmF64JZ/BgVpyORPhBEz9I3mwbU8Xw+TlKURf4jAa6jQG/AbSAylTDLIB4E5osE
8BtYKWG9fO0YDaCSLPnYlStyTr5m4fo/CtNwFbe/TgUMZThbogDMc2PRIqMtAQam
b+/ObyIpaEM/NHEB9SRDtyuzXw6A56oqcN0IHeEWtMgwEQMCuBmnOkqTvwQs8GlU
7Mi4uyRXhn0k09E6l336nHfpyEuGsXjc8OG1aic0QFIg11vaD4tAAJ8EyZMMpwNt
6RAcNj5gtHqRrlrfUgC9Lh4swPaZkEWhTJFfHtL910WsJVfEdnmUD0hw1Gbqb+8y
QIQTB12CIiFDN5RekkqQ6FdSd1UiyJz9GC3EcMd1dxr07pFd0ZvsGK604HWYty99
qeOJ75DVOuC/BrpNuxc+ZsVzd2zWeJKx6Hh6i1XVxnVpOOv+YE6q2HLdQlji6jxy
z2jJaaUSYgqVROstgT6X5yXGPWlT2PCvy38Bz2oOs0L9Iv/mgM107G/oslxHlM35
gyKjeReiZsqzucaEv4jMapAo2u/mQN/fXC0tr3R/cvx8Qkf6V/PwZrEQfpf1cwGT
Pkq1NBeNlZv+qUKiA2tTwL75bZn/gAimbIBzsYRYaaWjCG6AlhYrkIhyBJ/6pHuP
f3o78XJz6mJ/8E/IgRBZomzz2FTDpSJ3gfHq7gBAgUU7oCZbyiAJOUFKYplGUUxv
pDtTvUCXH7CxkYHfd5NWSxiK4ij8uBPak40eTCHme+kP1vNLDK8YWLdaSr1651lI
T+70haKyq0s0dTybJ4LILMKQZ0FNMcgDL9vz4XCfClsJJ7nZSYhdBfDRqYhGIkJM
qQvuH4I6nshZaUQM3nQzhCAQ3v+dyoLvQk4M+SeztH8y9mFxvU62IOWofIIwiCo7
CIRf0DZwMZeJgsrLVqHkV72F9Y6dMTpxmKlXEz/twLFqNZxqDGHGcCaHc8lG1nzJ
AZSeLdtXZNodOG9xq7c/aHuUNUKHR7FIyaa69csmn0fYTODi4+3LLQH1OyoOvPmT
nJ3vZeH9gPw72sko7Huivo1XPeVXZrGc6Ubyar/4YgNoGU9ksoolOJUX6hGcm4U1
HOV2H4dJmOtMFXQgnC0RMHzEqxfL2ZvpBeSJzVZx5uNdzmXl5WNfxck4nVbSa1NB
7hQyGh7W7nJHhw9DYRrDXZMauK0KFVBThqgtPKjKgcbyuBUzWuJTupfwiey2GAor
XO/YRShdQZXMbXrr9DWK3GC/94daQ/a2jJrgCx5LQAtqArcbZ6p7OEtwtgGu2V82
Mg/J1ZO74ssFhCAsBdntiY3DIz/IZX2QCtXCm8omouuEJC3LKJGB6M1giIdqcdIo
Fa+NA17sxJ3P4WoZWcVThlI1EzZ0MvU28pTL9uVdMbQbiymS41Syosjr/l3qfqRc
Z2jAM5CO+zThBKtqDxMLAFPQcs9cpzmg0di8NU80XflxsA7CLtuOebOpl8aX4vNd
Q8Cq108ZGo0tdt7MrskgVcqx+KoP6v72CQQ0n00TNuJyyqpK7yMB6Jc482skBl8g
u7cCmxS9fYlta3t0L5ya5NoOX8Eg1QKNs6vNMW/qqn1jJuDlrTFKkc4Nwkbi85WS
zdXlO219XangkVpBLEcG9UIliiX0rRVDrmte/W5otlBn3RwmyM/UlxYH3tzaCsx+
zpmjeQqmBMM5KrccBVw+qIDC3J1g2zXpltWAvn7rRz5oyZjWxqQ61VQPIshMZHJ1
kFVS51lZosNhAv1x5gM9UXkgL67OFFKRG4zuOvFcFaJmW2EpS84DhqqJctKBvO7r
qwkce+l1Xdlyk/SSMB2gJpi5j6dA6m3ygFyi8yDkWIJP70UTaCUuk9JZYssCizxZ
3j0sIh5nltIIEIVL7loOs4hHucqUBsEoEa76ZorKbjh8SojD/Fz+0Q3luxaDhc6s
2ecmr6/VHRYvpu0WuPaFmPN0XR3WVc5iUOQ/u9D5BxWGHw1FL213U6/t9+2CxYpf
lyG42eKEkFsfGvNMRfANde4g8fgMizXjYr/vMU+uVVPg0kTdFstA+ecthTMavS3q
reUfZdhPXIKCzvisY7ChBjmQrZ++E5WgA51u2POMkVTI3kFThHgACQLZ3sLTekOh
fzynQurYVKZS/79tqdoALkxDmXu/HMoz5FEphrx9NKJ4pSmY8B6M/Bzd4JH3opS8
WInKBGZppHU3xxF8/A7AfYnbnG7BXvSPVveXvC2sGfzSUNUitkRe1EA8apmfAQFS
9cLrnpgIiJ6r89FCqX/3Dz1rOh2O5DdJEgpgfm22rBlAvIAmZhXo3awZAS5StbbW
aG1cJ/bT+T9GxUZFJxOrmseicYNN5vqMtmZMOJEqhVJabtuflIPvt2SLQdrPRLRV
UXtMJ+6mBYYnoAlSDXO5RLL4uCkL3HoKVGi2RNUkhLTX13OLcIi+cfc8+RwioaPC
4Y5KmfZgatlV6Yv5ZPdnRmC7fSzWSQuo6M8TZvgYFMYGffv8BptMpm3ZDAFq4TDs
jWIrssgcxhQVhHzi3WXQz1/HXPIkQSczcgEXE51EGbYE/0f6d7LIFvzaubYM9Ii6
Rf7WMkfe0yJs1DWalcdH/xQuRWvbxtPi6414kspYwgkZogbcOR49xsJERox+7hoS
BSblYMVnTss1TxKMHwsWNhZIBWGnmlEJi7DEy6F4+6brFezN6Mv5bNNl//TWf9X8
fVnS06M9bL0n5SRV2mIRmsNx65nREheXko0tqWWEycrX9nEibwMb4A8QH3JWN++8
Pobi/wNxzHJNF2FCVvFlezVkVE841Ohkajysi0LAQMZ69r0K3/OD7Qbo3inOm+pe
0gPbOIL5NkaE8aN34Y2x32H7hB9axMxxw5c5KBfi9RRb6IH3l7Zx2TSIqAUtxSEJ
XpASWosH5YZtaM65GG+7LAYRIAZR5fYlc8BPS/uneOwu0qleR5cU8kQ2xvA7dyM7
j2IDV0zIuSys6RTBM5PF/t9+YVsQoOaPNDWBBI6zbBBkYYGb2Epzyd8J+mjqfxyt
9pOgnqf6WIRQkNmCOcyDu6OjdRZg3PURUKoyBo7+c3IIbAPq7GtbVPSc10EhSRnH
OiJNlCNYBoheitTGCd9RaKroyl0caWXEX3Dop+Hk04Jn3HqXmrgG1MOXyXa/YmJp
yDcAnjSIl9f/eAHAONK8Ypdq1XtqDiV4o8MoQgzRqIRPFQ/4X4pcEGt1wMXPORrU
erqUFETAiV4aXt42Cbq7x1J8xlrONRiTNDDWUFYZfZiM3Lmj0lmMk/aC9CDteFsO
JE6k+4EBgzv+bnu6gMU3AgG/lxbjkoxe7u+cNv8ZL0Yh9jYkNFmzVHI1qQWOwUbd
tGjCoAJM7y9nhIDgLw3oB/P9mJoUgHEinT5dcruVdbPDzrmI1th35XdUK7wFC4Bt
WoEcoCPART/tRu9zZwd6r43Usy/jIWRI4DHrYndt1zg8NneCas9lfvsgbHfkDoCB
LkV5V9M0fpfoWyfrNrEXVO23rM+YgXHRy+cyRQryIBSAsP+xqKmpLBrE1Nch7hmA
DunVMbI6AwT/GK0ggLXLJYdqKSXf+em8pvwprjBczhOFs1bPLKUHULpWm2hTd8Vg
PYVY00KXArzCrOCL9T5eisfRm04NdJvprxsu37F/hMMuUqHM4R0zzdvu5pqkyve0
4aA4T9TY0Ixl0SWh7WYkO6kdrnusGbZLZgjCZQUiaa2QE4lPyKjtYONVlDnPGamr
+1D6wy7076a7GyJXjTOIdNtIqAJuaFM4zBjG+f8JNufAMIzFH4/a8PxnpLPr8yyN
rU7YLnHRFabqWHddzfe6UYXz/ntNhYKXBAaKih1NLYSe21SHRSSMR+6zZDS5MfaQ
+ZLRNLgQXmj0ygzxQWLMnygVcNHyY+NzyHaZxcENWP9aNVK/oI0L0hhmv9G1d4dB
gJIUCTOJpRpRehfM/XeZle1VFM3URcwzVXI0Of1deJKxE56fL56jt3DST8i74hcT
smApnQLxe9MlG7jbpccDuXBJkFsU1b7hocyVepyXeL2HIRXbTPXh3HgGVuW8f4eK
AXxqeHAyCR/s5m3jQkSe1lXIVBvBr1+NaH0hBeJdxELDJ0ogVArYH1UascRj1MIk
XZDJyK/5Ho4gxGvXfJWBUvDqBDSpioUQglfsFZc2Jz/OxMELfcDhhueXW9H6fe5z
0RgPEuzq2+AFLvM3zjgyMsaJasHzMRQxWwmpncmHc2b49l5510WR07uF8xBYNQHL
3kbzRm+mVLRHDGLSFvHcTt98CCDa/HnEe/a/tNZfrIf6u0BIMRypiGdp1eVZfo5d
fuxu3PPr+WLASB8V7R9lB1rY/ASE1/VMo1DvuQp+gW2nd0e5OXujdt+vKbXZqFoy
gLGFvd9x44AjEv+e2fgIf1rSXxwPxilLtNp7SK7ThTut2MQhgcET/wx5dI3yi9DH
fYJmQDaSRlWH56lLnnI5gNPmdh00aXjxz/5QrftjoifEDn0B1ovV9iFc+aXeFtF2
rUK5MfG0M3QTTOGMrMx0MBeeP5p8jvxcNqTe8YZUYF8tJhpkpCCGC/+HwU6khM47
iFrbki7xKEnaULD32Pi3p1GG6lcKIL9zfYZX0YLdgDRoJcNtSEchuth6s9jQDoXG
HCtsZjwBWj9m63ENiP3Dff0X5xLkepUlfV5o8BZBkjZb9MQDkD9Ohrby73dF79py
J9Rb/76BovNGthm7IGcY3hNQNG3mtresDnFdFsDs564ITblFRbDK0GVhkchot0XF
xcXuNeoW6xOQtb9MwKDP46UrbM04wGhdDoWnOT4Zwd5hHmelMzOkW98pxo7uxeGS
neq+ey6dteA01LMESS7QvLaW5G0xJq78pacxccwUjtlaJ5TOuhmS5190tngsiFsJ
DYEOrg2UH64ixioX/gDQi+7mKdbHjQCO5L49lg4DptKiJfh781MfbquzEWGJ0opP
VYARKQvm+AdivnCsiuOrs+zyvfM+nEDW6rVB1GXYuQ61FMyWlZP0vGldpJM2dz/t
XHV9LCnfJMAP8Xz1qduAxB4+TiW9FkYfv4HnL2si5Y0cY4FRmroKwv1CQqxcOYoP
lYltgs+37BuFVQoQNQjqrJIFQKsQ+82dvROU+9pQ+h2iY7+pT3W0e6kXJYFWt5+R
BPGVeunHlgDQp33MOsYvyQ2UjM3oJjujLik1Zu9urmD1e0mESckf99ipfrxc4vX3
f14wQiUk7mVRa1fm9ns48yVEmF0BHmXsSsvbk6biWCE+CwoqjzZ3ICLq81XemCVe
z8fE+hVSH2bMAMqIoU+4PAX7Y49Q00nIWHuSm/1k3QUqBoe/tD2okOXOI57jlA9/
TtrGOrSV0timCVC3drKrQPb18Xn6YWD5bkNGJ95Iw6NG+dpgLzG9PG1RYcGSfVIm
2AlycXKV6XO2H92F5Fjal7OSVHmA9fjVH2/gTJc5O76cAsD3uBtmWxFdBZTb6mim
Qvt2huPeBZty614FuI4dy5k18Z+8oXYS0CcUngWOjoBQr2evuqPW47XTPnCIegAz
mgQAP2dGQmql1KRbryZiR6r6kF782UHLIfLDXeQrGcNSB8Pf7pGya8oalzfNv8hG
sZTQbeuP5JkZoQ55mw4k93PssTCmH0Q0+bpILu8+vhW1TtPNaUL/Jm3DYpnYIXiQ
6sCXIPKQfUDfabSy6+EMNS0qLa6bnfOXXd8ko0U9UM66NkFttZGzKMfjUfjW3lCg
LVoAb5q7uwY+qrE8G3a65VKoumfzfw/NxxMy+s37ipumekaSV8Ia6sv29anjlnEs
AiHpIMSKOT/oAHkAuCcuZBSZ1ch7BVY/mPN1qI2+srGw0u1678sPLKclGFprCSUN
s+L1y2/I2UQlRTuV8TVTfGqS32cCKfaznByFu7GovP5cowsnSKpTolxHHsgRZFcr
qyP8z2HVR07/Jqog2a68W+JTKaaiLhTtfOTNkyp97AfXQTXtDtNGhX2KCYwFLtRl
PFrbQS2Gj4zunPLrOg5G4mL8dbMnIXP9rAOcxAs+VdlNvDq5VMkh8n52S9MhyDCq
1AlaeVu24XB262SQ7AoiVo3Orvi0Z7XqKYJ6ZJMnv98riTgD1yMFScOFnjh2KOgk
0sJssfHNHtoBXzOCSYUU8zuWAupc7+fAn3pP5BR5+XV9wv0f2Ej+dI4k0tIP9P5g
lPe8c8tfpVEsaLe5EPWD1y8AFLb2sZ5VphzMoFGdRn2sH8RZZQ0vaZhkVAo+VKLM
Dn/0g1NrOff5a6rdAjxJN6NsqfAjFAEP9g+aBX8PTm9pZ+PO8yh6XgaSOTSV2608
AGnNqGRPGtesQ1x3Q+iamKJ7dsOOt8wmxQXg/C1ssqlxiYS/+aP0J8bfOXBS1JJ3
Wrwy9Xv3TqWR/I7PEPFd+OBdom01Ppgw6GKWT2pZAUYjPqwXDkEOIWDxZYoQ4F8v
p6YKF1jmnI+vyZ68HCWt+MBW15VJdL4LW5PBnvnyFkNwNsMfT+HWloUdqEIDrvxI
rMopNIsUvpXoUbspDRsEtR7WkOFqqgaHqm6gTr1et2Oe1US71AK4fe+iZtzGAlCD
jJAKj8MtWPiNh6/nQ3rUow1KNHSMHkCwWa1PqX0luwbZ31N35FUITY1gxkPi3ZpI
TVOnHDk+9/sRC2k4QiClVVMtHE0JoxIfy4pZEyb8Fe5FG6bXc/H53l0Ty3qhm+J/
9vzvJutnW1KzZR0QjX6WQYODkCEoYtFkQN0zrr1N2L/DOghkicrYFi2hbr1BRp0Y
t8UyU+0W7xmvT0qO6esiLfIJ22J/tZ2sPkS9WrOUySSihIZuc9durWGUSg1tstIJ
vtcA7l4vdl6JZVg77C653aXEhpVwjQyLiLEabLl+Hqo8ucbsJUX0s9JhVAN1q3RD
3mKEGAu8OIw7Z9/6kM0nwrwKd9BNUXOIzuwO3ei35nPu5wMDAvkpXGZ9Ppb0iZSG
olkEbUChZCRSufkpiosHu+JdUtza9wGjsbz+X32coDqYGHzuhaz4J0ln8dWqPg+J
z7YsC93vTxdFUH7Z+alkSIlIzz7BxhhUzuUuJyI4hJ/S0J1/gV14gWMZpR592khk
hIJmcuIGtnl3N9uhZamTyA+hPUNgjg3iYyDhNPN1H+jzA0jln4b1NwmO/OiJqZRS
tXJf8GlLM4j0GCumNHZxta2qnmL7e2c5eAfziVYh9S7LEFljNV5NboyZrB8jL1IC
EIaB4vICFh1t3InNUrX0m49Yyr7xmhK6hEIRdsRCcGjcEL8Nj/E3bSG7B7wH8RqH
sZ9IjY1ck10qZzkl1oOCBBO2GC+8Crl+XgujXunRzsptM84+ERF1QMXJuGiF2lJv
Bv/7xuspndEoxLt8BsuDPRxc8jWbz3sBbF3fqySC1sXRSKIHbnQvGMn4pEpcsxgP
MUQRaA7LEcXxXpU5RvtKKG0TrpMYmdY9EM97Q9bN7EUCpXGNwUxxhprqCyTYbrtu
7BZ+cMYyOCbDCpvbp/cJKn+uT8JPpnNa+mtuRtM6xeq4e5QZ0mdIDXOfCR0H334g
Mpp14rIQoFmcZ6Ci4FkvCo7WUZCbp05IGcLLp91A27hqzMSfTrf+9yr1ndSovv/w
dj4C+UD03aHa0ZXgKanCeL5QXqNz9db20VHJdwPhxvhYDpGMU7y0ZRvMyDYOI91F
hh2xrLIRsL64Ic+BDi8YLuyS81Yoph9gy7LtPbXI/6Eu3sppLffGF1wePwTa39cy
ZHSX5A9Zcouy6/bWsoEazlvqSb32gBVeX13rslMkLHUmRVBYP/JZETnIcerdD0vl
bxaUMsN2mwDPdIxVi/7PfXpdZR7THQ2QxG3uZ7gQP/wuI/+bOenVqSR+bL1OuK2U
n+Qm1KNe/1Gd+p7hfAIAQWEYfDmBz+rWN0amIzIFtVvQEMjAphgj1/kq7nusEEbx
r3uhOQIrnN0VtZ8ebVdMp0nRasH5TLmGOc1tHFRVFmSvNFbcjgBqrC/YQfZAB2IF
sP/4UT968vVWoTBlvoUHi857uZa/IyzesfMNVWbYfdBGqWMLofm7oEHRS1qtPZ90
XM9I+NR0woRhwQL+ykqm7mAM3pTJp3Ai6TnQyAAk+cUhZekOl+hwOsw8CiZyvlgJ
ksqRXzGVEnnNiIbfKiEnKNTYgTdJf+XDTkJvWbVRv4FcMumJoXJcNmmTs69p2r6f
68kqfqBttT8xyWSm6AdRhbY5F1zZ6QVKtANeujMXDVD8WFBg/6NWH+spYWe9hNg3
bTdN5w2SMf8trmmdG/AUHNNY/LwCijHfDtO95DTND0Q+9AyukN4SAD2rtmpYdXJN
0CP0c/w9p1jONQmAA3uhSv0M8kPkoBDApdydm0JPqO+klSVDzmgTTwPbewiDuCq0
AhmKmCmFfunH0NAYLdHM5/sZzAAtNxDtq2bIv2fJ6179mBG7dguSa/sDdGK3W5yj
DaRwcBiagI4+TuHnSgcNl4Ryy05dddlLULdu+I6F5hkEA3e6qdFgbA4r0y89HGGO
xdYIyd5Pj28noTYUfgPq+fmnlSAF58/WJtwmdpvP7lArqIJAMXHaz2z8Bo18gq9Y
ZGbbrM1WyH8s3cHqiZ2jfLGGtRusLqovejWRuQXVVUhtigfRkjeNnFBi4HFLFZCT
pmMJhA/UDjYF652a0GNW0dQaPUnUnmLCnr1MN/7q7HjfP7iIaPd+htqf9QKgsg1T
+rgpVYqAhVb/9BZv5rqF2fBfGHw9RbOIjwxU8iqZPW/v/OipicNd9kOWPFFo/E8x
jaIRY8D/4Cke88SxU1P6pjGU0lp4vdSQ8nlA8jyUKk+nUgJE9teVyVHeCFFck6D3
VV7o29U1UK0wdI8mBt7CvokpMMNywzp+eSwWAOTsA6fuYzU0HMhQ54LV72J8NXx8
NqwxYqTlHuvEGlzJOm/akqDPEQVzhihnQN0xEp7pjy8VncblMe0sft2PE0VW75tC
1tCHxyzZwSgvV0/NctV8Z9zPy3KhdoZqJs18VzCic1ezb4wCbQjTH0NskcgyveHH
7LvTAyTmnikbXqYhjlBX9IihBKTNRPf7B7U1cW7eXe1cdxKwqJoH2PDsAY/zObBD
GJDIvKI6fNucWiLuSU9ywPqHVMCrX3SZBxiAEjl7eLBg5pGNXHjQ7IGxHIyFYWd6
qcmjC+/+zFaFw+EOE9LvPN9jUGWnNwadTsgDw5iJV+m6yOM8mwt+DZDCFDLIcV9w
nwaU+QjngBqnVoejqqddYZZzgp6PrvhS+DnEyNtwcg6ZCjfX5dHjDwS1FOcAU+xC
jubqbBADZnsV4NIqnEB0KuvsdFwxZ3U9k5SYkHjx2dVlhaahkZgVIAju6dOU2l0R
HV711cOvdltc2I/Ed70HSxft6Yxvsv8I4wiYtlguQdFSkYWJ/65g8ECXjH24Gxfu
b5UChvn8YhAtIlB4fSHZKQcfqX0Ix/Gu7UEs+oIFCv68O/5lMiEvUWxDkryY0MS0
YLzDWVWQ29wlymhblnzr//5kQULPHjr0WIU/UoU1d7jT+9ApFlaPno+jvCtoh6tc
lEjWenZeObLg4qgEwZXoR6LIQ3ImLRu3eDn/VdEwoXqpAgmmXIKqpsMktpry6iiB
ptYT/J/+J+kmDKCDx4ekk12IIF/w60EQ8fR7YFFdsqfXMna3r6pXhZDbWZIMNB+5
RsrlNyGMF5VHUZgOcFCJgmaQKflL7QJwDN5pzwJ1WBLJ1UsiyVDcfw6etGdEfOcH
rD5S47TuatlWcF/pkOJLlSDroGvNFN545sXqXaC6i+dano22XtwPcVf28UuF5T48
L0v9chDbXsb5NW1OVDPcwWjjlGCaBx2ymCA7/awWDg9DPKjmfRqWUmmQdJWyGGfH
Dp53lo4EoSaHvXHeeq5mZ2hde1SGcagf7ATUxB7gSLYQpAEAnfo66sW/QyQHioii
o0cDUNIZfdllzopKp7b8dpTbjUiptXF6CLLID5zGqfFubmoQE3wrMMMTAOCwADSi
Iu6bEVWUYZiPhKM4mqfN5s7pa8vdJcSibXBziyO4v2jEhca6TCx+ms8pLQfppImm
3381Xblgc/IDRwx4AYEXUOOKMDfCV9+XyKJsh9B5Y6WoULB2DMz6SRBZ1rZTmEza
0FJhgeRQi8SBh8R4exFS52r4kyF4KFqFDA5VdPLEOD/ohmk7/Cbd4r/5OpyfkEQV
jeUNcnoj+oxAjzYnXmfLrqc8tY36jlcWL5IJtin8XZFtvajh8mBIsubwWeUawnjj
cTl5buUUxclFnOLpoYmm9IUvMPcyBz7Q+XXo0RBq3WNFiJDDCa7SfvypiWxP6g+d
pecoiAMp4VTwap+IbwaugXo3oIlCZDzAdGZQyLA0yoXtgZrewJvkUhxv2Q5xvAg6
IUQnq+JkpDk8r1DH7Gk0WNL8bvSTA1cN8Jg1MxdYYFNLb756wgAD553crmipsERD
E5olvG+fBoVIvBJ7jF7yRhXhcStfOMqub5NDuOHhDe8sbWlh0T8ip/KzAiNWqux/
6wwAWQ/ztFtuRAgjXVF1kv7avDSx2uiDFz1ryUuKHKyObTwgNGQ+RicFOjKpKDys
pLlDDrJMtjb8h5OnlhILKottuRAbOihRQHRUtBGfBEiLMrn/OkVlWMwTdCVvw3Sf
+73gZZIKopwDzuMmg6WT8amy9ZPzrndW2TIgfS/qdfqKsJnugxj4m2a1axYS2Cpg
/Eoe8wIj40ztQ8CVdTusYLLueDedf7X4XRR/BXx0QUNausK19+Ln+1+E+ooMXghK
dFV25d0wFYHwz1rpDwaupLobmrUEmAbsXE2pIq1JJP4+BvZBII9A5ak5+8k37H9D
ebTZYlJuzlja9aPpiSpyDT7KX+T5XCAYIPDeS3VN1uNbIEV+ueF3H/u6Mgcxnlj2
BQVlDWbkjE6ga9obBgEVyNCfvwM8W+oXR0AezklvSnwF3LCgCKddY0DjfiYVZeXV
5RXh+cLdzpZ065MFBDgUeRjC4ANROhItCraWfvbCZ8fLbE8Vzw3FKDAPU4KRtTzy
ydI6DmcHiJyv2UTkOwyN+4jKViTZjbcXYO2VGvqB/+ZURhzPPG3cB90CAg5tOaSp
B3wcwERrpv5zBYVydA3sqq7a6kvkNTsPVymL18e515Tc7uoLLLksSP77xx8SY0Wr
HOdoPyF3ELYtuG7xQ8waxG/j91d+KN7nX50TDhjiBYGzG0+buNMGAIayvQvKQaKn
vV3hTvSAu61lEzSkIvif7A6bH/6W+tbqAEOlVbxkNPBvJZfUtLse1LA6gCmd3RDm
a4KudhA0uAem+iAwy9qz1D0VIGE1WWPDraQ+6koL+OcI5oy2nxDMXCF26FjuP5Pi
IJbX3An+afdRI8ls9QaROWs/Zbzq/HYX3aW2fYBiM2AQjbHySVPteEYisWOr4dxL
rUuPD77w6loLZdJYK8fyvLejnPdbXeYeKEZTJC+MBcIdAQqloDKuMsncLskEdvGZ
U0lzfwRS4wwsLpBoUkn9v3bXibMSMiTUi5PGaLTYiEp9tRzens60rF315fYap15F
G4RW5X4cMPNiGuKWSj4BfaUOTsky4vjdzIAkEXwpMbDAK3nW8CKU+E0cH99nuvDK
RSqoToPAXyd9tEZVNykaHxGpE+6BZorYMZ7/v2EjCjoIDFbb3395RsBCOLOfjpaF
PLoetDw/vypnC5oP1B6VbWvBT/6xdoJgGQjDR5zJiZtj1OI5nrgnIh2w97suy8H4
vQ4ZYBjyw9Ch1W5x12Gjd5eGkO8iHfz3G0sarxfsZDWPXhWnmrarUP3zJxFaADSr
1CTzbM0kTfZdKuP4IRHqOpS0QEa1t3NFHD+ZNfQbHtB7tJ68FgeqqCQ84XVCMVQO
J26ECCV7MKdgOE8VzmsFGlwCTg0IbKliueNKoYI2xRQKAPpOWzNnTXfUXb6G1+F5
0yfCASVx2/aoJBV7SA6LWzDivtHpaOSi270jaDIetjzT7Y0xelQsO4/jLkAYTk/w
5+AXcX8loqvXT3WE319ZRZV3sYVVknEL20QoF4YEpUUkO7AThIy1AcR9xg/e+nE8
u7tIt9r6YzEiOaegVqA87H7UKtQxu75XPEsjE3w9G/9zBb2fywPfCb0b59Xc28TN
IcpmgJxN28s/7rDiuL+kU13oXX6N27JvX4W7ejAbOWZIamD0r63qtZ4QAhjnC7oc
mED1Y4FT/qLF1Q1LVIP0tc3hcxYsGpyU4kx4rCg2W4BF/oCxvxhJauh2KhB6+usF
T2Ze6bLXMuhhQ5n5G3vD1HtzqS2xcMpYGM2ls6ARXVkOwEZzERkf5Kq++hh9Cmhl
7gatqy0tPVtZfEfjWs8dKa2PR/9tv7kEzWMmB1SRe3udBRQbAyOMHn3o6skEEyxF
BPhPZ7ts2Qzb3frpa4vkOiyv4Z2cd+pD4+EpnDqavSj+vndSUMpWzsv1DokPZQ3C
2JgcpIwB+CvHjsPzptN5rHbE5oTdbv49nlhCxuPg9uRVZxaTU1Z/KlGWLGXQ7wob
iXuBQeruGmRHSkMdOE2wEz422zdyQ2ncYWMGc9Hfem1e7kAs8fgnuxNDf4DZODOY
rp7rPV66SsqaG3z8G+Stb8xqQ0y+fZQWSZXQ0Y9tqN5OK4K894gL1zFWpEh/NVWg
jmu1CJsVW+dlvg925PblCV4Lh87kpM+ZpyZjUEiaK0rlOuZeR9Enes3ZNQv4pQ3n
Kw2H2GUtqYJg8zD0LQ3i4VxL0ONWjR28omAWC/cioDFFH6Ovg8QdlPdGLmcsvTXd
M01bDxWwqBFjAKSCG9yImpjsd0IuZN8umQBa5pKdrMVT/6TGsYR8tAmfnBEprWF0
ynuxcfK5OdLS3Wz1GzhuL7d/fwnlauxFx6/tFLwxn19qeZXb+cs8eMC8GbecnSIv
kVi4ddQSVFdPBu0bWfVapv1k4llmqZ8ECKwwRIWvFYli7r5XSu9ifnWlCMpBsVCP
lswLxteFY2z2VIhcwGJIdITJnpy0eb0yVWZvDr+DBUkfvDEHOmL2rYUH9AxevBSE
spoITUW5h0VvrJqAgNqwnyPthH3hIuldJMHq+bZO6/FiqRRsi8Sp1S3GDWVHfSsh
KhRM5vI9BV96VquS/Yg7wX3bI4vv5Ok8ccnv3by+moCxL0mW3/gjlNqNNCVFi/ld
zUt5YVgDvp8TCccWdRbi+h9wpnzLev7CheujeZ9Esi8FrkE5uWGTIcQunrZUUxrM
gqtYvAWyIDmXrPJCJTa8zFQYatp8oFdtR+YfTFR5TNPuG361pJFjCNjrR6UmjWlc
nefRBiSAbp76DHSpac7TVe6DR7p9T/r3FR2fHuyq3va2OKsOjQSyKf8FIQkOzNLD
FhyUQ9wZiszole4mX3lqyg/DtFdvZnhqlUN4zqDcaaHomXu3w0nDB7ygqzj3wV3q
JlWFjTuPYwlDXGCzPm/YO8kIUIXNdcUICtbPyrZNZ2VdvDrzmAw87m5X0I4igWJH
LJ27eSBfu9GCYYFVwpgCAajVeg7dvMRTV4RUidVRvDLCjj8RQGYixL/EfZS6GL4E
v0KRshgWdCkclqXIlyt0aIg5imKOOWVTCFHbsMO+p2onyCfgv1g4BCgjPDIce/+g
ljNzPAnkRHEVnnv1ifcd30hpSq5hz0y6yIbP0GzWKs/PVMAPAXKdnzr9jUAZWsDj
4QYwlsp2HPzzsK6o0DSY7vPel/YuCyPQ7xK9XSD/jFPLEUf49mv0d6pDPSACvJdu
MoLbPxQsm/2ySrDOYX41tiHIvUcjLr0eilDFFesV2rj89d5Tgmhtc+96H7Hikgfa
oogY/xbVex06qb7AFn+WDFG77SwDYDTAiMPaLz2JdeDLGfp+GMjvBvF7Zo9OOtR5
iog2GFwmOeNl8s9NRSKyxGUJh3lB9/xnrfyrb9HMS3CQO1LxtwIloWjlHa+jvz/Y
qjwCC8B/Cp1w7rncfepqv3MPJhUZoWMoNoE9ckK7iK2j8Us+zHN+Ffw13AhvW55a
q+Pl2dHFLY4SeDinE7flaRt3KAhMs+RGIuHm4msvvlJuhcfeRbx7j8UHzYdALl2S
1PyPo0zX+AmeBp20vsJ+X9zt1rn3+3T1KAGyHVzPBjGEuXNUppJfaaDsRDhdd815
IBOZNwA0DbN1jxUOKTcxcjYHRwpgVdY4Cm3e/AzWAQRv8Yo+jZwBySnvqjWX8P8V
m8x1ILqbQ5/PFn9obpFRZ7BMyegKFCuj881veAfPIv95aduw7N0bPFr55xaEhzVT
Ax+Mio8o6ce3b4mVOERBJMDKgzx0XHkJoGqFce7xQ/e/71JErv4QcBNA6+duL+PH
XQKq6YbDFepqN5UwwPKJAhN3Fkpb283lhGaRYW/3UsxZemMOxjn68CKGw2eg+2gq
p0su4G3VO5tch4TB9NIEM3BPb937gdriWXR1O3fu95mRi4Qp/e8YNiyeasCUH1WM
Y4RRmeHXnu0I42JZPVJHdC+V8LsvBUJi8Lg1yqainaXDGNIE1ZxNiguVdd8EafVy
dKSdFVqsFnsL+M1XUtXLy6Izo3wduhujeuvzVjRdBeynvwioZ81xAnIN1cYM4yyL
c8TJUWM9atYReXNPH+VnD+zoSUotggSqxjnUQ04JZj9LW/buM1lTnY5b5rY0v57+
nibYhqUXT+qwvtD6jZZIVTt/TSNvrIqm/JXT1OX+baeYQPQwlIGTJYFq/weEvro+
hr9io47euHWlJ25DTZK+OglTmgrZcLqpwBl/YHDp/pbv5K2P2BGHUPEMyC6cpznA
r0xha5Grd0PUkMJaDig0JNDlAaqUG6B+cfpMD6cDGh/D/G5BAqk0geLniEqeqz+V
MXcnmdwZclHVSyl0IgFfQw/f0mHgzHaJhDMgnF3eO43xN+7NleuUK5uigjCAY+sS
kQgwa2bgjKiLOUBKCDrKMjbtiFXYDepjdZevCksgaWW1/a5dwUqOMPZLOq/SJUsr
uaBz3/WHWSyWoqHblcqIeRmlc++QBVAYmBixRLNNIL08J8Sv830hkOBjZiJIm0wn
xNLRfgKtnkc9A+kC3ZDPZk/IG9BIFzNuNAmvISVEctZApXWqk9MS5rcf6iFVjYEj
nk+EpAm9E9rMsoURnaBGC+qxUbRcJ0DRavmhwqQFWUq2gmIrFl5E3760XUkZYuuP
gG6/NZfP3t3kmTFBE8/45JpKnoddOYiypDT+xMMjDkzDiXu5IACr/gNb9TQg2erF
A+m3HvPnQWpQ7lcqZiT5+jZSjdTXlR5iC8+RBuJZoaBclyEGDkkPxrtEBKrhlKqw
FdwJDPkzIzX8/2wttXtDkltuksWgB9Cu76FRvY6L46jaoLDla0V/dJc8b1RG7mFZ
/UUOOogkLWjcXEQ/xoS7OhxR6HbKlcKKSIfOMD1d7IttyFvzTFnEQjSJ+3hNJELU
iRoggy3PX9uKYY5sInNbZPGMycwhpdjV1a91q9CUPOh29xq/TTSuXGOzgvQ4Eniz
NxTk+tofgl6WIYU0bVADZ4eAW8Vfl/iDJSCic/T3Ac7D4Tclm2o16mTIx+d79Q7t
bhxSaU+JgfaG8pm90D2tY0HT+1lxeXrm8IsU3C+l37mvTjNeSb9VzPg3+K8fqldb
cSQi3rScvctmpNeAG1ulp0CUCNbYcnm9vod3zNhvz+0oSHXAdbZP2SPlqtOXlzKQ
q3W5OpgBw+FdkIx2GHB2iPLHeM/5jdscpBLB6SyMNoMjO+ip5oZuGn2c8uCGBw/A
Mjc7T6pTGek0gJeswr6BJg2pQHLNgApahz08xU/GiufUOLriP5OPv+1RtKz7JL1A
o/ZECBnNQC9lVvZrED47fR1KW/4+mxt7auTT6YBJRbZPArqIQfYm2/UY8HiRkGJQ
xo/XfmN025sDyVpd2SpnPdCTw2f/WvHvNP6eRUTEP0dmLV1oNVnVb8rhs5t8DBdM
4q81lVTZ1q6SWKkQeyGCXJgOgqdUY6Rwq2ScBE/VJTrbJyTByIRRnaPmaTTsv1KZ
LnkKkmsFd62jvg0QqUzig5vethmsxHrrFWWV9Q0MT5bj5W4cWh5/Qd4JumySFazv
IvreD4OIY536MdvI+8lB/1minUCQ1pyH5MB7muQqU6rs/tOuB9RyYg6iDGefIcfz
kUQOaJDSf+TZT/4FQXpMFnJp54ZGlaca6OBVv338wvZ9rrv08PHm6c5yax9Jc4iX
6IxxNQnFwuBcipHUHQORcoEwvkavROklcqWQjmpHJDhi+LXOCDOsb7TYpTsfVCtW
TMaApZ7Sj5ToYKe+1CIlGB12dx+N4Gv3EuG7stzgCnXmmGvEjV2r8fAnzVCjPVSF
GbRiUq5eaFqkiSo6p341MXmvO80R+kL3nirPbezJsneEq5oppTNG2c5OYFh9b3Zd
us8Srx9uibaVzL9hdeR6RL7wdo6Zv2ubdWmAMaDqi9nbKoZAlUgRjJ+FlsRdv+zO
CSBWeUyV1pVKDG+bT6NENQ+JH8aGDzuuifnEERcdWYEK3IBCo3pjshX54r4CwLko
dU43JBZU1AHtog11MsBn0OfGxVlo99ZovpaQfIdb2My8waKXYo/1sxgK61YfANba
fIi6Bi/p69M34MwSUNtn14nA8/gOP31O8NaqajCiqC42bQ6mNvRcbTSwvt1nky4N
9VFkxZOGq8ODBNHlugXbkUpmrHbLM2cq8s3+V1u13fENT5ZOyKb8PiNeIjlZwrvV
paAOq7sUjwfalQUQEDpbg88PFJeINdDWpeaXe2Fn5IKjs/GHgMJWStuV+JM6fkIt
MAvHthJ5JGSiWlap878kuh6UDzj+vbTJJvvG0TeBIs4kAmIRgbffbF3fGGIXSOZq
n3zChDY6k1HS7KimA6/suZO9eKdq38U5SgdTiP0MNJgzC/EFFEnCwt2FEjABDz9B
9t57ruMTMJhYJmODtVPlHU+xvq2STR0gQ+hkl+dI9C3PcKBXQUXQ/89kuz2EwJ+Y
WjR+Dg9CkMdafCSHgDIN1IuVw7HDsxq/nQPcTprMdva6tOYutvm01cAovJReNPGd
CLsw7qLp3H3OilupwKB/SC2A6AEPa+JB6tu1cY8sogWnKPMY1M/dTqNogJxlXb7k
NXxGX86RN4AVJLLkeCNlbMz5Kwa7yeW+itiO+2KsPF+HMD2xkZMiDstvB7iZHt6T
5QXUjlRkGJJqL0b8wRPAOou9zd5jvt+s9B+V1bhCrEE5bEldsCgFTv3LZNTURn8p
YRa7CzvK4nUOGQSN6It3R+xw/ik2c9wPXfJWZPV4VlXzgUE1oPhk9AWwUtlUmk9p
dyTjAF/PjBwq6kKSabhMGhogyart+ZeZtAFdtYwAU4+H8RtSK5S/mUWv76B8YMZr
wlH/cVfZjN4RrcD5O5oXrBAkCk/6co5aGkeJxQvAIpEJVG1PFqzyH+swFH55HFZ/
//O+3eRi2jcaPXAMX4QdqhnznW+CVXsRJWDgmVtgQB4gfGz4erOVlyaCpd5fD0fv
yEIYp9JUCF70GHDEnsT4hfAQQ6U8rBuYV/AFsGu7is/3dEeDp/ovA8JlPD/n1MsT
QwX5Bm4sRrx2dit3Voybpxc8CGE7TfQdrs1b5F/tw2HRwlVpsoCBozQyI2ZRl62s
SKiP1rliLiN7WucQmUB0IfhK+vHRr+7ij5O489Qdfbj6mgPESWZ8GcvH2NDa8FCA
pAiHnqTgZZIvIy79vHiEKPa9yQ9fS434bGgxhGHw0l4Mhs3sGfxVjNiqqq5ycSaW
WE2CgGs6p5zPJliLGsbsG0qIWthsKIEJURqwUTeF+MtEPMO8FXyVx6KnVWQIbyak
Nr26D1GaE8UfQQ/vkSdbd3YnoBCP98VnAQOwMAGn0CD7GJsZIKzlsE/Uu3Vve7DO
vr54p9XeAXb3d4MyUrpnJ447keQpvyIRr2tMvXlm0Phf4sVyTG4xo4YdOn0kRoTY
002lDwIcSdJfRUwO8iQG5R0EggbWChE3NghFwpDVnqkCycnXmS0pTssrK677ZeQm
LETPSXhXGDpMTHX4ezwzflvmVgO5SxokI+qPHqn+wOkI0Cm5/YtATRgAR+JWX0VQ
HjNMJC4wUxCChOK17DHDhy4fkkbIUdm+6KV/ray7Pqwe8HhUKHTlfxv3RdIqKqa2
7GIIe3+70B8uayS6IHLJP6s4DxouYWhQcN6H8wcwoVWiAnWpRqhAMwpSo24TftoM
T41upIMOHDbhS2bQm9j8mE/dLP8lZwmKIoDywk9JoXFL1GHcOOrt1L5/cVsA6Ps8
Hw/7GWcnpe9V1kIrdbykR0Q5NiTNwSWVkdWGeOYf2N+LZ7AEna/p95o5yafFEYqn
v0408dE8PU1+qfAm7okJ/75hFG0rbbvLmNa/yTOQVGWxt5BCqAIppg3gPyK5bgZ5
hk7ID6hvAY8Z1MVojhXsjObmDE2SCiql4xAvOSKEXIpKh8G+fgVGZR0/y7PJ3IN2
RTUv2Ej5GcgfALMyDE/INJxoqdIhAyf36tDuN5E9QibXhFFKwoekwdbU8tcpSS/w
6e6n76Hoz9yNRscT343jH2bja5Y+nDbYnFbQxTYm24EpkwWnqh6lZSG0rfxsaqgH
P4lsZSAJ3OqlfNDF5PUy4yOVBjTdBc62VVNnocbODQ5EfPTVfHx253QvL4Tjgmfi
1jK8OFyQDiRvxwjDpwqYXaLFtF7v20c/bu5DpX5LYbcpyeT+DXQKfJAjVpg3G2k1
auXNeLiYv7wJzbEHe2cN2zipRFANpPsKMY0E3WqbCrP7D8wgBvXCB7DQDMPRSMkW
LDJ+LBBr8uKIf3H4+1cmsm8D4LG33G7KGgRFlpKfuY5yQul7uMpdPdeABtNvjNeB
RRd7jR9YB1eZYiOynogFH3W/prtsV40NmEETp15e/6Q7Ny0rF+dePj5dw0LN0Ei6
AyQHLzAsDYH96Z873fe61r+VnqU5Q3P+qPlyk5lzf2+6Dg1HfsqP7dbi3h5+AcMe
oAY/NVdN2x35NyTRcIxz8Z902YdtkMUU1MwQ9NVMSuqPy35MLTXaS0qb+mpiTliP
pqmMXqJsAWvL5WVqT+WBjx1yp1bYxd6HPsovsOGfD8O7aza/+uyyM0TNSJ7IrZSd
ZQBxmqtZn4DMwDU6DofdKW01HzX0LKhb2svT0Nc8srVRbkDz+uEriDYWpbgZl+0z
qunSIOsVWQ0cJ5nuqSpTUeNV+UW5UZ5nLuvLBHWAGpgqp6aF3+OrGihnyCdqTECG
Sn7Kr3ItFV24mRjFRS/8vTtCqUSL48J34C6TGaoeIc5mYY+AtVpO0FpOcB/bV8Fc
pFYkvZt5aPcwXFHVKfhYbJGAk9xtneboTBBrTxTV69DIIqKarEvquAmallkg53Es
x/aO7QSIryn3BgHIBOSJ7tfBNYEXNrLGDOalsNuJR/b2YPz8QElGPYdKPJ6RwxuM
LUBxbJnwNgurGzv4mevgrVmgaEeDhsoLtHl7Xy6+OwwpP39NTrRmWJNbgCkxz80u
sxa3ZLe/fSx6z/w4xs2eEE3qA7XcfrTDbCo9ewhLrAo6jYRNhqtWs10V3v29lBTq
hsEAqpQuKyFmwnhOQieeFAbbFNFvrmSIL89XVs2hSA0rau90wEAyDVxIdektO3P/
4rG0neObzrVA7oJk0dtDo/6WtNFyGH3sSj2xa62lqW2ql+bAjFYe/rnvM6ZnfwIi
Oa3Kcgg2IlAcKV6WL0S5+JvOGalQkuQ532NL1LoxxOCZv6nZIPXQJz5N1sGTnZWM
Jkku+3JbCRFrCB/BRUcQK5yltmV3VobF11u0bCWD37rLyxNJH9AHWSKytxsxUsV3
su6Bt8plSw0UXDsAxL8ypBMRhROr4ABD2PcwxFDEykgBZxr/430gUblBHB5qwh5u
g3OXoFLkxT5NnahTUZdvw9b5XIMJ9T1Lp/7oYscB52zk8L/W9wd2YBTAFFe29ogV
N0sYDlpR2+Yhfakv/NPZSNlS/pd+5O6zTYiMdTQrHMGw1THsHDrYXUrfzEcvoAOr
62jdGjyC/CP0rL+jOFvG264JwMwOZ4N064WdT4xRlm1Badrsk8WCZbb+bp8heRVy
iF68g1NI3IM2FxIzb4goM2FSAOfSVyaqyjebRkArw2yBwMC1PAwYOrXKujgYWN0V
A+pUad/Ga3/pnVZzSTS96l54KQXAO0EPh1B4dhegMEPpSpqQhHW30HHoabIpV6yR
5KoPlx3mcDcu3Bokg3/l8kBnQG1bjZ2T4YMpnfj0qG5FQqPqx+lO+gmmY4o4roat
HmvxnfN4ax1hsggziBT5/aQu08DiMqx8cJAwCEjIn/ONz3J9yIk7H/Dkgt4pOGwK
v3e18rIPQCeEps4IB+QDXqaUERBrUlrKbAv7Im3mWKOW4eS1OeYK00fFRFCLpFx1
PZEMiZ/e14+XyuNc9GpPAsV9NxSUsOeX5GNOrKArivOLt/9HdJqXrR+NdRZMIqQG
Fchy9CV7ONnzpNYVOpum+0t1seXhmr2qu/aW1dXjEWyBDb8LkjJbmmHfWhKy9jNH
WzGrzbkXrU1RxeULhbp75FONSVlK5wxtfhGUHKhAWjMyxwbp7zx27cNuFFP71eZN
dUvH7n6EUFb+ofe1ioExaoOVmQOjfrsFAQS42aB2HyuHaU7Rai/bAR57LhEbVn3Y
mr8etnubq/vHQTvNCCaMpD7teFEhy6jzSW6P8bVeojpvO3Kqp1obchlP3YXGlAQS
mP6F7XvMfHzgnhjLjojfJOVDHarxeKX9StqbEKIwC1wvffWb6N/5GxilWoSNPVi8
6IlJoHXV3UcVNK8FeAYQTz9hg42iDrb5jSdySGaDPjzFhzSRjD89w3icXafmu7Xj
ux5uTydJSby1nQL8UJ910sCsFlCkDBDyZ5OjyROd2ycbYo2MAITAqwRizwqf2Gfb
d8WfDqV0lIIEDLNyebRsmYP/tpNMX7C7+8tEKSkznApUDwOQYnSdN0Egtps9pMrp
VnnbUXX3Ok+s5sEosYC7Wn4mlHUTtze0vJMBIry600XlRF6IClR2fnc6E1PotdiY
2KfBCZPqVLcD/H20dfcJmHa24LCMm3MitmWi+KC+dZ+zTxzECk+6mewpR2mIGhJt
H6gKVg2fQ3a8B/b53RguN847VeH0DAmjx+ZaF3kLI5UJxNBEuEPRrhamyMIMvXYg
36KZnF7wCisV6WSyBNP1z4xU1owJCWnCtNod0AaclNCg8gUVUdRFSpQFk4L3ETHi
+ztfW7/0bSfDMHULFe7BFxvbOR+qcL8SnAPONgnW2S/cm33cQ+lV9tzuib2GjfEH
SZLJzK8RhDhWrdTzMg1IoONaQxPw6+cbsRTnRiEYYGipV6R0jfCX9jhYO8FSO7PT
Ea4APg9ABXvn9aXwLCrH8T1b0fzhsxm+AK0Pe4wmwp/11548yngiMTrwr/OUUaZo
wrNdidr0SAhS+3grbiSrbHZdeo6VXODlZUjC5zECBTOPhR1SN+GmfEHjnXeSQc52
suP/aGK1zeBN/cA108zZh8pvkd74mE/FxYXTb3z5ltNmK1ZGzJYkRegcWPqk9Rde
ThW/BYQyrZ/eoHey+LEQp+pLJoRR/JalSO9rtId6Ot+wGa9sNn1W+KTndjtrJLCc
f6/Pp7zIk7+U0TSPKEOOCRah6IVO6UBdd5fffWwKV+E88EUAksEctHbI24NwbQO8
xnQoh12zCo8NjSlHcou5Gl7vIvWO7XHofTXBtMGbB606TEB1AFEX/3qZGxXMgH0J
22eh2T3wdGegN769HrTrmlPbERyF7hsWUGJNiOPg9ptRWzzc48ypNc7zwKSNnkli
6Ml4FKcVJGCQRVkd+6mOWw34WYRMvw0YRelcF2/WS0A7WqUiNN/xRckqnFDNlvh1
6X8tovHsrI/A/UVxLbVGUJ3ErU32vmDoq81zPoy7lD28cSZRA9wQ3w0UZackkSQ/
QmgKnwaFUMU42HHm2mvnNWn2Z2eHNfRyeryx/NNt1jNZMjqtGU2E2mMWewvrItDx
plOMOe0Jt+C5DMrx+WvRbwPbVk8DoqZRyyIeCE2emT0jtnp0BdKduSNVOEKtf7Zp
c5vmMYY754YPcjrQDR0ANW5444iiWz9r9oXvXpF3oOjj+DN802UbiCNQVnjcku/P
VlavLspgRVAdrv8Ay9orRRewGKdM88NW9hLXEHWZpDOrptPXT41kKDF6yn8QSWOT
Y2ZCPZLPNiy1qUxiZBgRamjjCkPjjvdjAThaDaDAanO7HEuVKN10hyABV6T4xbOf
F0Vud/zruOPtcY+s9HPfnYFmQV9GmqrCUZjFbONd+3ktwVEQm1eBO2O+gzp3fgyP
YwWgPyXsZoWq+h6nz3sdJHxRX7mz5UT6jK9ioEoTBRMYoU0FYjGolP2RbSeMkgbJ
9TPgUD7fHVqnekUVx/WZY5B7spaRWq5XeGjSug2SFaWMjpqfhbZHq32ZJ61J9yQP
yMimj9ZbkWPCNd2+9TAI3WglcQcx/Yo6YwWu+aA9yznKwN4Kaz5TIjv1UBJaqXTB
rQmzj6M7tOhtpzXbMB2HVGFE1DHARS/P1u6iUS3lduGmNkdUmKNMpjYB14XPA/Cr
NgOCuHlDoSZTg9AQP+Ac2AQZ1DvNimtso/7kcjr/Q91oOaZYh58XloZBfWArL+WR
3Y2fv/jWlvUHGjfg8aKx9srODImKe5x8x3bgKAM++77cZbNfYMt9Xg4086AflbT+
3sAd35fVZBFO/SeVf/eSC5GKZbPShuWYu8Wxka+jrmRqZwzTPN/DdewioKhLgKyr
74BMJa0/usCs1dX3WXKLNvrO3hmDAbyfrEmtyVDUeLmGRp8fDZX3h2i4xopSX3X2
Ze0UROup/r0SJqHvZ7lQWia9AYBoDQncPW16nc+UWqwX/WHJTVE65iOSo8oxGWmf
tPbfaJbXK5GxVDdQ3793yIyY8zqS+G4PjFgbkmCIj2vyH/zoVs9+kCAAyMPQhY+h
BTqPaj21xIE5eumV26wbAw6UxMWzTEIxuKlCHfv279EXhmCiSJc0jmFFHkkya6M/
LSYSqWAIflg25+evPLE2LRShhLGXxRBsaVtcFzSqLqWC1NktCV7XchP20rxeVTs1
LCCanH0xdEpf55Jz/3TQlT4Gdjv9kiv63GOZjscOJWFbjU4aFtIzVHmbLQzzxjrg
MafEAOpEix3i7SzxmU1sJOLvJwpzPAzTzqM+OTrj6uQ90p7VP8cZChl1Og7HB8pG
NDnPUduqnXjhVb+mPYhCkmL9d6JQKttU5lSvk9blIQlLiGY5OAxfOGwT5wtFvptT
Q1gvISJwfRTgFGU7pexgmCSXBnIKkxwfOG8+OgnGtax0upNfi7iwmFBGZ+7WGv82
CPPUMWCB7sChCNAtCGhG7iL41oiUsZNjfuxHCWL6lvbN5wZmqmwGCiaAiquneUkf
WwdHFmTblekdZHYspNbUGNVdmFKTJ009amQYhmDtoHqjXn7X/RVB/7fxGQMdv/D9
uVdypHKIhfMENle+xzLVezARlnRehQ5DuhmoO3jsoeoxeEj4897dtZ4D4p+W//9p
xD/6OtEjg7H/HH7VmHY3D7GyJP0TsaQv1iGjnDlDwttsROB3iw0xotW613L6MsPI
T0VLOCXz6L5ZnNH7yhB3LrbLpCK6ff2262dhWCHN9exXoOh1hIfofS19ygbRwPJx
jpdfSf7zaSV7SpC0dMB++SmW9kDq55GZI0QUD8VykPo73xVRcB/2aoNju02oUnL/
6Lbux3FeK7gwNzGL/loBR0GOfHOIAD+DbCSrHOriHfQC3E+whKU3qb+jvzU0YVxh
mJ50rVAkS6vq5p435RLOo06m1gmuy5opzYiW6D0umEL3BGV9OjtBiSOMfl9hMYL7
xWOqicrpuZKq5J692d30CjZRrqLscxvgDo13jivrjHQfiLHG9cA1/k3Q/7MZUbIC
zK+jNZbG8FX0nA+MgFQp1Rtwti8qW4Dz7zfBzeMDYvMIrQDaoCSrNJgVCGPKvXHJ
uhCZu11BfYORBq8DtAPlFvaVq1qPxsQVZpYqcftbCZyFk6LiC0/exhKgHr6Q5YVw
0/Swwa5ilOmIkU790JQouVRzKy2MPlbO4M/6AMnX/msEG+fAHLhpXPdDIwIPD5h9
ZUdUu6Bx2v5dCf8ECNEneo2I4RE7rkDV9tQAEf25Pvujz4CsgMJKT/lWN6ftO0kV
WKIkzOa43JiEw/SOiUOiHxX9g8C4YmTXNHDGktM/pzBQnoBpVgKngHrV8dspthQX
21b3lj6RPG1U7EX8JJImjOJo4qE8qPA6nvMYV/CWINotKu53BXakiv+WJL4u/4ZA
C66JM90kwXHSDbD0PCf4ZZtmFfvEHO2l8YD5XptPpVe2PL4NIfiIfFu6PIPU/Q+3
biz9xVEbit3RFFvgjkenzcHpFt09Pn642hFdJWB2Evonaf8mt4mN8uAooi4/pkYp
byF6W+UGnm/nZmEmLtpbw9XQGtg9fUQbD4LhZdvsJHG0vBxm2Bpr5/bFnb4fwPYx
tXksC+vQTZO1TMyOLIqWNAMt86S8bU2NAO9zGi5WqXoK5w6fP4QzurHSEmHWKF4k
pvB6tehH0XUXemU54XWRcoU7NuCIGjTh4Wm4hS5r7Z+l4ESEbyeiMJUqc/nPMDk/
PHWWJYcIYIfjXZnWoO43Rs/Y9BKBH3mrVs2Gp3XVzxNo3zI12QtTZTou+HNlP6hh
Pric4hiaAMlKcSnWTi8hhbx+V2tsZ9V7+6lUdqlmi+NI37pwv3cdzZKPLVRXuS7V
5xsnSvdaiPVjQbAXT27Cu9SwTtAqej0dc/Ui6mspfNoMh+5LS+iFW/b1g5XOwO4s
QjOkTjAtspW5JREVYe6Q0ISGD2BChlK16fMv6J0Cow363yU/gdHEGeWAYFa1PD+A
u5knbApAtqVq5G/YAx4RZhBP/giLchCegKqtUR25WvY03HBSHh/27HGrXd4PIDZ7
5ADsisU727k8Hu82KT5nyG/ZtTb55ZVsKQjIQtXgTk1/AoPu2NR35xAvDV1vs4mu
Iw1tTcR7Rtl/8NKuWwfd21igmHB8DTrjtmGlfcX4luxOBQqx7KQeM/UwpAk3KDQL
o3pWmaI2OSBO8sv/HKN0yftD1Zf87zAHNOeLagZ9zk5AQVozxHme8Nj+XA7abwqE
EW9EpC+6mo4S1V5SyaTm8ncVGD5uTuQtqr/UrDiriFJOBYfnKnQSYobJNNKvdnKP
bgY0QGD1JgrEqEZFe0eggGLBQAG3kLqR+Y5tQ554DgZj8AEwnHfUr7Ns4Ck9wL7C
ifk6QsyQfRPO5Qe4ijVO9CxVqIoddryWk+gO7x0nAIb46PhI0MOubLykgXjR4haH
g2x1ADqJxiEIHqwgsvSac16NQKX1ayFoZcWJ0MbJt0rJotBNMYRXVhVoXRydgA6H
9HLMynhNt1+IRqdkZVJpttSBdmcCwHv1v76Spkec+iP3PfyWWbZDRTDiR2qJuv+d
EQd8UUPd61lDCMpulkmNHlcP64l3LpJqNYg03QBkisZsamH6Lkgcdcd18reSQSwN
WBCe9Hwf6ldq4By4JdBWc76CN/XPbT1IFe0HrpJB6/QF973k6XKkwv1+/8Gccrfd
v6otRrhIqLzlQG++OZr2VdnLEjX4ssZCluieId6+CcIP7KDOeet3BU2ti/h+ddzP
/opixj476GLMGPLbgfzGGP5SZ7MYJ0YZYZVExIVxrTTe2nkBLHqMRMzlvx3hTJqN
vMzx0rcraCpVw5x4umZIVSm54pGnMM7LWLefX8cFhnTvRzha/nqyW41aeLrD8fTX
RBqf8CX7RLOf9T+aYlewVwX7HcMRVURWF55+2q5NckN9h8yv9EV0Lukce9d5f34X
PPD8sA+tWD3INMSgNKMB7Sma/l0yiJ4uIN02S1DHg/b/rqtUGbJ6OTCx5yczXqzT
B3sdObkt7wYkRrLVr8JQ4o3S3zJnkbK/8dgUtrtyGdYeB/gpku03GJt36dVImV/2
OlfSAI2CaIfZwtxQ0wc3e8j2aTLpyHQBEIm4Rkx5rImaJBEbYV1Q+eK5CFhc6PG5
O5BOCcBM11grapL+gtv8ej41gUadOh2AV+fwBwovaPqUnisI2JecPke+ppc+my59
7ijEDXOPmp5csEvgv4R7UZBZ/Nkh0cHq6/37hWt5p4Q/i6wYCTvOTgwCcIM59DsY
vOxZS9ptxJocX4X/fJlFgicIZ3Zs3W65o/kLHEWD6V+QhzXPq1TkafrMnjOOfokC
K+CIz5aipJ/imkPUIOu+V+vNH9kHvLPjXkXMF2OVuzczr0GuTvxtFvlHjrTFKqqn
R82tlhqjh1k834pjX8R7cY3uLdIC8bo+8cq85hu9lpOvs98sK1b47jtQGXOvsE0k
sajS6nmlFEPwrX5eti/PL4tphsRmZtIE+Fvle5Y0E7Bz/906rGyA3nkSkfb5+GdU
QsZt4Xcw825LniXZVuXcDjJDq51c/n6zfx4K8CXeEpTo2XeLCp82Jp02qUrb620r
bTPc8iuu/3TDgUBOWEIfBvOV7Fr9jC/fGv8Q1Z5ixxTUbJg/xACvAUzIXYFK0C04
WFmTFS0Bgi1Rs0g+AJ1q0yFJGjlEfOuzHzSimLoLDvnZs9Ie9rhOvcIsBOh5DXWG
I6YDg5H1/zKkB5zdoXKweRuiGawHdVIQnIsHy030RZ4IACSoEEJ2T01p+7Ufpxcy
J7C+L105KBdBxvKHYeDy2EH2HTRBfhVNLrROEQjYjlhAA4Zx5JFaKjF9D6P1J7N8
hipXXYaINYIhf1kSbAowWJrI62UV64NxJvn5uvUf+78dngNDSoqe65/pbaq6Sr+K
F8IsAEQ4j75gt6J1ma7aLA2mrXNGosNeJn67yjpjDKn9O9E6I0TIXZLmFfEhrCu6
W0VFw54OoFC1H4Hgy2UBa86dSHuY8jfZFbKnVfLIRy8bNdbhX68xho0j7X5tDFh4
2zltGO9pnnINiW68KgVUuE4ZYPPrwjfEX5V6GActqqsUTqFZyMxwyX4CmFrPmvDQ
rLAshjVFo99ERTVTy7lNWh+GrXbovQt5LmmrLxwNedebUXbBPPMzoa96rVfB0gLE
f8ya88lODwSW9XJLBpA6vpHQ2vj7JsWlBgMQWDkIuGJaZAHCEiv9AFY20HMdaPkj
GpqD9YghBMpQgSyASzdqWa4d4SSN2ees3ML09CKxsdqaJKxUuI0zJoQJ/BA8wiBK
rj6rkDJ1msXQ4KKsJF6rsdrCX7VMMfD02QWDRlbmqeQkuNbeonzrXPZ1cfbbGrIA
UeGHezJFa6kB6HKgrkWkoYXbLM3YP0ukVUroXkEltJs+FNQMg1C2xBdQZBvqwTX+
aMWps2+Ddl10L5Wy2nw0AlJ1zwOxzjIEFSNU0vflW0LTBhbh1iqk1ZZAU7rpnaKD
0fKIjAQGxUyOPgoLk05dgbbb0UHRBXGzX5bJmP4sk6ap2NY5qwRAA47+wSiwtScd
R4v+zsd7sGEpLZmrAvCpSaPsuhligxl9i0GrE/sAk3CQFlDhQwnVolWQKgV6wjUJ
V3txlJqxYHwn3N7u32g7chpAVyCKLhXGKiD1Pn5p001ERiGIhwV5rhtkZDti60Ut
4mvF7933PnW86eq5HJxo6jc61YR948dtTYqS6V1oNooDQcVYKV4uR+bIHzrvQYBW
FDA7M+LOpf61fulGx8uWFgprDTD9jP4HfZQcoi84paH+TJEfSbbQY+7Z8tpv7voa
AvZNh8wDuCfRt24E1XSafugfpfq3BwfBhRDjDc+CpGyTZ+DQr2n4lRvwexNqxben
XHfXdC+hJbqctkD940OqIN53YyQzFVd9HrFX0R6xmft1QqSoD42vb/KCM9gE3ExP
W0Ekw2OFDE15U2nBZ7FSmFNGlAzZAEH2bpnn5afLTg/7TY3Dz1yEGwWyCTHvQnHk
TK/z7QIT8GkF3NUPnLKEKYi2hlUAQAAFSucAmxSSaC/KDbnmy8/M3MD2sv7+n6IJ
z6ga4Id5/2pcMAlHYAxfvrGN0Q8if5iKkqEXsjVCAM6oPR8A9v9dQ29AcayaMUt7
fdcllOlksCW+5725Pfa7pPqr1+glWX7Wp56Cyl8wwpVov5TbNOuc8S68Sl2Hr+wE
5LHGXAyfGF2U5wTmf3rBew5lajh9I4DZh8DxtgTTAB2dMLs60KSZjDFb888Q9Eyh
D2giHjvITzc0c5Mx82IlMzV9/Yi/SDMk5iB1qJS9KHnvZzkj9xma4W6RgMmgUN2P
oBNbn827HxgJtVBKnjf2VmoWrryHoinB/FhvDGDb60BukUeerITSD5TD1lX6+fz/
xoH3sdCLPQe9lpERwEdNt83UbUTBN6lL9g4saKTAX22jUxLX3ptYzizDitejWHsB
sddw5ZHcZGtomG4LG5wzQXvlD5UG550tyzqMogb1TMgdWgayrWuyzCzy39KWHqAK
oVg+ebdO7GDYt3K9V1B8lA1f9cA/iXNf/Ya9t8k3Q9ATzBWQ/6B4B8EFBTdKVMCR
yyKjax3Q3tp9XF7AYHTHARWZrcLTtT7jvWtUL/EOTpnAuVuT5gIP0VbQWsTPJiKP
WjBRXbU02705hSutb9gFTxUNeBMLWY/Y0CxNQSTEX6MaOxl0Zt+aRWO6RUVp9zgP
w+WKOXKl2KTnE4x1q0aWgeHQe/A7n+za+c2gyfQ6mtCNEjLreRFhk1o5Qgc6/XBD
7ayvjMnqHKM1+n1+RE8qn7uVgdrbLfLOoE6dgCwLkIvpGoGjqYiRrY0gCOqR82on
plr6GXVOuaC9h+lRtxnZBYmkCuOEnxZa4BvhmMEsc72Jc/ZahslZ+zw+V4a0rmY2
YXL159Oshj0u2xXwX7H3SrgoyibV+rRjcZFbgD+DQlN3+gXCsxg7WbT6Aw0ZvfZO
gP0sTrzfhahV7wZ9CoL0J0OwGr2yaSovvOLhona2kQqOJ79JVQ4WdHUOBzVQWCoW
+ytzOBlWaLNX3274agTwoJBiKNFL+CGnv+zORCqZxnPxhTts4jxVXauR66yh6UsJ
eWEG75lXgx6tV/t0nv9/7bJwhA2Js6fr5QrmTsn+nZf3DxBs/cTqErNNrndNG2md
wTGqKERgSOrx3umh8hNaF7TbxOkOVcHEQIxU3VRXeRbmDO1M0lRrVYqaOVpBMZXm
KLoIjeSKJ1aSvJMxNqD+dqwTwGecQSFvoBQXNt9yXr69AUJ7ywC87b7Gsj1PTwJG
yATyYbtoKis+1HQL0v1iY7vOfwQdCnPgRZPd0544/YY8L66lYcdH2Y0aqfIvmJM4
hUPy1Bt3wuFWQlLnakPGAwsxS3/PW1QF98cHeEN3h5rJePkmPlrWcHfvESA/vMb2
wpzw32xq0Ps6HNIV3EpiJeOCVARRPZObuEh5QbxEUKsLhS8wRRRHfm3rlSQBRAJk
Wa4ZwFZLUPebKAYZ8VbIdSjtmX+uGVhtxMNX6N+PJItcyDbAyJCMbhSDoRKofwHm
YIyJq7HKzU5gjRX1ZCkhH4zdyzvaF26y2zCJDFhWO+MJ4jHTb2aXacaG6OIbNRkJ
0oMASXUacJihYTV+QkhpHtL+mdcx2gOA5iSTBG32Qk35jbqeLv4840/iTGBTHMSs
/ZDjS35Vckb7LZOej382QShys0fACOszZJowZ3zsHZJlljTuyk+2u3TrFIGJdjAA
qr2Qodn0ClBfa0pEc5D4YWjdOErDHhkzcW7KCbdxVDdLQ/1OgSRrUDrb6qltpMKe
enZgg+uS3tgzwosoaevAx4QNC7aTKP+uh81JuyQTQawo36ZjDvrFYejwn9Ez3PqA
zgflEefmiNeYxQ/CSKNQlSheJ3ZEMCGdWIlMEVe3d8iA3J2+TXF51fG2hKDSWfWd
6ID8mUQhYV5q4Hcb3u1+PEhfxd8RyquvzfqOvdTVLWYTkD3KvktoUXjNiVfIZ+ry
rFtkKayEGZqOUX3usS0d58pVyWcz4h8QAw75wH0TZ9h6V91X6ki47iSIYnIK1OS2
+9ebr09bOIFk9UsEZxSKJC7+yxF/AJzIJ1LdeeBupMBUCVDiOTlHa00fCSEQP2ne
YI16ajT7IzVTFLz2K6EQGekxG2ahsBTFqzige5ucF1qp31reMMIKdZbC81vBR8t4
nV/3SaRY7Zr9WGU0q79TnipjqNRtpdRpBbVPlVOHig3e3OUFjzRQ4+FjfAdWOuAW
Nae96vJyU7OM9SU1y8RdVji9wFMDWjzBhqvgjmBFQLz3CoGHDcgdbtKRCwwrywxa
sH1XnYhgjn0q3jqKmXjB8KyXpVOvnAiI/VNIz5RtKrYAN9tvDhTCPiRbVNdxH+DI
LfpwjFsMRCXmf34QYyXiiVdzcPu7FHH7KmkoqtzzErQwE7cTcg4f8P7ml5lCX0Cj
RNca443gQU/atSoF3ZWlAP00+RZaiD3XMHkjJu7r6wnV1bFqKQe1lUwAdVMx3ovR
vphd2RWGjheNLiuxTrAKlS+EexniQWkMLAsy7hA79mvRR723aLEzzRefulEW63c/
mtEaxdRAqJXExczEg5Uj6Q4tPWmmHA25VWZcR3ViUrzqlCvXjoQoZlleU4XGklR2
WkI759s4PzFO8IpM1M6YBNG5qtAv9/Uq6CgUvbv5Z8Eq3zF6uGwnJair4nxoYZrC
Ud9xOR/QUowLVly0lc97PT5RjlhwohI/osy9miQ1yaD4dDsZEnligJ6k+IBmGZaa
5k3k+ji77kO7NZYCSYpG2fCAB5Oi7dGKy0qy5PudzFSTrz9KiqnZ28FiwnXzxmrZ
b7Oj5b2oKEMRjM+YUFKyvw84aBpVjMQb7bk9O0Mo8wENtemgbTUPpdWyTBO0DIvm
KlSCO1jXpjNUb/jTUBNnBzlix1ccqnTvgjYGDse4kUqSXJASOD4lVsn0FBhhu8oM
ZCeq+rCnAWWAJ9lQgO1rA/VgLhTJ2+gQ954HXhX3Jwr/s0Zq0yUO07+E+W25Qf/7
aIOy14n+1e67R67RQNDo6+NtLoYracL7yyfONJhM3i/djVSPdhZuvCDKLy1Tkqll
z7hm9D/3V3ajCdW3XSCPYA9bMrIHOaL6Ocs40N540QDZfjt40+YGV3Xp+nzmqnVN
fnHZQo2ThBhs0fKMTWcRXX2EQvcj9yTTC1sBTnjgCSWkZyiOB4P7CfefWJ4Mp1MT
VU7lt28FnttO7ffsClIu1ELnqmHHBefZS/JwNspA1eShICdSZdZX5n2pNG7+E2Ai
gRTh1fivpEZMOZS/WyaByWNdapG5k10mF3HQygijXU4/LQ+hZ0uMbIQ+tgQPv0NA
PLIFK3yLu6J1uB5d9U+yG89U0hg+Mq67PUXyy+SCGtbsER408bhlZEkD25MkUWrO
2aQZLpE655HGK5bItMLA0eL0d+ASG1clGJfF4F2QU/zJ3YyBrM6Qc4FRL13qg5rK
uPeMVVVwSGY4GAv0ap3TFHq1bnByWmkEoXNyjh8McKWtiv0Q587kKGjgOnz1GWjz
0qm2A8ngZO6VDt2wXmFxge1Z8TSXobPuTcXTXkAiIAW9nI1VXZx0849UQ8Z3uhAz
0nw4B2iMmNU5UuZjLM0hYjVTJxgXSxaSIsJbJA6dbDVI5wfqWz2XGrd3sFPeP4QD
O+9GPYKgAnfCA3LxDpO4JV0og6duDMLqmY1XJMIezDlTVBi8sAbtQUUMkVhRda7B
XIEwT2TkiWoQWuvIR1jgHxIsmqNmm6ji9NzAl5v4UUB0KfYZMnGUM3ZpvuoWV1F1
Wqc4TeqK8fiIVWUy+vX2aXDY9tTh+Iv1i8ZENQWbgyzJ3eqMtELzUfefQlMgZV2b
tzZ5l8A1n7KcCiAel5AZkJ6m07XMIo/Xg7XrhLoFGUYYKWktMgXvNHN+t6/n0Uzr
6KpDsGNweyM4jUpkG4peZVPWt2rnXtY0HARURmRkKbhyjl6EYzbWHVrrTn1JcWDu
/uI82Fd+KogxtwVw9DTQqaECNqcJ4mt9slD5XbnqPDFUumALTFbWu0BUqP+nIgiI
S+WX+OLig+JHpgAK9bysNF7yXfCjbueUnsWbPymQrjkRehJyPjgrruYGtQmPqu2t
vwtqvm89cNxkVqiNIiKs6HejkiSoF8QIdEEGD4T8pXfl3s6pb2Ekk3H1FCSVBVLz
96X4yyQPi2/dA1rQckMfQcKe70X26e04esEQxxeER1pAj/qDmMMdbDEUnaBEpc+l
ixnGjTp3lqsDI174sqBVuoQ/pTEdm0dJ+mp83f8+H+lZc2YiqCwo+LNAONzC40cM
yNsjtW+Lbhs53AklhVyE0jyu9MB0AS7w81uUXE9DsKKw1Nfo6Zku07yUxgy8fwQt
UzHx12OVOp87jWdbNwtuFsDpO2NtBrnIUuP+MOvU1qYIqGHaUQmpX30YByHJA5vq
Z5X7lQvqVSDXqDCl6Sd77KWd+UmobjToeLU58t7htk0b57emAHV6m4Q/Zy1pf4nv
bvFKiVSrW34XOEaceUJmdJhFtUdjGNrzVnkI8mJ2GeoipcF9rs+3b393JFYsz1ei
WYuM3jdhXd380Geg/jLu2451o8sT1qa5ywvtrGJzfr4ryinYgJDOPAbXYNkrXt8a
gQi2z4uKGyBPJqaSf7Nsh80TXK9k7Vi0rBKNcVlGsr61a7MGoOmjaklt4o9rM9B4
qXLbmeGwqleXOdNKX00FfW525hYEgmeRghZcLON4IFsnnHuazSuP+XjiK9r03NJ+
A4zQs5md73fCVA6UliIhKCrRGbOaV5lj5Nrpc5dOarWFMfdHkGTZwLOPTC6/nxwR
zeNSTztc9Lx0zbZm2lZueR1NzJoGY7+VxEROrOnwoaCFG9aiQn6yNbo288z7T39z
6ce1sGWolP1lC255k6d4OtK0zuIu3cE6zBBEPkPvRLShv1e2oX/B1npFeqi0YjMO
8m4ei/UFO72Jw2TBs8nIjflL/MupJrgC6XYJtNZ5obGbCP/ffAGXSke/ZzP4+lri
WhlG4Aa+56QI+XcLoQnvQ7qvJgvNBAhmMZ1MqDfZw8pCtYEQ4G0J6OUx/S7BrN3/
tUIwa7JmyNRU7+ZKr9YcqXf8T/D/fg4VHzNrrM/CG5ki0Bn8oTX8t83Qt3KPU/n8
KwwyGWZ7OSw7rLPioF+3h2mV8d/CFys3jLCedvbz7Ays0j70/qUpE1ElabntELBX
d7858AXVnqp8Gx4wiCMgWQxvqdrWkuzubnkWFmtTTwmca0Q56ZhdqWwKYVrlCyFY
7wxBXN5euETbYsAYeW+fE+Ib3w/sefQ+kmDLgxSBOBFxh24SpOL8NB8FLT/Jc1hb
S/FOHAKdALWDd8qS0QXnnETUZjBoWALJ1OoHDu43JDT+3I8ef2evN/qdszvLTX+2
KlqhgFzDWvo4p/zdBrtnjsFGRMb7lk8f+ebVBCVH2Mt2+ZK+6fULe42rKqyQ1nUn
eSgJTeFZt2nWN0bpXPX5NT/M23Xv9vF9zFVzn5g7adYXcpVmzUmwM+4MPTTJhKNh
rmfbS2wdG+18rLk9lsA1yKUyZylra30XNkjqqs/eP4ayL89PcuSef6jAHjrUS1Xn
2JVudeZZayRh3adnaTSvVwPNSNCR2SD1mkmBCjLnPOlrp0TjuQ+ndtx11lx0GHII
txYUVBWFbV3Reji94PEPMLyAORt9Cjeg/cjCowxVao/DxECjMiwp7YfeAm1YMhxJ
XPFVQIuZ2mDmTY4Ma6TXpu8v1LDq6pNWjLAAVrcPTRvo7S86WyZgcecRnDPyf8C3
qnXNsyR9vYoHLz1v5XUGAV3+0rCITdW++M/xXx99yr1Y9alsHJN89HZaOtaVc+zW
P/CaJyQA0JoTp7F9oWWTva4sTOkAAf1GlzOF2qSi2DEQ7VLjTE7FTeGauhLxZ+f1
tR7bZDbEH0NQX27xq9N5pEBa37FcSqLKPEO2QvVoG7V3jYYZPZx1I9ugUSjCMbMw
zo+YxMthnYw9brHuBcXNCB47EcViQ4/bjU76XsL4VfGkTmYGy4QQpSJIW/G6s74o
Kf/2NeDVGD3OX8GbFeHK1FNMLNfPu1FUnZs1wRJsBJFNz/WpIBFK5au+DcHFDz0d
/H5wpxyVaLK4QL5DeFvL09IX47bL5Qdp0QOH1lGFXDaSd3RlzoXruoHmgBiH5Sa+
9ZOXqOeHAA+Q/9Edws9c5vI9p6DLWVFGmvpiCa9g5SxnkGHfOKTD4NRPqOmDQ+MS
sX1dmrBn9E3kTvS1NLUZqz4S3RImAv07p6A2J3fS1tqvv2Z47Btew05/iwzjMqez
NlImYxmwTlFChM4XBHFqgzQrz1mqJoyWfN1wvH/p+Kv9hRTuoYIPQ3MGrlGSYbVz
xY+SogTf2tNqbtW3G+VgM5RiQg/fPaizQICOgazqYmnzlVXzktThMfsA1fGOc+Lo
k8eeY0ToFeprpGEIp+6pPyus+XcmBwK02Gr0/t9WCIVcn8t5qRgSOe/iwh8Szvd8
wzjZOQuFr1LH1pdMKb4SA982BBw2DQO0F2AWYXK9CmYgr0Qw9rRf1dwRPTbxGlXS
kyk3+Sa8dqIMQ8+R0Tn7fR2rsy8YYkHR+0Hd/MDD9VrICwE514Perp5JNUcXupQB
pCs6h37s7sC8NkAz4Klb2o/11j0+JNBiUoWnNBouH7kidxC8K9KIeQSyuzpktWIu
n1aDGtdNJ2XGETZzpApbd4hws2+sldzVaxFu/PdYPYObArWWhRkoTKjbVeAzD+aD
m+WwJDZEkVFXnsJuFv5Fdrjkebpf5IiuxSHyIiTOG4n4z2JgW/UtX63csaPw/nAR
wEhIY2ZFkchGVBY2dWGHKC/MPYtVctQYfQfeeJK/iz++NrJl+n63IT0zukoTbW5u
GNRCOeJeNi5Z7AiG49K8B17Vt8gbAkXFQiLFFlEmzpG1Ud9Vgnqg6Y0aA4v7ogOi
xg44og7mrqnaeu3WvfF1jkOq+R01ZEJ1624golcF2rxW2kXQiNR3RA4EnABNoQ1N
ykbGrsTb7P9xOOCe5mBvs4A27dHADmt/Gi2TNgORHGjzbm5BifwEuWGQwCkRbnyZ
+AQCYi40RibbgzZMKOY3rict1PzdXJKnrceKdQr0ttokuvqjnGvU1WGXWvVpyMtk
/vo7bdsaL46x4CsgRuLX8jLTBd32nOfL3CCLz26kaPsVmdYsDXBzCT9muke5wXRT
CaGvWjzDynk3bptsrm2VJAzvaryt9LF7sIxb/Q4sRRRjBRnyjF0Me5h3+w+01Db1
X0ALj8Hk2NqW+w/qVgxlGdqWDl8Of8glcYd4gQcKohRB/AsHUpnjvZpkiup+e0gt
4MsQV5LAH296svo5QDKyq0Ii7b3PrZTyUd1JS2LSAdKlAfnsQ2JrQ3w3hDtSPgN7
zTO1/ghl4dyPtsHzkYYXVD/0K/v8YX8h77JTxPNXf5peyyznTkqFvHtVUoH1wK7a
uximOjQSVK2TrybbdHBT3ALt3Rb7aR1+A+cpm58KOn9EZOXKTHwWc7htU8W8QhO/
RdZZhZhvBn8tYDwlfPg3rMG51Y0KkVdHzLrJltKoJETQfXDyFZB7/ZwJAywUxkMe
qOHZxHOOGfEITJVrmtBmzoh/wL0r/AkUtzdh8xyQzAk3CHTVefu/BbBSmWX1xBnV
uhTj/5jte1QiCPDaEul+0TG5ejTe8p/MQf+fCFINYLFZc8ZwO+driuGJaI8x9Wia
aBz2HZf4u5gpL3whCYhqLp4LkT7ccfcGDiHGkAIx4QVbsebDi5CHgkSCGXiFEzIZ
HvU54tPlaksElAXp9+4hPUdbly+COIv43SJ2fCHiHopYDhUpyHjCIB7qAwvM0IaF
GgfVfEr2staEd6C0ESDDa6f0GuC4x0VfdYDmYQ3JIz9UuJMKD6AkjCyUIXFmmcm1
l32L1kNb5wq1RdZFqvXRSErCYFFbIsV7OiHfvkOhWWJxlUlL33EhigXYFWFjSJ5h
h0TF6cxTYvXVFL9ZwlFhnDEX/rMAEyGo3XukU83If28bqSPWtFXo6TT4agEYoA+9
T/kBJwD7w8WMDKhnUsK3qEK29ngTqBT4fRM334gBJZkf9vVxttIYaRlaTaD8CGtI
Hx+FhRgSXYgpEK+gf5xqWtWQORgPktin+ZJrwp+GgbZJmLHKe5fDu2tkCDs9MPmf
In3Xd2WqYqyyidyGpodXyXchLqtVpfxsU/W9GSonCVHS3Vp/Q/YtBAirfCfBfdeA
Wk31I7s2gMn0xrAc+lN4+tfMBjUWoKVKDD7Q+xI5HhOkurppDT65cJljx5u9hFfY
BiFAYsmBLLeiomUNuyFjBgDtM819PBFVL26SBbGA4DbW793erv1DOdH2MGsG3JMB
Tc8Vk9W6S86Q7Wcwb7UHlgkW6OVFGepgLAOJA22HqtH5/Lo6pCh0ne4IkzwTU6rC
ULMbx2N8hecrZeVsMiIyIYHruT8sM8gzCl14MPO8sCRkBqsDTJdmWmppLdLYNlOl
7La9a0BYQ1SGQYJgZEErNXrdBke/qsP4UsZuDPjsM0Yi56CfVpaujBArzfg3g+Qj
yNLTOuoY1kcvkbocxDmRYP0fj3cVN3Rq2zc7UGeoCOBqiupARysV13a0XMDXuVHj
lA+G4TVu9dkw2z5V34M2osXZ4a1c48IT9G/7QIzvFlsoShbhc2XaQrySDXH8whQx
kCPjsdZoWcI/YdPCjpV6AHrps4OWsJxjUvfPlLKrGIIpvwZTalXQ3Tb/YrtLy/7g
G2p7EyKlb3DY25kZEC/4BjGz9Jb7SY66AUkrSPP0nLSV2BYsflTo6qnr9V1aRYKY
BKvBlY7qEMAur8G5uPdZYM6O1C8ke7fOiR8rJRw/1PWY7h61az7CJnrmwgmGyjb0
L5GJPGUyBu0xw1P5ZD0dgIMIzqw6t4gTxzdO9OXqNDy7ODF9PUnFkCAgS4tJyz2z
17/l5G9g4P7vkgRa0HlkD+8yEapp3KPuSueaZpXDQJ7Ux2VdqAouw9MqUMCi0ni5
u0vOwgLqHAw64BK8oBteFWHezCzn6Og9w8JHcV3ntyKTNEU378R4/rAVeRvTavNX
w5h0Lsqtz3YYIC9lmWVcIHSDqT7MZNhLiNkyvyAVqGyUeufcR34dkWFok9CtfeMk
AtOgVgCx3Ciifnl/xlqIAN+NYPAauap0eS3ihSx9SoZRwRaz+G/QDK5VzoN5oo0Z
6831EP6TCwub31G7FFcHGktfAzblxstlz0uDsdr+aBhHh0OO+cpgj/5w62A6r4fN
8ddzXiSlU+NIzXCKfYbpdV95NwPBoKaD2Q+bS7C63RO1OTUQ7c11rm4hp9ZVdYC1
UwioRJCKf/JIXXGQ1Of0h6SKgCLynNpxaMmY/sCGn+cWFEmykxdavcfoeEaze7NK
3vO1HKlBHmqc/AkrFtQiVGE477DzzVkR08MpxCu0wm4ye2CgBhsxBjLPo5jYC9BP
3pzb5F8SZACqzJHw6vMY2J6LoSXBK/lkjNtUQhz3eVytoGdo7oX86Eb4mltiqBo9
cyGk3a/FlEdfu1g9Lw9ZMkODU6ktC69Q8lDiaDHNYyyu8e6aYc1mExhB6F6fcqf8
2LbSOCIdj/GPy66QyHJaF2Pz971KrURnw565SfStt0fG5AGr7jMnc47QPoP/DypT
4nl2w8rRwQPx+pVFb+Z3BCU3nlQaSV4ANWhVurl1nMkTvkHL/v/MVzYZOXVrri8M
Nbc2LkKXg6lJo6/0b4Xsya3zHIlBBjXkxIe4ewKfrbLRb85KsC4F3/2S9ifQLdxb
Bl/uqdWBUXQEpvwGl0JnZ8CI7FUyP0sgTQ7JhjYZO0cP2EHYGV7nfAqtgF8LWeQ2
0EqRQc3hFpofPZt6VeyevB1raU5QFwgIqK/o4yndrMYldKne6FSQt/rHftP1NrNS
W+Ai4GLzdowxhQbdSObVafhvlraCqENazUGcG3+OwYxTvxKc2hJ2/hr3y7Fye+Wz
zdzrNfSqSCO8XfCrPpAczqrCsAsrm9HtxQawclU3V9Q75WLBT7Qyy3P2jxTQ1EI/
S2amPqhEjE9mwKWcZ5HQV4RPxz3Jo9ob10Kasnyvd1/F5QoCsSods6YcVnt6jAh3
AO6TVv2WEAIQOitUlKhuI2/BsJOEJYXty1GnudiyfH9qgwg68LvPmSvxHYANQ0Ei
veu61lhKiODypGwWtC99+yniBjzySiKEdahLHnhGZZXzdq5szWfakfstJcw2BOaq
o5xBaYsL5zuequKlnf9ScqJ/NS1ZEWweIQvu3iF5LI4vT0b1AgyUvQqn0JFu8osx
qeBzimXLwVvYT78CkgJLd5gVs/MYPwP5n1dL/O4063WvvgZkz6HLyyPUNll8ZeUh
XfE7M32oklsIa8FuyJRlcFuelIRD7ATXItAwOuBbBM1+vySapJe/+s7qBBdDJz/8
6/FKSRGEdMU+dYZJ/TzEVgHZt89Ckq6EDE86K3rfgRQLn+vcJ53pvLYiwVlZGifa
6IgrQshme/vlZ36ZkjIgB+ZRJOGW00+9pCed9at0fO8czohjk9YvZ37JJgAk3wpQ
hv+kJ6lqdpX52HpKM8nJsWYlc4bGwnVTGBZ7CUO/tu265qDChkFGiFdAw3F84+kz
sV/nTsXskWzOWbkocqou0mF++DBJqDQdn5/NKW44bBMRdz12WHac5wSkFfPFKunS
mXP0W3YoGHlmwunp4DdgjTWTrWl1ogXLhEqk/MbufUqeeFIz6Oe2Zbm/U/UPmb3j
MB2nRoaogRh6RPk6oKEae6IZqB1mtcU07tR+j3pIQJzk1PFqub8K6Wn7EbqPXxjl
G4fIQI+Yac3A0Ah3FVQpp74pfqXJkqEKPnrv+9rnl3oXOvP89m701ZgbXB4MA8+N
6CVqDZhFLdpgD7gBDkiUve/6gb3dtfAYxmul25FFKibVseI9sYbb22IPXIsdeSPI
smVDkkRToL/CqZrkrnwfyL73XL42ggiiGUYLe3ov4UxQPjvL3ez2nB/iBSFJXkWE
ghaRx4NJEbNwkp4cecGk1IiLJMDiDKg7xWCFSgJK30waIb381j/zuZ9soMaLTjTB
twIfMhCvei1cQqe3gB+B3+hpNDCv6TUdVWdYL+US9SD3upZhBdfXqgCJny7IdFhK
gfnDrMVd89UqHAbb0zuCy54YZGQCwdwxC1Jd2tEF/ng7tWUM7E7S2mzaSX67MsDT
dJb6v0juUsPXGeG7jkK9ClxzvjhjEpYs3LM7ckw6PSN7XCc1GgUka2TYEmheeJgi
A80C6Exjbq7lAmBqC4evHNw06ImmMPuTV5lXA9WD7BePX/nVPBNGW9zEmDZP+GIX
9XT/RZ2/sUKupS8AOAW2XN4VNUgNhJsceaJFKg7SsScrk+/Zc5xgXOiRD6NgX0pb
YA12sCXEb91oGuZ7nwCBFmDyPMxUQaRFUQ4DOiFGuBxZ/jFuJdbLPl4ApZoYvCQZ
oA63utsKAowY4kZ70RXho0xJiV/RaqGJLVnXMdcxX/EEl4G6/Ebuo6CwdAAHO1ok
nHuE/y4LL3ZkbUXizHQUgGb/m10gQrmLC8Vc2vFpp7iztCgMf9lf1huS5Ck+q7ri
Qf/QUrVwIGoQnflIz12FAciN5TBAr3dDS1IdGp6TUw1WbgJgAcrvY3+ta7Mh/xfJ
2aoMQ45ymI7wmlJ2PkhoD2HQG5wlWcX9r2iDk4KyFVqWekD9E0ctGMmBLpbhPaoo
1zD/IP/SDzCwdeMfGSoQECLn4FJWrxyV/4z2Qn5vy2M7lHxIFSj9vLi6CGp5/A/o
0WpfI/vxR5wEhA3H5WcCpg5AQfYvFEymhb+qzg7BKJnkDHx8Ur5IT8Wg7aZhJUeS
fLjnj8JuFnpcE5aqeSMiEgv632kxUA9n0q15WU+Gve1Vtj2XjcGRNC0VocAo1i4d
ReLk0F65hwNeh2dlufEn55bzjnqQzKnYIK8qwQQ2pLiwURRdKkbhiJgvAzfiWeIA
XVAYUb508xdkSmp7LKKQQscIKv2Ke4EkDkctjzgZ6PK1zGzuFAIEV0iQqXLNPp/X
og6Gng+IQ/ep5s5IK68Ujb6C9f7V5SXZe8sVxKerJUBoIhkjYHOTuLPdSwNFQlQ8
1Hc8hthi+o9JQJY4jDj0AOynnz9HS/0JysdfrEs69Rbkupmz39ZmhFPVNXgUXfI2
PhbdWsvlwJ5RmXiGxffz2Fj1wJTWJczD+N4wOLyoh5FTymIVVFr6mzQ28bz7WztK
UEN8MUhf0syGKZeNV2R7+yKVMMPyvtW61NYLnLw3yxt4KHAnsD3K0IsMNk86mN+r
6k7fzswLSnlu8CXeKIisdpxPool+5D0hjB1G8IRpyTqMiiU1/JEMBhQGV9w/cqdQ
ezwBEXSBlbFhMFSLafJOwJlb6bWGJFbK1q9QIisKl2QvX3SFC4Bg05IrdkXY90PX
4ff4Jit9NI1zjXKbaAeD6UFWGQ5FiiPFqq6IdW70VsIJSq/eumGELrnhflPxb2Tb
HKMthEszlDkbn8iXz/t/LOm145TmhyeyWU/oNOHfndjuDi4YUMMCCId/S3ArhnQ4
Q2UBXgIULWeAioR387G30PsDvNxpnY4BH+cCYGqcQpLGm/rUnCCi544YXsQKf5io
Zfg1Pr0SmbTpV39LN/VmiDA3ud3WRdhOMMix41h8C7YKYQKxW7DNjQNPl3hAphIc
bkd9Xn2hbqlKzYXTHbTNI3CYZWTdoniJlApHXAQhbemGmirnCZLU1F5rgK1UPtAo
varXPSX6inXOaLwGSIB2cfByzRlD8Xhft5LCeLfu0hIz4KqOidy6a0nujuccSIkG
8E+x+fTws1uSWYwJF6C9iFGIT3iyrXiLVvtLB6mN6OtAJdifIyyk3CVwcyk+z1rO
VFF0lkX7hCSGCf8CtIEBn+pVH6Gg5btpI0YFtzmDq/Qn0Bkl3t9YegW54xQ6wry+
lL1++YSQC7kSVhrY5GmT8L2gz0A320aQJBbeXsNSQ+RI7rZMtOWOqfITLkQGvxmd
rE8lZmwvSFdOyaqkPAvBXvGCHCnwkBPffew91gKabjsxrjXwHapWpYHqOnBcDf3l
1hu0UKwtHNQOl1U1buQ4iFRI4fGPxCRVtlZq+Im2F6t+nPB0BxJMiWlWzVnbEhlb
eXzJGkG0J6HF4g7O4fcD+1u/Dq8p8f9pHOAYtTaF/lN/vy2XzUZGh5P4mHcN8w78
2mqhNytcc1Ykd6PA1nWc5feUGT/lDLzaMkqvs84J8dPYfPkj0oNCpk5e3c09AJfl
H2LR83BPCOkIQKq1EV9Yj5knx76YYRX915VJnzg+BUk3T0V2YJhq4mJUKH5egC6C
G/6cciwAGMtBAKVc6b3QqCR0GnwfAYH7zi7rI2Gk5laQ9PTHBMTODzY2JIHz6Q18
wJm5s7x444oYykHPbCdTZ6CWngJCgDIg8L2p9emMWSPj5DV6XAI+HLPbmjwRyuIT
PMH2yC4F3XovVQCDAO7S4yvD3z721xr2k4P9jYCeRiH0AcNINdbu13wLVHpqREDt
D2I4DO9eGFzBVqow65VJ7Qx7ZRXuZfQRa6PLUYcrKrF+wzilYFFPCAiARQezy7Ah
lzmj6Qrfd2aqkhqv/r7/DGxz1qD1ZakuW1/+Z+87/bpTHIVncZK6m+bQPz6q2UbI
lb+k/NFijw03pOM0G3jX3o/+hj7IP5qfdsQodl3e17ESDXBAfQsUWQ0WinhBYtY0
YA9jV9aFxcGyKT7c2mpMqpJHrUzFG4+0RSLHELCfG/57Gx4gNXzKwNdJitVx9RUP
3Gop3y5ZidJ3NTgqI+igDAMeNBxwBRDz9aiRkWj9uYs6W+eD2QmTDAIWL6yDKkhe
7E6M1j+OIqsyFR9bXtMA0UrwH0xMD2b57ldENpShekCE303lYO22x5xmgCg+ah2w
LzHF9IN+jM1sh0M+udGsiWdH7HSi5DavEkdkOniooMxZ+zlULCdIhydiTnE62AzJ
4cuUmkDCN5k1e7boSSibGFtQMQhXbr+/Dknng5tut78QKxMPPjqJa/dLKEy+i+jA
2XeRo+CC+RT0HjBqUko1LpRV8owx2WXWIUzMJsS2fdr/osILMWWRaU3n1g7pExIL
9M5iNhIPwdD7Ki6kKJmKjRt1qHURo9Kd7nX7Wv7Z1ZufHfGc9Rua6iyocIzofus9
uU5NZUFLvliirJriaefaz4ELauG8jPybbRPQKtVamkHTr3eqR3htln0o+VXBXYmC
8j3MhBEQge5hwwqJMygmciD6TkGnUAACfy/pNjqKmfNG+DLYq3TDmE9RgxwZofjK
OGc8HIH5/hDGijv0qKqAjc0KxlOON25e5nS0bGt/t5zS81FbFpmRIQiTv2yTHEQD
utpbxkmJVp9CL478H4Vex4cxc9q0+5LDd7T8LxZu52cgof1jIy5kNzLdoEUhQ1K1
HAVjpjCa567t0RHxkdtPDb91MpDiPQI5ALZqGVCgKVPVjIabE+Gj8sa4Hh3lwVlZ
fd9MRrLpQrWvt6njoxxgiBuh/TWwV8BYHWvt/THNVXA2Q5p2gjZhJ6rlVvG2gEKH
XSBvdXo7E0r92W4dRWf7s8Poc/fDMZvLMNMBUKYErq7vKOig+A9bmHhxnoS/KdXa
+fWwQKqeCxVdi1NFH6SdXsBkmseWoc40ADVrgvKu7KikcrKoyZZNOs8a+nl/koG3
IdJAAyLRBNtONq1vGxdiVN8etXM6rHQQlFKA3W3+5QuOsVK0fmbqqp9S3CkqNhO7
HKFE47gyFu7/pHfD0X1Yjx4ZbZTWIAdGh62YLluosL1GddKBmICVEyX6STvR9lc9
f+GZHBgUf12AbmniSxCPGjXeonIwB6l/oY/zWBnsqhJyq9lCLROCa3AI7oQVZm9+
heE7XUIZF5zI5acP4dCzHb7okPWiwy2gJB/uVRHFVJU+eyp/4PPEcUmKM59YfL4W
l3NK4eO9C8ljBttPMXJyuu3Y21qcJJfxDKA/wyHtubXv6ySC2AlIS1K+aSyeoqEc
PlwM/XBsIQpyaGgZwe+ciAStPpLqkPcW1L8nTrSt5ss5u+104QgEY2o1vKDSyIOb
uBQNERT/KvHL4/bFRvcJE1yAix7quQ8ChfoGwaQyEC6gjuKGCUM3C6e4hKV8bMt4
aBYpXtZIs4mXGsO6raEGhVQLJYqONd6K3xmvOXUgWK2ASTByEJsn8rHGCXNBU5MF
3HvZf73lZjHrTQVD+Hl4patWGfxfWn51HgdLp05Fkr2ErgSCmLXPHEDLBFGhUt/M
AoxnRmJjY6Ahd0zMJz6Jdb16GVoPZ/0RndON4elIj0uX2YqbdLUbkZnnp3sV7dPP
BPApXtfVxGacQfSkWyIQ0/zUium0v6f+nBibvO/PMgVd9Irq3cdsGx400WFcL5Qt
lLo3IuKNFZf8wjWNEbwkpgDfZqBjCnkm3QML0OmMH1+WVtPH7ZbQBlWJ42eM4aet
vCFBNVnKgLsNrzPMr5bg0niwx4s+TJ/gDnccDa4tNQeELc36zcxDMv+DrVyRdXVq
f1bEXapecC0N91o2BfxAZbZFz3P34sx6WPH3gaVUmz1PgKzfBz+W2WV0DJ48tQ4B
HAvWRhoPaR2a241ZqnzYcvjjlJz7OBGnwlaMI37vb+drUnN4VFeF0NQUd5VhDgye
IljGvuVh58qcKKzMPbiyZqngSaCWxiz5QoON0DZ8NvpbgydlOjHDbVEM4zZ2cj5F
kRN4BTSDMP63ENHn/B8RKOUadNAcbjli9O7jMVnkASg9HoEi20AF4vLTVKVtFh4k
39xpALBHZ6Eq+uEC1UaIGwfdIPFSYojo2LHb8IS+FnCXJmoxS7f+vpr9pPCdnYhQ
KgbbHMxCZ1tOnZs0jvokjQoAAJ34EdSmLO+QllGzqkGWl5ObWjluS9vXIAilrhSt
RFWWe5XrPWKplWCpyy2rv/ej9IzxJh4qnr7TKHWYXw9rNKVljpbyjYi0uwcB4JRY
Yrf0yuK7LZex26U/HLjeNHmDDc1NXDyDcQxbopToKowl0ra7ik6xqBpoLWJzOkHJ
Rp0QYSuCDFPaiaos+LNjgY/88+JW5/SQpALOnzwExTwwqC63Dz+QgCZLqjCbChn0
3aqncN8Zs4kCmX/2bpBg9fR4WWdt9NXUtnHM0me2IuHShoWowzTsvEGKVI3p8epA
4vfIW6vBZFJ38d7ihkYa1x1PYOiM1TdW6wUu7RP899zn36NCBoE8rqupAiNeUwok
PpNaMU8L7UGD0QkGCu6aEroHAxJLEXA4FIWUeLvN9dyXT5YezFzy9YqM5n11pOI1
dMjX+DYVAi9lTML80ZpoMNcX5WzD2FSt/ecSchaHocLipB6OpJD7rHybfK91saz7
ilr/QUf9Kc8yMPTNc/9Ef+ATpC8iT7Dto3wqBhtdmz8B6aKc9OX5rSajvN9Ikopr
vxRjLl2wD9zOmwPxxoTt+ZsnC6FdfgdWGtFgTT2C5KI49aycDZWle9lvYc6RSCDf
A7wzXlKoSA2uC9FXdJLPh08AClNGiujtog/7MIbUdKjT45Yk1yp0xsCl5wZbYHTM
PVYGuoRi8O5W3ao+Ye4B0mtkGGi4MiWOKd5f3lxQNITDAXeqgR184ZANqRDhUdCo
6orHsFVCYVjC5EMOzRNFO0zLI6+b8uUX48Ur+e7KSCeud5qwPlmk4LgdJjAzyc4u
RWa8k4KS4B6XIv/+196fFWje/Mb0+l7i8TfDTNqykokwok+fMCiu+zfE0+xoCov/
DoBkN/M5sfKzJqA2u+mVeCF7uvhsdlPguRNFbEMA8qfNftec2J5HXxKDJNvO+6yL
9tjc91wfowBgUZJ3xT8HlU1VfI1jn8BeuoFrUth5S00eetSXyHkJrRfh24LuoyUW
P1NEtYLYm9eQTaNcdvA/eDOhnMpLc5tyz/ClpUcABshB8VChfOzg6eOSvWT5ijNS
4f/7eAdHJrAq1JrTEsqNoKbGSe6Th/ZW9xNcYV6QUffB+LrxwjyTalh7RKmxOcLT
eBdpGVbRYHRsagYhYToyCe5Qe2o9bsBRSC9u9xBexJMmQ9xCeFX39qvfY4slWc5H
/b9ji0WsqMNBUXEeQsxuuVWTiFyS9tEg/yYxX7LFZxW9nHsx5oweC12b025w9o6T
WWCwFRP8YILHFs/Sw+62V4XXZlJ86MRlitfOrY20nBsUBoXutv7n9seIaK/nNSFQ
7CEPj6WGEmojhuDiBwUsjEx2+T0XtDwK4/Atyo2D5TBbtpSihVEjh1xDK9a+AXIw
VKsn9LJFuyJ7xhByxqqqOW/ygELmMPQ04QgkUw9qzb6QmTYmYR8t/Wiy3tFD4fHD
ovAMrW//a+0hhz5n7viUcDz9f8yEYj9ZLuCr7ZOWJ5GiY4U+GpbD2YBaNLmKBwep
Eyl3U6IIgdLLT+8cY5jeyRG6Yscc/mz2uB1AxNCHkXsk/Yj2LAth/nDUZ+Bau/Bk
mK613XBaEZs+pUIFuLvmEqtY4xv35lhb2Q7YuE4HO26VgUovN18Z9xOJusei9Hdv
2G0hKh2KejN9H/y81gfJ7s/0wItS4L173d0UFTP5asnMyvAKQY/ebWf6GBSB6/dp
ysDS7YbBOPn5n3Ld8qX9NIt6qqP5YU59tPc9+T5Skl2ureE+SQyceZ91aVJO1oD4
o3A5HGdbygcdMxE/fs8UCMcIyhhzCwpQTfD2+1BldLuUCZtwrdxNuWNC4jND8Kdl
cQQrajGDC62Czxo4LUle9wYy+Qn2x8Ylv0JQ3M4T1/S4OEHqPQZYditg80MBv8WS
ouZJxEijYlDYuaKPn3ELw2NGEOkZqHeVlyFACuyCgOmvesqsI5OV6EpMPoYWzDip
sSAR0Fhka26aYG8e4RDTc9DJeI+1Xh2Vga+7DFJDR8WxC7jqcxE+fBKjjq7W0Ne2
8BqmtNwgDTGo5hsxhXCXR37qEjczBb5zPiIXb914N4DNdufzVFh42DetVAlsPE+1
P3cGZb0GMEGarBAl6tUE8Qo94sDy2Um4QxbqAP/n6XLaCXopH0U2PVTbSTw8o/Oc
TeiL8lD85yyYYKqhQuT1bvIxoVBRbIaKyI0/mN6K4Q8BxdSjXgzNNqb3JGm624Vo
s+4luaTXW9TgBT9cOeu14vYsbor9hTv4F1gUcCE4Nn7OhBsqjH7jCM4+WbufNIZ2
Dz8RLBXuR+WBxkhuzP8IRZ5U8SHnRWoLKjUZOufnTScYggcPmMCaDlQZOW8be/z0
x9TwNonRLu0RGQwZwTblKovR1aZ6ERiBGNUl4c+wWhm3ek7Khp/XPFJ1aht6Sn81
HCpXguMy/r4Xj0/KoY1/q5n6vUrtEUdOu2UK3lJbEa9TT9QaHdjVfFhVtiHU1EN/
hbqRH9STjQJBSt+iRLoz9PbF3o7iMmajWdlVjrDX/zRCljetEmlww2X3wwZ+elk7
LE9xyB/YjAxNbKogcX9N4TlzRF71HyKPiY9E3jFCJmaqCM//y4JP7+FZ7EQxqSoJ
BvI8kjszDGroEsltII1MtQ5ZTG3cU3N01cz5a5iat0ge6VPEuOacnESASQrMPDxZ
3NLeemcXKedtUE8zGOyGlx4KpQwpaO3X/dvcOXX0kk4MtJ9/tRHVzz/J2GpGN+k+
F6PgU+ZajUyjSDy06V2+2Yv+P7XaO82d+BBX723NlorBGwbZ3WlRgStZJLmlVnUN
qxm3JPA/gCPqK3ZcfhaytQZwVQ++M/jZnjzIHx5uIHdN0mZAq279TtMARQoswH2Z
0nkyrVGdHHqW50pwq94aw5CzjEEiq9VP+LQdIvdlsQiz71KnlM26frbi7sTxY1jc
c1kPtveWP1U7pE2iX7b/6gLfiYCuJkzo+LU9psK0Gz1kR7kMQQJIgk/gNAs7xEj5
tQ/zPlXc6mHB/LofS6GqNBsoxVLjueG+tJTWf08Ne+V3XFy/x6sgShNwj5VyV7Mo
quoqTS30CJpYW8PIF/wfxEe1jsfaII12EFjr9LHo4WL72an/Rgr2CFBiW2cPHcNJ
5KlebouL+ONWOVu59HMpDnr5OV0hybtX6b5fwXIt77cwqv4KCAaGTV1RmgSDd97k
Uu3L8jfvDh8fr7yHhG4my4iNjFJ9rMfS5bXp26VLAmXzdftBPMDy6aBUsPYmEPa4
14lrQQEzTDFogQWREEnrhakgNYy1B61/4LFVPeehs66DJ8fQ4CkFRYxx9FhUXqWI
h0T+Bcp6D0ri8fsEF+jIwnQXlaP968KUA0xbhqeUmCurOwLnI0UphSxb35hJFsGs
wcAKL4/WHdobOCnNOdTggL60DZ9Trq7ORw34AmROnqjvc1pXiP+gmaxAlii4Thmx
g9HH+GVShQBN4YSSOKbLK0HRceRaB+RdN38XHIElFoABLS2xmKU/x9z5Xqt0RqKZ
7SMFHilMVFtwDJTVP/jIUJ0xCrf6BMGAyrZ1Lwv2VCJIFmU9MwVLmEwOBWQsy/Mo
s/uTcB6p9C0fg62KvEaicFtTDPi38/kUm+vqz0zzyky+nJTTlGbODroqQKXbniWa
HNxx+lGg9FY1jrGrkpuPmvJIpUKMYWr9wEP0MWK++UCGEmVOWA6Qqp0+vQNiL3/I
S1bl5IfrZfgUOGn553O1LCGlzhtazygEMR/CuI8QgLYYE3zLTVpnlAgXhJUPmEta
OVLmN6H1SeQ4syvRCsKvuQ5qcYH3GDRo6oXmv6d4CmltJyEZFcBq+GbGJ16E5XwZ
VhBlzKoyCcrjrSfg8J7oRwLJSaIr4hXNJJkXKU6kxJiw9/U6NWzl64tFwZ740IZt
8n48B5u84enp0IUWU/bo3kUaHWL6Ne+UPxe9Jao66XffyhrarOYr1FtHpCK+rFB9
DK8Jf61tOpyt0pfkLEABDCiRMZIqqcpJoGVVwMCRfiQsshZXWjnJ7uHdhjlDmsgo
gBZrZU1lI683wsJLzmkHcGHF7itLArLehF9IuVM32/UhfH7OXU6lYsn+8YZTXMhu
hJvDtgqNPvH0ODMcEyGHaJMuZPosf7z5qA2i3Tul5xAm3IemN/ZUpOQLwfoMT6xO
tfpaXl7cgXF9Dd1Yd/6ZgkzVKzOqaCN7YHD9Zv34GrBZwMvJasJkrxa8ffHSp+ZQ
1yOyBKAD9Yao0QVr5LEbjpEv/+/ggezg5hVNiQcosgpQjGufpUHtg8R7JY6bgAOO
cvPIFZOSO9scnyODdUqVY4EDQRIGwrh9TGI40tBal0gDIcYiWHvysepw4WdHhWTN
bjr3JkRTbCN2DVfChcuIy6bmVeYI/Pmi7+hR9MobHbh0A2gUNuAPX1i3FxhnX0Cu
EUlIWGZQ5S9SeFZxMbcDTkupjgnMNLtBql1dJeJFjTeKposznXqmyb/NGfZbPV5n
jSgVQ5SR1OrhWYW4DfnpBD6jJt3OpCDHAQlkQeQ2fVu8w/LLEaqViCAWSd12oWlQ
ieJSlwmkPveFgkamvL408sB2s/1wkZpSeaMyHsfNUMeloyGFHSCgaK4GQTxcdFyF
V8HsHnrZ5mW2diXgbtnkvGVWuzaya29s/jZs3sXdflRzuhsz6FXczBdsRCb2WRZB
mcX2GHnv17bu2tHbYSEDOo9HVAettlYpmlBwIgfZJp8LzfIcWfUGMfNZMNbAC9zQ
iSSKt4moZnpKGAQ0HC7hWVJdvth+c61uYMPoniaI7dL4t/FNrL+hDt1aKJhL+8FR
jtzcXZbVO5XNZO3YcQ5uaQWWrRzKIf+PrvLlgP5/QZwKGMlre7KIUVQPNq2lED/E
8TJkiKdexlDQ5Iyf/dVh5yEkDykc4Hm7BxRCVHe4TSNOROMPxjvROww2B/FZGEwa
ZKvlYbS4hyxJ3gBGn6oXQYIsPUwTur25eNtncG8+f1CXSf1gzwu9RxOnWJazA8PX
QUm8NO21fKDNpjRJtyfyjUSmn4likrNBiv6LLRUC31xftSroO15yLDOo49MjoorH
WYWX1W6Du5jUucon+RYFEM7Y9SVRmIN70pCz5T6RiEx2kiulZahBpi50eSGQCz1Y
3fmOBBrntl11trZeHw+buWtO8GUrkSojdetSjTr2qfbgOQ2uDeCp8F70/L2WmXXd
3tbrR8MRS4iZimC96JOQZG4ZYaDiuZ7xH11fOgloNE232lVc4sYie12+txlx3alK
2eEp/C9aayLNXTKs0/frcHuu1fQrZjVol/pJ7EE8G1NlU/Gkhnzvr8GIUoGdgNJq
sefbqae+N2uKOD1iwbicc6uC3htAOuYIarXsJq6XWNYED1xnLnJGvc4dHTQFkCOt
eDnBoImg5UYMFQukoB/hzXoN2lYORZI+bZ6Ttq7a0pvGwwRlBvEBt7ABhfctNgfg
1WZstd1QfwEDfIe2gk9M/TgFxXsmYtWpg2sRtPfSgCIs83SbkpcNCayKcHuK/eCU
bO4dyfP//g508eDsr/MTpZRM+aYV5zPqH1RzkmhPE2NcifU8XvlG0tSYP2lfae+H
g4RkXEtj8Cxvh2nFr6bHbrkSNusUR4g3LauOzxXu2XuMUvPx1ria1EGRZ0MW01fh
df9GVK3nGNdI0PHwWy+QO63upDSwVN8SFA7FeL73sBjLI4oYLbDvwDzcybbjY+0t
3vDizZHbcTxJTTDrgLMSxQ/icNh1BQbsElUoSZgElrQ/tIvuNhkfDwPTcjHeT1xQ
kfdzPYiUw3zsgBHkRbTKuiuck/alBtvIeDzZ8EjiJHW4lpCtW5fiQmlCIH4DiHTb
kSFw9dHgavJQvZcBPl86i05pH7MQxgpD+c2oZvdaE+3DhFBUSoc9ITsFUUc1EC9I
w7r5HAjDU+okDL9PzFu2j7YggtGvl3DNJ7nrNY5qLM3yZyo3h/h+uXGh4Pwqmwbw
7hrhMQ9yacNF3ffpmYN/icTVxAhTTkOhtDoRV2ZhHLxSiFKVXqyWvjoBx0pu26HT
K1V0HFFwkFmEt1/+WeFCX77GcnYL9dGzM7tlu8KFBCL1daNQH/FSqt3fP4C7Uo48
sn4zrDwkWsFfZwOv820Wbb6wXD9sAvQWVbXPsnO33RrgqL1XVnOovBDHTgHMwEJB
c6CQb5Jw166rwY0Ug5D5bubpak4O6lVV8Yylw4fzzqF2TxjhN+OhFYaQ2HX/MWHv
oIJanDE0iYPwBYA5+3rWLNDLsR5+0zKpu2+teHDkov1deylonGUJE05KRuG42YQ1
ma+oaY6+rqh+KdN2rDkByYT0cOPTRVPQyGuKx9+84d36CMPqMDyQh3Pi6ANNL0EF
RjZhtu0h2XmjeVQABX68I/5Yraa3gRVQqn7kr6P9QzlipFhZA5nDdffAULtUhXhm
1aodyi+oc+YXSchabpMj842Y8YyfRDvJ8JdQrHt6OScfRyTxgDjVd3AyO48WK+ux
O7JNtPzD+0KDDRGdSgbaZ+VDP52wi0m822V8xzWLkSloGWmjMk1UEjHYF+yK/a2E
78rX8LeHGBcA0w/O8M5k9pIS0U98MYOvabUM9ZhxQZ67++MTMC2jmsBrUUcLvetj
UPEDsGR59wRTpICGdqL2boBjrjpiIsEpIDMLv+79y3bzLTbpvpGHYSz+oxYaF3wj
8u37EWlmP9A8ISej8bHnlfNVUBvfizgXeWHxCvzPiin7wmz8lhxRY02bLuDK4YEt
d99qOT8p0ywEtZXAr47HEQuDio1gVr/w7oJbWtVma1U/1U6sgWbE4xEgTgM76T61
zm8cEsvZ2Hhyt5UDJ/rbuRQ3IvLk+teKthvTREqPU/zAWB12gmuHkGsvD8vSLGv8
jSr5Vjnngc3pKN/yRw548LPymcHQ8W4qSVsdhrqU28gBKMhp4nwaFrQmvotBlRI4
TBwxvDSdSRPdcoQ6my+PpZTVkdgTbcOo8V1JDPzG1Z4p5OG5G/KnWM+cMxq9fH9X
3/QtePySg+GoRkqmQzP+jXhcNhzY+MZJcJ5jL8y2NOPzRoAlseAB4fqDFlY0zgJi
6VrCxdhwFbJ2cQHkH9bmesr+ZgmPNMO0rjy5M2HF1YdNxw2OVh7bClkzaqIDARhu
8XT7zkgQLrVmYvAaqhqXjglrLGOSmJEZuIZgBYtsnifMv9xQ7pLISCTDk4Oqqw5w
3/ESztAdn3SiR/V2yxHmr2iYzYoJf20mNMGxyw4sqrPjEwI9ZBJdLDww05HHmG0d
4JAnQm4S2w8a/Ur6luGttp0qKdA7uaNZpmL7uNB2rGQ7kwSWMul+2Zg3traaRqGA
ufPKk8j/RnRjwY2nN5N6gIK8D8ju45z9VXIsYhTRxi1ZZiiL16fywirWMhiSi2P0
og91ELGk50ZhhxYyEZ1w9xh/DjBkX1rkqCx83azHjuRNELv3YlGA2c3/nBvUuVzO
yKB04UQDmAmOCMtvTqxZ0pxjSTQocl5uCVxARK2DtAKx64b8Mt85b6Epk7ch9Fhi
VSkT0N3vhnLFEB599W8NT7YKltIiZaHOHocb+SQPd/P7cwv2Bzxgk192E/t9tmDI
qMIh4JjHxcJgIamtFLcxvv7SW8FziGFJQri0Yn/7XgyaMYEhUs48Ewqu0+tQ7Mua
HyajI7ULKTb43MisPxaBsWY04MT8WFgmaEBIokxkMRNT9mID4ARkE4EsiAjVYhFW
CrjruH1ChyKkC/svqG4H9KBwhjgeaHPsfdDRokvKOxL3ctW824x92cVTyafos4e+
82CKxDvzoDYMtfiK7DBYkPgS17W2o0mCPL8AHhgt2NrxtVB8skFDX+cCzJrBywwI
QU/93OPw7H8AXW0PE6kFfqazd/+Kquj7JLAJnhRMHDDgUAvrgj9xGuOG0o7GZ0fx
1w+OnAW8QBC+ctP/gXUsdoVnRUXlHpqWkuHdaMfFhLyNdxKFYW3Z9FyWQrMnLMRP
npNVHGBAZEaa+5az8GJSJPPeGUdt0LZDyPcuUwQui1S2D0YhctMX3xRFX4/bEFI3
LWXYct4G4iJXDvmW4mfahhBqbvQs/L8NazyUIC190vmhwTf1sWfVW2zVN7O0z+rB
f2EwZoml7Ho82qOvXFL9xF7g3BfFDQBiVY3BjdjygLzLAHR1mBEa3vDKfdpxk/xI
EzlPPoZ+30UbvHJ1pTB8gQyrujDwDtywAVCgv6RPAeUIpAEfwKYGal1SJUhvomMM
Odi8ghSbIWPcYveK2Q6QLE+Cn3pan4gabgtt8li+5sVk0NSIjc0WDvss1B+7IjjE
9e+kqS8gOPIxZw97CjSboR7HlauIyVBH9KMjTuZy0zDzfYuVKNxc9r8yzYRzBq8F
kOr0yH+p0J74eyPgxttA9vMKZoPnAJ84BBNm3NcONjBY0QuRVmQEtp3dVw7kYS+l
E6IILPOqOW6Uj66Y1f28hw2V3Kge3hp6w9JLtMqI2+1YZ2IGtW0L0sZOrUj8jxja
iULU2oEPljXOMyz6nAaVwwC3mcJ1ddpuANF63DDBciaZHs+dZ8Yw23sNp6mTvLuP
3AunpLQPJR51NHpIt/VRriQ/zODCUAFVsfzSGZjMSYJdboHApHmcLbiKYzv+wXDW
HwL2s9EASM21QKCstpTkwyq9gTTkWi6jO4WMBjT7zdn3gQj+LeKekLOS8N0zpnLO
qi53LnwM6ga1uX/q8r2qzvLFZacUmaNOrtmvwWNjFzJTT9+gWpsaVH2sCKjWhZtJ
0zzFhSH4Agh0e+ppAagFkdJaf+bbx6ubmWSycWrx6MWLmlhNkiZQUw8WnkC3UF8O
PmNSkNq9BYw/opxt2XimAvw4BUQ/sQ2CZ2dhj6olkiwSBjHhFEKuZtpCKgmG+LZV
4mZOdZxBiua1OsUzvxvNPz2e1kezKODdtS9yyoaVjJAoi0PzbGFZ7is+jMOU+Ift
aNL3B+2UAqb0YpCaEVxshX8SxbMQGrSxyXAImdLLk0k4pqQPD+LModWGTI0LSkQH
UrsVzviRwzHzI2a+25Lj/zI5vPLQ0T1TqjbDzijmu2G1cs3J5kAKCHAudUpcZjlf
tj0rZxAazz4j7qGwtCJgCSCw8ELBdlGw3TboN5v1TG4zh69xVeT7SsnMDs0rTHi/
ijZulchrXjePt3+70NCGnCBg7PV8HKdvRKNng0XroV0ZZQVe81iKai0N2j0nhqg6
sqTOunjJRXIc+tLX+kiPDt2JSkAx4ppTMUsF7D6g3m8cJkzFrCB5uf+WNmHN7osN
/r8uZfj7Xa8zVtGhmRvLMjM0LBNsaepjsm7dMS20/KCjQw/TvEx9RdADC5coar4A
W/+ZxuQfKflzi/LZdssf1fh41DdovpNJxSpJSUghokOtnYsPDjA8yilqyUIl9ies
/wP8eUbe2AA05I5ukYGikI830sHcXFCiegrbocoOcBGremeNlWs11v8fuX4sJ1Po
dYIjfyR8fth+EPHML3VQdKF3V3AmTZhvxF8HaXHBJ6kWXi+7MY1ysscy/Oa38T/I
F07ZBhyvmy/Nd+OanhaI0BRkA3yfjqaumqOSH8PKJ2KqPgN55ArzgYUTgilMZB6O
EKV5taOyqi3rx3zJEC/OE33u4y8rBCAYibYct3SF4DTyQP0FH724sQ6QlexWfWiQ
pv14lG+Ti6Pdf0HFzz1TlZBj1eaz03Oz1vFdWT7MkB7QAa6sLO+DpSudJz1aMW6A
9ZYJG+HjUCsvhUgCXf3l8yGgi5z+kdX9Jm9ou4XS487VBmyKAgPNNAGiUzIaRNV3
HutXjE644liLFsr7mpZK3PkeRJUhE4KfBjyiF7heZShQ4CiBY4Cgr9b0HgVpv6nF
UrnSoPM9tPr3BQoNg/lmWHsHCkROU2gDNoCbSnL4Ri6sMvpUwE3ds9nbnq/U8jIQ
lsfcxrGmWqc3Ba44nQ4fvpGk5hvYq6r6LzanKyC+zpzYieqAv8kpj+HtZFnlj4fY
VYEcO2Q/wWYqzAsMnLiIwxR67awVmYSdZ9mwBI9boefDwSeVzyqxHYcr1/P3FnFl
XWZU6WRt+YBa1P1janoKNyuftcFj+yzOHY5khyGzY69spNmv4/QufDwR+S9fNPq9
5Zs0vGn3alHwe8qvU1lji+0HLRRpykQiobHfuZXRybZZdu26p0TtQmfHUuk07vDP
siEp2f8uwWdO3dk0Pc9n9/DesI6fHLl4WL7Tta7eyyImrguIS0YJZ/lUQ1+jNady
cQFm+EoexNuSopRbutN7xH/loT6KLFm5bLo1nsmGfpHQYjuysHLotyx8Cmmcy91a
YAJzUTHSL9QXWEPJl+nRDZRKV3IRUwORMOsBWdq7vHsU8TddHXyYyPGNcV4ESCNG
JC784roovfREZTREwUnJBrJ7fB53NfKxLpt5Mn+yBFz3Tp/cenecrbB0wr4FFQlK
osmDYc8wgXx7k8AWoXWqq+tPIjVOJo5Fg2M0yCy2APfTmpA03zZWb+OBIZ5YWGUY
JfqoXGvFye2CDaC40MM6DwqZogNY26u9ylc2HIYxR23glvsjCny04zNWK7AJhrFT
GQjq+uoAuoifCfJFrn2yOfijJ0OUvxVsX20Dm0AwyAIkacWfqqTeYSW8FKlN2nVE
Y+Z2kQYxC63o3B2jJM7XmC4yrUcx7mD/9BuDfLm3F9UWCQYw/Bh8Lqer94b/G7D2
GNaakF20HA0D2omxbpj42lHjD+HtUZIlUWPG6eW9cuewhAaaW0Cv76+wnUgmjTqJ
BPSoy0o1j/DSiVAF5gBAfCUv4nqRYfUudBtvqORck4Bdy0MAIjAngP5AGFzz/wRE
Uh3+Z1L/shOFIpQia+6NcAz6j77OuXSBT4o03H+uzG5xD/oARZFPnQf+qqH/Hi2B
hb+ISk5h+qOjRA7VnbpoNt0PIOiHNCVYED4JyeU3RaMZo0V7L/ILOCq+6/G+it7K
swr/X+mFQ/P9hGxDB5CsVdAAVYNG/tDIjPf6FukhDMWTCyiiuXou6qbc2TEFoP7L
vf4HQExhvJJAj79URllppjfYloXTdvZsGoUcK5GcRe4tMp+8RUQMv0Z7uJQ61aLV
1FLxsomg41h20w1Eab5WbF/E7va7gkV/BSALELs1dQtHJkNUabSoJf9nu0eKyEns
ueKZJggR19ecrMHLnGzWRH6xgdNxbfyx07h8d/JuwQVb2Mh4ZnPpyEBvyKmzyZ4I
dnSqyXcSPFFW/0AtA/c9UFWmqwPclvyrIqW9SsOvZD9M1dh/ACnBNXqSjnBnT6sz
rdWfOQpfRwmB1EZ6ll2/lLYFEYLF+PUoDYwwvflnd3W2s+6NmLebXveLQCKPP6sS
swK7dWxkyqPdyG7+pKstKKd9p5XArT0W5oVhscmDeDEoTlpI02gfticiIZVFq+gp
Q9744FNglXZOQSb214w7BmYes+D7hvcisQhsz96jf84+XprGgAr11xOpEhNZ2WtV
kDDDmEIJ+2qgPg2q+V/CwGVU61HdzMQTLpCoGe5TmwuQtJ3guebJzsnN2kWgMsle
59VW2L0w2dcUdx7MLC4WCbGLcpt2/TSZr9FtWCfzp76UOnKm0OCXTmr/NF7VxK2l
4EcYTSjJAjtdw1MZWgobPE10e+pzA/YXyCplRKznpRItsBnzasiufnXYNIc1nrdc
2t4VnkebI8tuaujG+csh5jgKIk/k9Lj+Gs2mSRFcj+UgBQVaaEncm5XihwCEV/U+
x8W/EPIHbscRp8FT181Pi5rRTJafRRQ0kLV5Gk6ATAh1XHCpVpc05mdeWUWSGSN+
nX52WfXtILQyXs5xU0hdISjKnHdBF67H/wcU7NrGv0e5NY6aaRa3kpWCHov7pJqi
OeO7vCedncYGdS1r21c9DWS4ykRRbjxNL/25LTprRnpMY8cvr6850Q6W3EGOUbib
flPoGA3EQ75ZYOtC7iKi7Ezp3VNkqZDY5DbPLpYRoyQmIu8/GcwaBPSbU7LbtH/z
DqDxDz/oO3L0MqW7RXyDTJnigswywi6M1lHrlsJRvww8ch7J1mXsG5wrTKa/8IFm
wWOLDnstGXn7GfFrTfpUMG3HIiJ56vwD5KrZJQy0bamLah9SWwnzuBgq2sSXQ2bP
myBsA/0Y7TViUiL6e0DWbI5nkJWdqoEMMwllOeaapAQS4OpdHKkfj2uWuf1QYNI8
gLqAdOHLKG4U/xr5aBzd2ZJN83SQfz+8ko7lhEwqkN4luDPNsdJm0R6ACOMNstTv
+Z1mtMBokGwqTk5ItDpA2rObNgbvOr+G//OVEJbtRazq68jMhROTBb4Pl/H+mALw
4qlaewPZCfhSu36+Az34kLVZd4/Kv5Oua2dQyaM0iBBbbGpJliro8DTcKuh7SYV1
daH/TU2Lp0c7+HQ+jGlAPMl/8KQ9thqVAc2B+eic2jP1ZVsaqltjMydbtEhN+smv
sJHYGZhiGgEA71j23AXVn9lL/5+N7NW+1DivR/M3WmRUK3VEvpqLp3ezGqkJSWhq
8301JM3vUuDK4CRzo9Fb0YMbchKGk3ZFtYyw36Vjh5/dSK2FcCl7bnFEOZSaIwuO
9wSfpmvYy2EswhSBbVVrPKNFIz+/mzcV9iYiC9WB7R79pthWChioMx7X1TZywRrh
YaZbVCZZqN/NeGwjfvkavMI9Cds+ofd+Zdv4bXpIyfakvwFTl4tAGkUuHCQxgNH4
Tg3VHUQLXdF0rxlBXeTvv78Vy63eq2Q8XhDuaQkyh/zbjmDNvmIANw+sXDc7UPoo
S2vNwYuwxyvA5H2LnFOQMhoc0Dr8dETq5b1L4qYh7jXX1uSDsS+A+EdhWC889Yla
+sKlnhhptP5HPosln1tyG9mFjFFyECWKcp1Qh1d0jUa0A0715g8gZ9AXoFEblniT
MYcHdOdZoPqN9aujha1ATmtb2fBxb/YIQ7VdmZBqkH0oEDmOpCg1Cyl5goxl2ZQ7
7QzhLCI4CbDqb00RY93HJ4oMSrim9wn2e0jDG4FyBJvYBJtubIUZZiXTO3ZEKzWV
ZrQvD5Y3rfsYo+1UuGy4b36S0E67CZvQPdSLG7CMo4vZa9t95HWruCEHQKyVHcqX
ZXBgpwOknPEfEm5ENfEu1puTjXCVu88tEBRDVQzni97QLJZQ2aa/1GuDTUb7mAP2
K1io6znHEnGuSzkRCO0Kewdf2MwF6/eOPIf4cxKjMRh3DMkP7/w84EwJqhvBl2ad
hKJ6YOlishsJeleXd9nz1ht9nQ8u3QGKbsl49WYs3kXKB3wfj4D2h9qk0EmF51MZ
b4NSLnBKt+nQ3Is/AC1veOg/7ZK+FrP+nnIolN8xC6xlMHoEQtgIz25IM8gJFwbZ
PQVyZmTlFj6WSwHkgIPGe8H54BkdtkJ/LMMZcjJAV1z4ActVdon/CXTvUqGCWyeU
fvjJZz9lroJyFjpp6bidubXjbua0QU7dAItWm9aCrOkVSKZC0XzkMDgWmW8wH2il
UtnlkDP+s79x+U5iBQp9eS6nKjPxVRX90nyMnMSDgaMlDjW0RbNl6eAlZpNatlnH
2M/M9dKt7vrPYdXrrHdYEGFNoa2rPv150btPtQmc4rBpSKtq7eu48ARlIgwZ7XgT
NxIo3Edy0+TyrPWqRAOqQJKqvGbMIM2qIS5/ptMPdn9U0QaKIhlSKUjBjEzV3XTD
whzOXvcwHZPEdisFYoxuHd6gXndFPR9lu4+tvf5I8/41DW99kNHqD+IQGSAqDMzh
VBjltwFnNdmX82KdkWzcytdrJDPEKlx9E0L0DumugQ1vPOcmRJL2hp4E9XUWj1MI
8T7UjwouTXHyPPsmHQ6NVJARRD5qbzOJk+U3r66rhfZ4qG5GGeQNn91Co+09oL5o
5Z5qiCNnt8CY26abPanBYoIfc3rU6cYax5Mp2efJ3FnbylJ5DQsZ0kTiIcrXzAdm
r8CxrDftrKjoMDVOGn5xtfn/mXEVskDX4sUUOxj0qmRsb7dALVNTzhBq6Wx4tYPu
65kcdZtAK9RK2z4/NI1zyziMVAZf38qmkHDuq1FXGZIsiJxv+0QRycKyCQ6TNt5J
dbz5r17NfZTYB6+qwjA1MoGutGtqyKhHkT8Dvly0tYQ66wrvKHYYmfbPnlEfc/6Q
Yyxwjr6sr0x9N1EeFHyAnnv8l+O/xJUmeoIoUY0qrzf75cs2eDYzvYiGKeDsymuJ
UjVWa5mghsDAZnchQGooeBKdeqbNWMEOeosR0Mmqelel+YL//1LhQcKOSJ4viu3R
aDYcZuMZ3hAy5s8EfDSQ1lcVcFXj0XnYTogoUIojzI2IXKNAF1pTGaJi15Dn5eJx
mel/MnUsjQm5HSBZHpmtKLSVkM6vb18vzH+FIIu4ii4pngs8hKh4PPrspq4kfu7r
eWJ0OI21yzLsXGOIVwrgFjMcui/Lo2/78Q1G9imE1E2J+d2cTab0iNoZEQTb606Z
6qKVddVEZjdwQ+Fo3RZ3EuIXGIzAgOPzvPDlnXQo91tOtXTHsPtnDZ6qRVdbQnK+
/ewr1NF/yxN0YtmxhWHX6iSv2+pSzNUEEDfsUHbsUysZazO0qUpNKEx1Vu7h9RA6
gQgvhTFj7ul5LptzEh2oAixOPqbT4Aae4/GW0iFvErAMqBL4yLV1UkxJ892IYEDH
inS2QVq3yYMpel3cxp+MRMEQX4U8kUcODz3kig7YZbpCrXkAbqrYB9kjD51YDpnv
VZ1bFIZDIEFD0cq+U+oar3wyfwjEvYyaHx4USDudjJjpgO40vlEt3o/G9Prl/THj
21BFNJ0vrdLaFMYvIDDz4e+bVA3uNk59lozr/a+6lmWh4NwTYJsl4GI/MKg6XTam
+s+xx+LeOkWZQnsOMKb2wgRuAQKa4qdlyUZxwY1fn3ZLIVcicQ9h8Uei1VHz3z3s
Peqg6mTodaXOpM9PosRmKTrAo1VFxpAaAIWgeS9J7Sg7QYCU3YIS9fhPkJ+cf/C1
rWUoaVBfGfubkhn78gLWKXCXQQPOxPPxXUZQmUNe5tki1KkL0Wl/SCC+brRUs+Zw
kM0ElPK6SBR1CezhYYPHHY8vGwengzIvtXB0DuTnIn09jcr/Vo7sjH23ZttcxJFR
0ki8vKlZJFW+zJxOzpJPCDSdLDRgaLAChiD0B7mDyRqaFcfq2rjxNOoKKMoT+XyX
IfOcMi5WZ6piM8F6a5gY0L6RRYr86zfYQpr6UsfmHsY6Q3DJF1IODrHDiQ9/6Yx0
+2aWkbsgejiDvMlturgrsZ0ReIJMZGDy1+T5NcY9hysSeCsOBr9BkHzcWh56X80N
RMAugjfQYhePVZK0VcZ7VS7iETU1aKVfHuAYwtGJ93eJ4VwaF5HZlGdjlueLBjTT
i6zB7tq5IEORN8ZjDZwk9vShPT1QwQ3dnRxsxJCt7VEmM8EFT0VRbFHVJuNUzCqI
Fwvdy8KLI47GJC7qNTe5rioAaafeQsCvBFgcZQ6Xipp3/h5mf0SgLYo0Wao6byAz
+80Kpqc8SzpLnAPaMDcVEKmx0zWm3pcSik8o2C6t/TZJplG1EazucvSUKsBPZwIN
U4dGEXRNwV4z6MBTLsac9PNy5HGqKJhUAY/HHC1YeaJ2CpsECyjzZ0ThO1grj/Ot
DO8qKhMxuznHU9dVRjCasH3QlXQ1+CT4nvqjYKxrFrVOkcYvfSktIhpzxr8zZg+k
S7sZB4DXkx9lt/VFFvTD8kVebRncO6dMnFwSefXd6Cn6ChpXxmXNO3VDQRqL7afj
XECT8lXJjkWWtay0bq4eJ8FG3aa80iNMy5egpu7z6wgAbxTQG5Q0xabmN8OiXdeU
7JOR2mbOVwVMlcNP7dUw/AlaQ1xX+z+KaSoUg0+iONECYFUOvOOIzCvLKmcKmt9B
Si9VF+a9QcHANwuOE7wpUxUDCUQoYNARc2WGpq4xhDs6cjpqwIgTaJMYaUfIbSiT
CS9SRuR+olv8TEwqminTXlmIhKAJRBhFkGR5ZP6aKUmIKWCqTR/JzZ++kfF2DXTA
vpdgWeaTUxE1F0XO/hSGunsCQDcp8j45rlsJuJQ0MV8sAm8bOTiDZF/peYEEmpVd
SDfpALuPwWwQ+h1TYCee3rqt68qYdBBjMCQ5F5TOBMQaOJpsuvFYa25sQYkXGHly
JWTDmYZp5Sar8n7wOeqSWTWZfD0ZRu/E2ch7MKx0nwir49JhcB07T+BF9eHrRHFb
FVnlebfIBKY8edV/YZw2tNbsB2dPlI2tvL8g9o0a/U3FsU4pPO6nO8uO15CRGZMe
k9pz23j4AfmNUn+VvuX5Ejlexze9IHVjOFhaOtEMYuMN+7Up+qD80yTYiQ/Z+u0m
ut1cfTL5G34bZ0C4VXyYDatwLSvl4Msfop5A2ac9/Mk6A+/4j8aDtRSwu2jyF9Qn
yjsKRd0mpxTutjkLVyFhfRU/1fnvfwwnIprKfQqfpjEwUtIufEpc44mQ771VKIQz
oxQB9YL3W049UiY2hnYNLNkH4gzdL76+il+PMP+aXSV+a4nypI/Y3rv3UFqrRZoB
XaRrZ+NOEC0TgD1xzkrDNkiSN8tulTXHl/JpYVtwGrDUEpUQfP5pl7AAnZQrIHOC
i1C8eUIFfrB2M39VF7TJirpvGXOqqLpDEkiEn5zchknpD+DF2a1FJ1baulBf6YxC
BTeWwQt/Mh2g3uYslpeknIkn6rIQ4hFgtLzIdTVPIkO7+Row+pJNrT6EbkOzV0T3
Zm86sL7DcEVx7Oq1j1OdGwoBxkVO8zMEIMXya1Oq+oGZ8eF1nnhuj0ML3035JKmv
V6gJUrhu9hkXP48ZPL9VKCfyQqC3QC8oqdj161jYN8pATS/zIY4i5dCROge8Awpl
BjYYvSTLPCnJ/XZ85kgc3dwLEusD6r3RJPVIr/d8qAywkHiVkgtAwMLyt4oYDzVd
ljhouPA7yKof1R6cZiGgMVCXqRY5wCQZ9SyUMDZItgNctX87BqdKZF3gsnXVinWl
j6tnH+atYyQ518GOTM7Gnc5i1L4dOFTHdQrYRI/PkCFNiOCE8OATIMoQ4gUl6iPz
7vXK6bmhG/2NVjXiqFKli8FohA+ORA+rO7q4URB5sFmCWtbh9i1ZbP6kkYJQ9nTL
vBHfDY/hIuGpj/avOGyw/PBYfzWvJWzld8klMCFlLadpPELacllYsvDBM1bxq61i
iRDtCDTnRnK5D4P9464EYGQJAKUHNQhpS7wIbHhJIjo4U0tLk0OnPOFxLesSCpqG
h803qjgAIgiymBkDJfJEgr+M8gXuTQ8V9g5UAVtHI7smE2G9N2rLkd+dpPty2IUH
e86uwefucIR0btRyg71LkI+V03HlBpNQrkpPIjsyh117K+R71dDr42uc8AYiuFJp
M7l+50kjPEczSdQcSWy3glEno49mbCIfQbHCD0Vq0xD0BNNFePOO67fnm49JzIUh
wNBdmqfI9GHukevHO57ZQNn+XF4n2qnbAO1+O6OAseMfzEtCFbsPseGYooL3yYlN
MrHGAZmJm3quLyp1O0D49o6wcoCJpa/5+zxG7dBijgEGEqynaACA1vISRWvXR0Ll
MGljmZ9Q3numGu5R/SshcHOLNutVetV2YYz4ijZABiSUOLJaJbbAghjMvFHPMKRK
imOo+sOl425WXqJLnmw8pgZcTtWTJq0c1Gv0B+eM/wCzRNplbNUFVzC6GkK9dKM3
bpROhosaIr+yLx+eODttmQENNJQXG5vf5gl74oCa/vfc+pDPmyVtE3sOVdcXVVIU
xUUO4wVPicZbDF5UQeWT2JW7EBsrZkUFlutaF0dbB+r3udCrqNhP8j2aoxK5+8jc
YC7VTM3jg3RW2Y1u7ee0hy1rDCv0wn+Np9CoZRpY+tcP+uqZtEgaDMnio/eO3CFu
gSBUO3/MQm8Av7ibxcFuL9ZefZekwUGKppNCdjCxubpieGs9C+aKTbpCgZme3toB
JZleBGN7r2Lz/ts6qzyr9gZw1qIodzd948B6kuZcARarX++mlxmvO9XRCPiqsoc6
BMNxKXOisgIW/CWj3lZZaj5pfAsuUX/gnNSm5gLpkaELt5iG7Rq9ulcu+N+5TQTz
qOKL8/7oVNALX2ip1CsUnej0qxdLtk437nyHs7XAGSoF85iiQVZtoAPyETxKEzX6
u+qrfUwwn/qaT98UHO4nXc3IgjusXQIM1hR8cVFgDnYXxp9z8kMq+O0p7FdeFZue
ffp8PUarZG+rZ3o8BVTdAwjJ2OOqo1jxnP7gXbXnlMKTlrO0ChZEkj99aJWqHdXV
KLOeSY9tboWCIBWDeGR4dEoX7x3ZwZkEakZKV8eixPGTEvjQArDG5vvJUa7Cc8TA
Qi+3bEmfpijTLml/UavBzSENnpX53ys/No6smSNspHRFsIuKWrgZWmIMsB8+4ubj
UJcjtNYKG7lSTgntCNe62WuOxQVpC+iqoqRU5X0EFstlgtHOTnHofbSGY8L5OLwG
v93B4A1q/Z1bJtR+o/cfukBrJ2xX5ebovt2dpw5fKmxRZ6zcfFOfCIIA8SJS4/7c
R0+PicCk92Mm3stzZUhEce189bGK4ZcHPulOFhPnSNc6VNUFykp49XNyUDaDyCBU
Y22yy6t81Scxeu1i5IQ/mmo+YxZ+RWaL6TTiNFPG6mfTLtc5cG5mHqWnDXXCxhPR
qgW0kEmR3CEek05W5Gg0dqyzYxfKhA0liyjwKW5cNTVnQmhZGyS/IiLLt9eqM69c
yRi60A/mNE2t8qnZYA/Ghxd9C9QqJ2llRviiR+6+UpXI65kklUpQnSIGCf+8EZIP
Fl4DLMLkdKNfW48rUUIFCxC5ydox9B5QZtHbUcN/65Cu3PN7c7nEDp1J/6WDCDUc
b/g1EEOBe2MmYkVLd1pet3VUfFDx0yMdHGuv+YjC1+EDV+WL9QM1P2R7C4TAINK/
3YA5n/5HBDITMgLulsedQNV7sXb9C311/EnU8ezhTXh4VTWJDoG+3QD5KRZkJONR
I1IYITpnlxOP5foNlf/cmuDJxhYwCzOseyc9M8pyk9F47/Dw2Sqr2NmqpiCcKput
Mhp7lc20eQT4QomAc1D2b8M8nk9c+6qX+32qFJxXREQiDCsDtsEhZGkF9cInXsFB
VT36N/EQlEX5kHJBA+cWilBM6iGJuKPLrq4boZqju2L0hssy2sIfM2CM7rNQ4G26
U1isH7fE/hu9Ayhz8SJ9j2soysK5LTiLRczQnI+apAbzifF2ZqE80oxTdDdj1z2G
bSzFsazAU9NES0bTiklXy7/pxWQAgax7YtLI8NyETGusc/yWa7iWn983mxa/M7sY
dnyfjCpzKUvq5Hw1UPzynTmAA91NIyFwJQ55gzZIl8lSeLpnnmgfVMfKt+NkJgmZ
r5KcGzsddcJlo1EsKKUAH5AD983/wYyQ6hjAPH/onlYSKuARQaS747nJUGJDxI1M
VMEU2cwCnl3AHl4xZDDabBxu3/AYH3BSBedmMvLCwkOVK2TfvAeRamXXjZpaqW6x
OSKXaamUDxi1AoeiYxZ9kGi6tGcIXCuEMjOuasZaweQCiIwzvVsBQAKPUw2d5t9e
Xp9I1Na3+mZVjTU0UQFwsSJNX19KQj48mB5zSd3d59KV+3fWeCdpCEJOxJbMMbw9
fXvGEmUB+Zei5vQbTuknFB2WMSFLcsaZQMAtru9D8vYht5QRvK3nKa3Zlqy90jfw
gJlVUaAdHWDxp2nz+7kJTl/tebOv9P6ZriMiaZ8O3V51dxMK+A/n/8D/Nfi4t0fm
Fcq2Y/oMRGcDiydIhr0Rlkp6fqphLeodjXWrEjr21Y6UWrUYT0LM2gmKmdJsE3g+
40mBioKZXSsmcRnF+YfspqyvHvlHdXl0Zg86t0Gwu/aVGZyJh7fc2KaZ9fdUYKtQ
QKV9ZljUBZdrU6w/Bw8Om7aWqxXhpe0kTFTtgdD3Tic7dtU6FVKiiUaTZFH1xx3M
r6cqB3PfM8kxWoasOSCq39EW+WeZqjbEXawb+Ibid+YrCYdV/2rBYXmlebKFAlRc
7YUbZfHceRCjsjKeMvj2tD4QKn8CnAG1G6H63xTQ1NPDrhJVlBNeTmGpLsg5L6p8
TDTvj3LCvQnjA+DH+K2ZCqokeNoNc9MNz/+yl29KC6ubWF6ko3Sz19/IsK8fiH00
ygz4ysYDA1NxP8NSouJDzwBZmiTuChLfaag6xq9iWXICkKm2w2ucTMbfYtDjFSmR
D9jZz80a3WSldRyKiYjUaUULYdoGf5hHlZTonvHmEo30EW0pE8FbsrUx5tuTCabW
nc4MuACiW8MNlbANGDi/D0hZyCTqShfLbO+f8BHg7I2gd+mgExf+wjXFaNRwSGeu
S+pLqYlcXwqM9w6DWMxdYsrfpkuZdA2N0kVVjeptZLGqO5FKq8wJmvPONGJys+0r
a0VfynuPBXvMXyNrPZYbJoPXXJEAkwbq4kGQS+vUugUnTMd1DQgX+NzdLEuGMtaM
VvGywIo0TXDvSN5b/vOPgg4mFD5wMA81ueWykqPvhbHy9WmIqySEN/+RG9uWEZeH
/XdmD/adoEOgERHi3NHUoecnpjuIah+OYHTtIHaQ4Z/zmesp+0USLeRjOD6HrLXk
Kx9FTmiinJZWXww+DZdndWmPZzOTV49S7DZJ4lDDl54HpD8kBHDSOvzuEhkyr0n3
yGrAwICtmpH3BUQemxvCsohCmGUB/pupK/vTdfEptNYRnvWNqJj357imivojR8on
d1rLJWb6YN7fOnF+ORCEON/ZF06EmFi1w5ZnagXnEwuDrmo1t/j33ibXnbsDHTVP
PNrZTDcZ/E/h5wPqStKuz6fpnAdRcco3WqbriClkhdh4XLM1iDd5VMhqcHPGH4dI
bjde2AZz0Y04ZNluDxhkEjwECM2WTeB33s0q0RNGZekGjkEzJOe7noTVTml92Yl2
Vu3JL12nW4SvDIAroZgyzhLOVHemeS4KIlKeeS6kVm3ybNfOVsO68HZOehyie9r4
MMkofBVblC/pz4NHOcnZueHs4Vb9YGDglfORJHWzP+uLNycOiUCH+vWMfFluTI2p
5ss8L4bTo26sMPqei3va4WGS+DKSf5L25HOTucz6dE+IaZN+8ZUWTux0aNnBJG0j
CRaxb5yOCZEi9WmyD5nJShVIwGJK1zF4+oHfnnOTEpQadR2l0vuEtomzipXg20Yg
0brtE2x93gTP+pk7PgZjsSTIIfM+HSeymmU5UnIa5aec+XbnfY/1GvzkK81uItN7
1xHfX2b/3cV3avLhY4JgP4mYoVqX328/0mMAi1+woNwB2D7JqHUs95L22BR8/Yhr
K8PPro5iymLHpxsv9GLiMHpiH0IjvXFTIoKyIhMLJsML9z8vG6qRjoPwoHAIF08w
tLivAG5rhLHLrHw0vCJMYAYl6yc0E5I+1njlAy5wAb5sC6x55hW57jp2XaI0VsR3
7Fp6ct8VBcY0nWerTLIiTwkikLkuy+Z3q99Qb9+i+mMMrEa+864zT4gMcRdrtZ6D
fy0BtvgrXBo+/oAfzITgv0xPKC7y/WLxFmQigwGkXvHsLx5Jivg+jUBj+uzGwdr4
jxrywcIIhvoNg6PJC291H/ANyL97A5rwb/plkTdXuyyHNzlVpXqprUqSVrnCql0d
Pk5YGMP5Xx7AdFcUuYAad6XnlUmM4U5eQlpSco2BqQsPd369mJQuqhnwgBJGo8dE
XDYV/aRe5HJrqpAyTb/7jdGv7oV6tvTsKdRx9RSZ+6oqaNg+4FlOmXWfpqwlY9/t
O9RdUioOo3GT59bSjzVsXGdV+KjwA+l5EPgziFikzvNAOkmS6mBIX0TcXxN1f97t
+Q2K4ZdbcjbaM4vyk0QkBoXwM6+qB4wKZMsboLFQmWrT8ZS9X3qnuWJXeO3V0EYa
mFX5n6AsudSJ4SDC1Z2AooOOmlOwa66XgiPukKsRFtRK47Xaovzsfj9aiwr5LY2e
1if+OcLAwkfMWk0Ml5llbm3JO+OH0S+FQTLhZIwLG3tayv1y4sVUSpsc5p4eJzux
VPrJwHXE5mMCrqMv8Th692KUbMVVg9wQ8zfp2mxpW+PWyShTM+1Wr673f84Xtf/a
pUNoENY05sOk6ZnweFE7foZinfg4HgdB1mFBxdX5FNH5DuB8B/uRVvzGCquhJijx
kZjK+CYtHmi1huq3xVLqWM7s0z09K76KVfY0uMpDlNqCO9oKPoDvlt+yuYekSDHI
O8UOwqqyCqaJvUp0oIZGsNHfpOF6bx6FbU+UEHNTnniMcnOU8QauFZEf/QXfnE6L
50fAtF+w+C3XFWriHVAJYOwzkmbQm4Phk/PNNwH3hJUd14uxMh4Odx1iTnEc+jdY
KH3hfQH8NsX415myks+VJ9yybKYbqWcQzf9bldpW8W+gtKRHmEF4Api7LsSPWvUn
me85eRsmF7grMyJ9/v12apcPk9vH9PUnsq/lGrJCTjIq3eTpby7zs07SjjUfSXL0
YWHn6gVkqEbXSuPK8bEosvfEujrJY9iB4tP6FxRcbIx2gRhRCFKeF3mgQEbWovwJ
Q8z0hUMl1B9DfPkYeinct2b3SsaACZHPIQ7mrWQ+7Ruwgl2+8DvfrD+qOwRkOw3K
4RsfzhcxoU0jjyZBrqQ+hVjn2r6KfqVQclxZVpeO1bowZw9PQolpqjvnkHbx2J79
OQzxDH86P86kWUVfMzjCcjmKS73ZkJPVvB5g+HkR9Z6L6zMiIhDyytfKvv8Zem0F
4oMWICMnsUoCPfpiegtDYA4nz/X2QyMumTSo1WWosKE1kqBsGSqdD03BwrAATPAl
CrA9d2u/kbtC7f4RKuc2uvnJH79AR066csi1lL6/Dqoyl9dTx2/Bi7ffPnM+FBVH
Bx2PBMdaigGHhdeyccoTak2lINXc2xzmRtqg/+psheMqfjWCjxqBddYnnuJCiFds
SC2QAUQduGxqpQ3qmvtmAtAO+1vb0aZga0cIAIk2RFb6hUklCSvLQpaFRHSG/GXi
+W44ZRDJcMhWuFhy8x81g/FdYDXT9Lkf2BiWqHPqav25VYXtwf0+EkBsQ7AL3kg0
J13HzdnZL9w3UD1XhoJgPACWyeKCub6yVfMW+VP/nSUyg5fIFuavS5/zlTXKy/bR
DkkxrwilZ2lQqMed+iaFIEklLU7nckha0wbKc3D/lGg5TW7A6hhpkglAgYSE1DGD
IwJyABKLmmcipzIkkSJbCjwa/nY9g8FhBWs8p/pS+x4brKKdVQs5r9W1Dl1W3SZE
Ia86KUzfKbdrjKXi6cCBjONjmCZovwI5+VqDWKQA+HZUtygqTyQaNsuoDA0hg/UM
h4vyKKwejoNub9sjfM81uOgR0TDjhCpkxxmERqTTsZgWAOVXcI0CJMULICjqCdin
CsT+disaKLDt/WrofcEX5/xuqBOuVM+cLviF9+VCb49OpUitDWmoUo9ti53tPC3X
tr7W26mpkpffUVgtfGnrh7O+SRhAyBheos+Pq3Ig5YY9G0hvTc6pqEcGIfDVYPeH
5Odkrmrqz9hraQP9yHgRve2siq98GM/F7zp1EnuCOpUq0V/FHbE6wwMvz5QOqsgn
2J4RagoImkqpRH702uQRQnCWWE1lscZ8yQkpKj1/1iVxWM1z7PCGUM9e6wCqp2yr
NMkTHsBZ8A+vwXfzBDjH47zkaOvmAZHbvhLiamjiW5lT43KSeBPqvrKC/oWBL/rn
Qi8MPeQ8zlhHVv+AffUCEAhY6/f3maeIP61eysfjtjjnhBFTtMVlr2qHIh7dFtd0
141KRSGM691dsPlTqhG2a/V751Uam6ORqiyWHYfkcWIA1RV9oBR7pBHv7h8Bqh1E
Hc14fhxsVhlyiabCtbnwdaHOS2BvM6OzgtA5D5Mva1BlQbwFXsmX3oH/ph+qzQzY
ViYWA73Sx6+8RjjgWHdGTBtrz/x7B/UA2ZmmWnmm2XSgZoI72wLiFqopg1MLNFXW
Wonli76Wt7zXEYeFQ3OhVNas7Lpi+7rtzUDgPl+YEhWh7H64mkM7g7EWYl6FqL6A
5bDTSDSYGobPOH0hks1A2WJBxtcNTwywShw4dz0nt2oA27dqFEu2nibUByetE1Aj
fdlvrFYIVgOXlDNkzHqTeJIvg8aHWr9ZdTL8gGhvbW83YYy+D6Pk0Ur9A1pPr5Vq
hBtEGrM76Qm5iy+xeyubIOfERKJptQJ1iMnBYoEgbqdkZUUpQAlq6dg9PeqTYjcA
oFv4BjVagFFvz4sjnrkuwkOJ0R4c50cVZJ3KJIjgVD3zOobhxjYn+jKJMFRcS4g7
LEWwtPZ8n4LeAN0k2EvTbO/MVfoXRxmwyXiF8jUS5TS9+HV/ByYF2rXXJ4uj9JKn
/+2bviUcDKNo/iM7205ImWShvfvR72pxBF0JF/nd5/2iY88GYM0zDHD1fyhcJQnl
TLZP4LatMD/41Uu3+P6J7TMCTkm7xKAIZyL08ZIVYMSOqO/E3kOjCAYo6Fspb5qa
biHdbnkXThZJaY55WLGrnNk1iWaTfUnnV06fPc5Dhsm8HOLZzlXdRFg6sHmHRroD
HnpF7fkYkPPtjSwpCIzXSgktwIomhWB+V3IKYaBWKjPowoNECxrD1u50BaNaH/c8
AvKWCweFqAMFVYooyJrm+Yq6PWK+4FsNhkroxWjd72cxMXbMqRHOAB0DCqwhWaI2
VqvEIYUPhHDZBSl5Km/R7n8g+u0a05qmkbmPzpED+9U9mqeMhUBbTrv2oBq/eS25
VcSjhrdbKXnyfHUwn1eNHSzpwSplgU50sDoJzZXJGZ/QP71NZ2tE54QfLDJ8lDjx
G6Da3JITwjp6x6w9TQiITKxn2S1g06owIRYDjLnBwLUL/8q3QNpBG8Vo/kz+DhgI
9CJyRxctMw4waAE5GBZF1N9TIeH4TUJqlKeH89hXqFgLgoVGgaZ2M9Npk9dUl6i+
bM5CWCYZ8UMzkpoRW+Ji2NODIq68rEIOowsPKO7Emg6edX/RxKkObrBLE8VfMuqA
FjFDcydrJc9bd8/BX+KYCGya2eeix7lVAt1qTaVT02wFTSFMR//C2s8Oo+rAbM2O
8BGX0ieEROwhY6ytYNVtvShhx3AdurwrVmGnE8YBX53/b7IJ0Zieg8bZgvy5dAyb
O9kdr2NtM8D/KpBge3Z3hNDRwKwBdv9dFHxpAcUfq8+J21hmmzjZPPa6Ym9s4vKG
XBF1FZpbvpBkRYELc8z3cjCkUTsGkWKT4EOK7CvMW3L7E/fxZO1G/buXa9swB4Dn
A4EXXleIXF+VrG9n9NFSScQPweNVtNFUgbiTJmea9hHQzkwRqKHK09o0Z1NqqOV8
A0QpQOAvfMPuGEVfM31cOzFERUlMFEO182BYGIV6KxxIwZR9dWqXUhE77r79EdxP
ZLNBU/gM5vT/Duu36NtvUfHFTk77+y7Htnee6wE3wghmhaG8PMz2xu17zZKe4eGj
JZ1vpEie9mOA2nrPiZGiRNBxsPbkdhqZpnSk/dEucNFxUpzXnOwy5uO1FpSJZENy
PjdB6/9Y/HfvB7XVYShP7rUO/YrZ5rkuOsJpJRAt5GE46t28Patsoy3GvZ5EUW3w
Gis/xgKLKoHvfnsr0xbXVEwASUFJnFbMu1SXPNmilMxWIBcjDv3SkLLWzwIBqb8y
xS4008eOL3kD+29BoltOkSY7gghx5bQ6bsibCBBk0D1Bt6z99zHiIBUF41h9mRrm
bNT4DfIiBhs/32Zm2IHq5RyRrx72BRAQadKDIeH+uaCNRnh8Htj2s6eu3/R4sie4
RvKiFYge2qlJghsBznZzABvyMMrmKm9M3wXnlN8A0uCo7Q1dy85mfZKov9fAF7C7
Z5sQyfDzQbgLaZeeypiOCkNVrXcaXqybUE4VwzbFjZVb5S4+mLjBCHtScLtnTH11
HOFymuxA6W0cVB3VLxFm+MBiJqympGTP1JrSh/fzeL/yIKgkkJLfgP4UI7ET4BOa
yh0VOmnB2fwfYsHOBGl8UPWsHEhXduXeK2wDSEBxXO+i9UWQa/Q8mgIoeN8wjRP+
A58QEYWuCEeou2aCQI5LOIP/eaHPB+Q8WL14SOrrVYrvTGA2JyywIoatNJKeANFq
hi6UvhIzwd8m9UAOqDfhxW1r6hLaxQDWpjFrdBtOgDZuta+O1ERcBfC6DWPfNdzl
2Pjsldd9qwSPYU1bSikLa5xyf5Dsc+YOk1vhHtVLJBM7SVgikXf4KltgIsE1spFg
ncJG1dTYMe5PqPIsrYNf+9w3PBPELXCmjrTeGboRJZYw/loPtao8zF8f+Hb/+hjn
xhCLg/qhvZvB5PHIOKGBLddKirDIGYyxltQJJRdqFnRtqXgJRFiFumqbG5hUAXoY
DyDk2nj99b07OBdIQmXe475iqYXi+GoXIuK3xvOv5rP0JjgykMYI+Lou3Zqf1TcM
R379H8RBexiE0tuKtVVQY21F5XXiG6DJK5gWSVRCJog7L/rdtFN2zJZ5SrcYlvJ0
42/ao/xDkxc3XVjQ2DwWP8cuyKpAWAW35qxUD5L0lESjSLGuIzKcojd1bwyJSrOk
7tTVGu1vgPOU42Xe753plRmuz0+cOzO7xCYD+ZWGMwBmgC5+wg6Tu/a2EZpF41QJ
Z1WGIaEezt2H4crcgBqlhA3TI9UIR1m4149uf3ody4InhmXUUHqYvlRnkLllK4N0
4MyNawMDAIEEdUxyHiIWPUDxA8DMYZLsXW60J/1CE85SMh+ZZmh/JIklt8S5OT2b
dcaqFJEdrGdw1EG3Z3LvyjAsYXzDvmPu79Hm7Z0b+JnxT/1PRpSaxj3ao9Cmg83O
HYt1rQot+EsZcuKd/1sex4IYH4NA8avQPBDT+ZIpAOc06v837TI33YndvuXW6WNL
rBSDRo+RDwVNmWAly1XbYGy9QJsZy6397q+WKl0HNcs+hn/ZkD0SPYeVrONGstGf
911rXhYjHnbcENEJKgDGn6z/SWpuWTMLlbf/6VtICdU/WMmS30baDNxUYCOY33fR
vM63qjmcVDxzYtRnKuBlzIMnPx8HRlymajqOzcqjActnYHj6nApg1JTFvJFwRAPT
8HB/7Q9Lc4vZok+d6Z9qallcY9+Ab4uSW7KjRU0+YPTgXQv35MWlXxse3sp/X6Yb
AswrNCmbZtc2tNdtLkN2oWGlTEI2qSLkGyuAfWJRTiLlryP4j+wwQEGBPvWsEt0P
Mi91z9++YwifT94feRInF1JJAtslgTDSfh6pcWggNX/fT6RQgoEQDhLvcPEZ6SO/
1OXKoZJ0NDaauA/0cOg/rCyBDqM1OearfIRoluLtP1z6ajO3A0gxYkcQsKsLCInV
TENubZ4qlBvvFFCa6F4YOgL/GUftM3SUS1ZRkHdtI4266qnDcSNh3+S8a0qqS4hQ
r2L6RcRG9Y6lksfU2SNAdKUOQVocF6X2ljA7QG5QGNkVOlz2nOOVvf+dBOsM4XaZ
d6k3iwzfRTfuvNI/Y18t7KGquPae+agunyTb6eyl9LQZwe19EpNkZZxLYgmPx3hh
oKa9LITyccRrk0HeXOT5/t93jTbFWPoXS63Ywl8lfpKp3g1pLHkVMCmY4dli0mO4
5xGS7KJM2/P0q+lpXMnLS+vEkC52ZihNdsq7f5fExgfnOSblsTsAayhhlxPo0Ep9
JFLN33RSJTxtw6odvK9uT8SL4Y4D5Bs3gnwiz+nTN+bWg64kdCXrE2B1J5qC8dKR
+9/1khITdoVTDnt4uE72UYI1gsLLyz5QnRCVPxMmHUibOPpVsEKtutTkHF3BwglX
W0MSP+YX//oZ5Cs3ZkwmqclptCtHpkqTFk+PZ21GxNrE6btnEGsJ3CB7Ne8XYsJ0
7h49yMI8UDKAzJGzkkTUrxjyqBcNaUcCu45dzlOeBR/JjsW6YrXIQhzyDlnaP00E
GjhuH/bgI5KS7aWzPIyEvVm8kEG3aurzFy23N4WQj20QvRameGluzVrYqZHl0Rx0
SlLp+8xm4rfS1/CrE64Uit6FDCWu9t/EI/xPRM4hPUHXrTnVEel2e5UrgN557x8W
KYkSRAbZuLhr7e46rBCYjJoEv6UFCGCTHzR1SaJOlsELip4spKnHDTRguD8EOKfG
kn5vTbYi5UT/mca+lXWQmW9xY5ETskfHggcUPIn0kelfTWYK4N/JCEwERULcSJp9
Sx3APLk8p1l6pKiMwaZd1Xp8tkKq+WlNha9Q5lvcrXHCkBPp+MqglP0duU+QOn6C
B2hRujqeN5w46K5jvYaUvrYL32dMQhkj4fP9FUXA6ONkmVagBSnNE+CX+LfdjhTZ
5mJBKgBPlsxtaX+5W8F+JTTn6FZk/hFFyzF7P/9eFfGDG6QoaL2pCDtXIxXGb1/M
tfNplQz28m0BurCtxyMImj4aEqtCOcpNQz6VuefSypzv84qiw5fVNjJsQ+VnXPIW
IphPJKQbcvZN9mL12aZVkrvqWmHwGrhAgDsdE/b4j7eQ8kFlDAMXGY0f/Q6htFjp
RBa5xgutS8Ep+u1Vmq4e1HGUFWbDPa8zSVnTUSReVg9y6T2aImlW4fE7YuVEkJxd
n3WblnwRb186tYAiStY3ooV8a4RxIUv5BMV7ukn5Egm+4D1KAH906DWotQn+bdfW
J7a6ibZrSYkFGn4VE8FjMd+0/VHVFlTeaBaAmgIQun265vYA5WdtswCQN1E+12VM
/4fN3VRvkslEWYv/aik2XH9/assjQX/dpxZIXH/0qOMnTHjuEsX/C8ZPTM+h8jfS
P+SLMKLEkP+/xZWOP6b9LpM7OThPM9G9O7nztWC7EVIkCRfqOgqh7+J3tyfaabt5
L3NTLyBcJnGG+IWGApAeO0T5jT6wsipRa4XKKkzosvfwdTHE5D43uI4zH0lpfQm5
R0pc8MrBvEf2eyd49+EqwDvjudC+N3sJUMTzG3/yezZCV3jm8BMthFLOpYM6+x5Z
gphPnN1jCRQTxOt2vS99SIdZRz9zL2+5GkBbYBS4o+aDMZdHmvFcdETXANqwZ8Xs
Dbsbwk4SolwHVKBsXP/o4d9zzbKSrXTd9LYUgNgHOooAB8lTVjIIiniBcx0cqy/N
ZiVSYOwfgna/s4D/a1H5I2uEff+N8XMng4X4P5wxki490/eSWki49GhdKD5EFNGN
PZRekUcf2psBOJI65cpFpsFYBJntG72txPrL/UUWP2RPNTQxB+qQfhXbVXQ4+wL1
KFrcofDmLs/80+Fd7W+AdP3sCVvjqDGSu+5Eu4bOCEvM2u5biXiISUJC87EICYj6
aVhzuXXJERT4DLr7rGB0PYQvQit7qR8XPGXwEgEnoobiSP55JBN1npMPNEL3irxs
q+zq8utIG1Td3Fn2ICj0dff8Gf278HSfN09YwNvoBc6ng+XxDhoulfDwAk7UcVcY
/W22JzQByfPCH6oKMqBGnDfP00xYgEpskV1/9f5nnZEejwQKXTY1HCtgRM8ar1uL
SxPOG2BqUV7amD9nvEWidLIvgJvBXGPn5+ULOD7RxJeFWwXEbkgeoYB3mvaG2gGH
LBB9K+6XQr63lsbv5enSan9HOloxN6NOBeDKs+jVW7Tc8apxxFryCDI9EwbRsV/P
AoKL0+srbxZUrslDAXhTizmV1UrrNBpiOfQ+Z32nncslOnQMXNqKAQ/LnDro+ZQA
RVkpof9VYyhMd0viFZY2p/QNUfIzaG6iTBT0zUmiq0kJHfOwp++bsaIVnXBkZvqh
7kMziaX1py2mgaFVz03ag6xDnfJiJ2rgxN16osKtNZP0q2wrBBfQ8oS9SAnBLJpH
+kJPQTCTmhPMqu/c4xLAkSAq4hyfWiaYZssc2Uz9FXmS9KLrzbPHVF6u3Y45L3Jr
TuHKjUTS5i1jum2bW2bmeZ3hxc6v/pBUKZ7ypQMk+OFYMBXtQWZsv/+al4gwnoMQ
GREMsRekX6XZn3naZrTEpL4s00pPsLQjkiTQ6hP13+eZ0NTGqYhcFx3pDaG6N8Yz
q2qs3d89nQaDVXVhEqWB1spynPlhep8XzmRF9OPKC56YvUuP41QzkP02HrW5eMIo
8mfdZ7ksbx9FXIpalRpJjkpBcuvlkJ803xO0yqmBaAsEqp1xdGrxo/ICAfHHezZ6
tsvEo6X5E0xy57jrLfoknfuPjjPo/nnc/IZgcwjGc892vx66QxWdIbWuk9Xaf4Xh
WffJRUROYeG8DjLZpib2UYe3b/951LVOfzM8Az1ECXb7bE973977qQekvgD61p9L
Z1Ygea1tg9g9/9fsBWey/GhPl4FQ7jttcSekEYTg2XEk68vmxUZu+ZBBNzpmWGXO
X5d9IB03v+FtjJF6D3VLMuQwdLZic3HGcD01NTXLgSPPF0WYEyhS8pu75YG8O1pG
8TYPtXvD6NDJHfu67YmmhNt19B6sPPQ/IR5/rcklEEjM6UBeZ0qwT8DPkdQRDU1S
9x04+SHc1Bdm0SOoPCgHkCXi4jYS3+kh49pZvQMOVkkRZHrcBD85PoQd4eGPwmQk
5mbNWeXKsRAv3lbqKwTVi8/9rEXZZNv71mdnWzwLxgCnJwqcGsISmktFyFVv8opy
Cog4ckMbOWveOMi7a7vfhnusj5wYPTprkrq7nCbNSPgtHMY2wk7f0A0g3mGcNHgQ
l6rP7Q2GJiTTHdhqLNLsLVKwlBBLhnvCpIHN8y4mIdx6NYvzCsJpzRXAMKS3nwl4
HLJCTTYfnZgRNDr8nGszMLGiCYaCVVrkh2zFcq70xiJf7KxYNqIqRd6eVROIaBGW
geyKnAh9pACG3aRoFZ11qHOGt5ZfbmLAASjlc9Gm0oWa8abPbrDZhAjybPaaTCgH
BVsLOqATWfqgadxQV+Xmh1qDfNKUpOT1DaLk6ympKIOQsW6guP5gWJtNDrvE87ai
3TVZUIknh8clUIZ7yG8SU/xoSMNzjR2NThybFc6RgKe4l0cd/6RuFqmf584QT4qX
92/QflX0NDsuDPxQ7Yl8AwKfXLrNnLlr5lh4QgDG/P9XiY+md7+E3WWJwWvNAaQN
i58ol/0PyEzf1GkS96+bequ5jLNesKY4L0TtO5ZNtHjPIYZZC+4hzRQp8wnsE23G
bVEL20/jnx0h7b7mAKm46V/5+VKm9pwOf5JJ4Fe2f+DlPCINDnsyCzQsPkJRP3Cr
bB43eORW5YLEyGMogB5aDg01IIvpFCWPHONZvEahHzJ6i20cfk5TLOS3ghqYdLaW
skwBYPtOBNWsyn/V97ds7BDlGCEIwOSrXtLrzGeeJ5P0lmCfLQxTT6eJe6LUuc8Q
27UKVOZkxE+xaMqpuFMteSd/BbE4ePE4b3WBEZk2jmmTHDB9qtPWWNDmDMqm1qSc
K/eDgTXR7ZG88VQP+oWJvQcW0iMZQ4sJjmk4GUhMSTJZSjxwHK7PtSaGRlwn8atE
3hRFX0MZjZGZvi7PFdyrgVBT60gInlMaLziGn8aV5jbRvhxFATaOwaHPWKkWQRF3
W7V54HNlflCTzaBOltPlr0HluNK5GqT/V33FQLqXOGeYLnvlL/Ox4PAJP9G/shkg
sRnniUfqm75TcWlBEc3R3cu38Ea6Pa+b+qF6fYg4VIANa5q2MDeJN6jEh6s1T/Do
2g4YANEY021MqtD16TxmpbVIL2uGLxK6C7FDsaqX0PKOLTrlLi8Xhci3ohdsacmb
TxVkkCg6OLPp6eCLfa8nkWcF03UCJTbmUZeZ0lOVEb6c/lj1qtXe+AnMvNpwFe9o
ErMVo0JFnPlHoRr9K8slH4MwxLDOXe/PuF5ntefnxpYI7jjiyoNvkWJCS/bYoQeJ
kTwxZxDAbNcZIvaHqAZAOliI3XPuKjwi1uwHtLuzsj9gG9HUgVYBem9LOEhIqv45
njnZbnEsoZ7Xh+/xj/CsfTDGBZ78k//Dn7vUAIicsKfb1Etn5PTp0EARLLKoiL7G
NUYLueNOzSvd1wHe3mG7TZPwszxVqLE2eAFhTv+REBJljfcyhFzS7keHLJYYdLte
3Y9ORsrHcQxu+1RFhu+z7yLv2VGMQA+JBIczeS/LWir1efGn3uQBLLcZRzJC7D6d
T0MliJ97FEimXSRgRYhJmawfsA5yFrfbqQMiJwFN7J5phoN0+uSi1iLI8iGan/+F
O65ndWB+Yy5t+gLFZubvJ543aj7b6giuKGC4D3KlCiyHbFJjwr4IbtyrJpUtNiB+
6wkUJgXYUJYsnU7y3Z6lgunaavo02jrO+4Wuls/4QiMCB4qXD1XqRSaRQ9lAst/K
CtWG7mecV6W99xDPUngXpC9Zn5XOpPQjimyhbaYhfyKPduR6ygDoAJJMAyTxwe+F
q/PVrrS0AhwaM3EIlrBlx0PJTAgfLD16R/PQ1v6swlD2MGSvDPmYN4vt17SnZv4L
oj7OT2SMrkuFbu0mbr5OilZ8Sf1b5WVQXWEKq1pP/pegwUc21gd3x/51AcrzX/aq
H6OM9q5W29fp6tB21R7MZwmvMMNZ/3I9WCJ5nsxGTlaL+CM8QtHlCfFUoOD9l4ib
LyqxToyPsLVGS04G3+JISY2rhVSjLwBSdO8KYjfo00gFK7tGKuBd5CRGCS/Ozd9Y
QR8FIxvKKAZx6Iopj+dVtCqZaVKig5zRpGaPoQjWH1uAK0eaonZ6vyjhiKr9Ubsd
EYGLzvn1ntI4dEKVZySI+mT4NZggxO1hw7KvbHvCkIp1+Z7H2qPyuE2urg/OHw4H
YM6TQ9/ePlrCuEH6+vkH0qZVdRE05uV+yaUCUGURl/dkKObW3TVuI1NtkxaQuleh
mOzfUd+Q5vKcQgQm0Ua0et2HqYrKRfVNE7zTimijEjkJ1RdrhezRX9Fx9zT9imlh
XZt7vuRmlD2RV7Z92xkZcdSMNR1jDMjUvonXDgh4jmOcemMnep8B6Qg+G49rCNcE
mM3bfQ8s+s/6pZALCfT9dPnmt3OVX5IxbFTQ+L4uhvrkEPYvdnT/Wv6AdG11yn2W
c8AHRb/f2M8rM1QMhag/tnIHuhEomhba4ydDZDwnsVR27zbeOJn9H4rc6TfoxlkY
ma08eSlI5fVKDb49FVrf79VIJO1Mgtu0rz9gVIKlOkoL6dASItI1IgJSUvZOIvbg
sNGIXtWzoErgbDfP7rgulEHq4Z3THAiBDit+JFCraUyAt2kW0gybtpoyjpLxcBra
LMf0JcNoXiZVidMinJoRL5UBdVGvvsaKRGNePnVou+izpiv8wr/pYalWySLk3yOT
P6duXY4ktPJ7Ft+KYCtcy1dy1ETpPhly48mAepCn5JqCVMnEhWcQ8mtO7UuCjGKX
7h+0BiVskJ7q3gVCIAUg9Iy85sF/ri/+gaKuGJ1kh+spyqqY28C7JL2EqSMH4P0a
WU6pqkDJOQMB4veot/pq+F/higkuH9RJRs+6P/gBJps9cQtMEW2NPoAlib0kT63H
JYes0Exh/Meex19OfhvjiusClDkKo8vhqQq/bNN5rn1EU2QGgrH0ZwJzwE20ns80
xNkKBVd1YwO0mJ9IyaBEQGlhkIyilECtVBmz4U5cOLYbtflPnVOzx+Kw1TOcnYwr
IsqRRIbpWmZi3NTqeYiPKwSPqBR3G7Wkw5urwF+0Qo76uEj8tZZa29N8RQ0Pzepd
NmL7cD9WOX06td9NVioWn0R9IFLpSv6/IKnIVuc+xos65NOfAoX5xZmSL4QvZskI
Xypi1bpVRLUm1BloaAWaMg2syOBNvddQ85W87MrxFfC2k0waeY9OIzRJTOQXGAJ/
g6nWWVSRVALaPaO6Sh/qkZT6axqLoBuzTCmdBfRoNn73gBpUqe6YQjLTA/H652nC
XqYaEN5Hm8q14yUFatndpWmFwI3gOZyTcXCcg17OMqoC4nxneK5XtoAOa3uExWfy
o1xqQeQfcvVTMCTVErowSjK9xgtUwiQM/SCOQ9+2L2dEGCxrAlqei1XEGejdyd6s
e8B3Neuk4SHjG0/1aV+4/gvnPh6Odrl6Kfm4utnrXKjBmvsfsgWTymyvB2WmCdbT
sXk10CYDv/gAngaiuD1cQ5puo8QEovKqV8henPHgWu/H0OHpbW3Ej05+bIZL/Dmw
wE4BrxaV7uH3vajzlVNpUxR62ig/0kZN4TMW3ktShBZMU/FeX3drLId4IAR/nT1N
f81aCY4dH52KbslL0Spsc6FNnII46mfh+w66QhkOcCUdR5VzX1va9hp7nFwVDmYH
6ueZ7uJhgNIMIuNetHkehfsui+UQCW/gd1MHQDlNh/EI0Iuk1MFkc7Wr8AxBSl3M
HsRcHxMrkmwqn0i03BvcYZLyFO9U6iSvI5dElCxiPWyvK7VeulB702RB2RBoaZ6z
RkUOVPEca3/6z/gKOuEesyRvm/khN+QtP0au9/SN6DhgVv6oXGnAMHlURBvWRFhT
rJyufTsiQW8sKiExpzgm0NtGZcY04JqM1c1zpLI+UjXPzfMK0NYtFCax0q+lpzP6
DMdez4Xvigqf18Qh0ibDCxMu9Iuf5AJa2Kk8vlPUCzhBVKwq/aalMbL4QldvmqZ0
fjJ/wb+RFb0aqPqCQ4FcMpTxcXX84UpUQiuJRWObusP4RTc2u2UWoWYqh9PVOjGZ
OHXjrwwDFKo0vjdiJTUVmUWySwsdA9ENI2s0QSFyoXcLpX+NM9+fZZXhNDsscJce
4Ve2oeMI9Ab86bVOqRd5YndRKxFE/BuCEriREccMJtbDu36vMy48JHV6Ztqkyklj
Bgp+4IhfWRvBg3/UAfu8tG+DwCAKa0z9DL/qATnAVOBNE1kR7DFFMxCclLNbxCqt
kMwetoEkCknMMzV0ZYJL1ihWF+TF5ghBV07Fu1B1aZZGy3kf8WmGUNwQjzjKEAzH
v4QMIJuV+mO1qeAwaTCdxPNlB+pWfSnAwsqoEmITkvKoqfbHkyP5yPCb5xiwgspq
EQShUVNnOJ9UfGx5aBfZFWBf1T3AFeiQ1ysgH+nUtNfUDXOULvMAarFzz9XtiCho
N2YBM/ET2ug/ltdVAXnj6lAw5vAMYCG1prbfqqWSQKPs0h2JaxxBXUS63uzGUCpo
ei8s8uYA24DfQQWsGxv6PsLHa2C/4v2hdKAGm4Y2asbYTd9Me3ZxW5yzwHMGfvVo
75U3/U/GVDR7lzk2+rOHmI+ziCsslSLp3siA9OaeYqgGI74ccb6NnwmueXs1Ej5U
yu9VWg4C8qM6+cqmVsRXY3VuE9r246E1I9Oxpwi8rnd6Ow9wMA0mjE0wqCJ2sGDl
ECws7PaUhbOyw7V6pIRbQ6yqkbf5TOnaqpF/m/V07PptXkIq6Jq8J5t/IuP6bOI/
mSpiFRvKGypBZYUBqVyD27Q6NJuGkPPmmkhp8/2/5/JqDA77ZOMzLOGnXxaZtIk+
iVaAtWD9INJ5UlnmKn4vLTKloERD4nv2mzfZrsfvz2LSSiqvVrLJRWwnppHpMMs1
/T1k33Jzf/3RSdWBk/emtnbreSYBqVoRLi2ior5V18rUmpmVzbkVwAGaVzhqnYkz
7Q9maJa0V5iTFic/HhYLQ6T5i1gY77cYWoO7IAceSoW7DNaN2h1d1wh4tjWqljzx
aWPZptw37y9qB75ucd3fPnI0UCM9K55YJ717F7tYtY2MBiD/C3qdYvS7xbOjCo8A
wrESru301p/8gyj4CzmKnWjzAsBdcpc/3AKI0wVAsrkb/Rba9WVsbeYuiJbvyrBN
kTBV/AgH2+u6QY7ac0XV2D2NnnfTHb58/AXQnTQoI6Es01LbfAbBPVlmGBfRKEG9
3TBWlZreLOoPJ/N442A3M4kjl7VW0tKY1Ax3z8gKIAPChzyBGUoLI/qDQnOAwz1o
syn74uN5756jsQur88s6Jk/Jv+3m3nZnYHmQTxuIAShXN1vYySf9z8qYV7brDWtl
mdloyTNIHQSpZtVkPaKGQ4k/IMMZONBE/mbv9NySaGTEmj6pVc55/QmFqvwMzEWE
ZSBzTX/WI8zga4jtrGbDyFmUmYEvZY9fJKC1Z42BrWhwMFPRSmGk5ROn9IB3uJDY
6V+/mxzXryHWGmq5ST7T76jkq0QrQqdzOln4KJ3JWWFnoc8JiCIIKZE8D9PgK8Zv
TuVMNWHftfW9VMNBc1tniE3ZjfwS5u3Y19bgXm6dmBsIZx0oV/VE9lXFrO39Dg1l
M1HhFTL3D+ifDxHiE2MrPBJQjjOiTkDrEg0E14xl3ZgBavv519hVWYUJr5Rb5dEm
NkFjHnum05nnkjWv/jpb2tlQU/jFDwR/6xR/OP9aiRhumrQAdBtLr03o32WzKX34
t4xSDDNfvm8Rv29qlPXA62ZoeRd4NRhEJgMoO17ouI4Kr92OnTMJ7WVMO354PGDb
gR3HDw1GhtUwTMRqaxBNfYOmV0YthfCSWf0uSeGP/qfWZCOmHGsIELvAS7wZiRbK
rI+munJf505STmwQs1XMhXc5Mr8zteL7K2scgKF5GKf9luvwNOc+x1uMsgjZiCIY
I9yMXu0fgphpX/r0mZqlFAYN4AgAqbZphA17d5KdrGxndewYS9GJNh27Lz3LrV73
HMNAYbiVsgVMkh1EY76Qr7fqY4tAz6D4vjg2jpwrWmUXpfNklwqjMFfutFfP0qKj
glD23zsPxdWTCX0t5Lsc+RARYeqTE+MOsjZG9kROtAK23od2OWHW93wDyFHAnTGL
1QUmJBbDBgu5y0K1KZw3+oC8uTAI87dGyrkyS61DzA2YJ+Iiazgi8FakO902Os4b
nPo7WGFcc9Au/F9A4gGzrzMShFSSis6tKZXDgIWFv1/+7v3xTf8xuCVmxlscHmJe
Gu96O5wp99CtyF+teJFe32yM2wsozAQgMiB6U0P6rIy5lgsTeNrNWULVpFikXLbv
lpu2V5trhfDBOKO81H2PjAugceE0UsQ7S9bfgSFE4LGnByYb+/LWJwabEply2STP
OxmYZMxa7k5gHnTHeMI8PT+izlWrARN+yf6qHVo3Y89yaOKDFktnFlnx4tlr4r+e
xUG4pzzrf7H2+ysTk6I1spv31P1cgDZgmfLF15924C4gwegeOcy9ATdGGQe0+R/x
8TMCozO4McEb5D9zSBm5aS3LF+HVpqjbZpLk+8tpi0YdIezwA0Lor+cNAo8ItlfM
+Y01WrR/b8yjqFHdzTE73bEfNowB/lnnp2JXTWWfI5fnk1OM5WxaP4MQymLjbq4F
X04XRpSZx4ogoJZ9l59xL+FK5/RGp/8A6gSQEt2SgrfPdQ4o6hFhvyyMzRW0h5Ru
SrKjQdcbjsfbbdxNfllr5W0t4EpxShIZ7K7dexnT5FR+1vJ1JM71imP9QjsGCnAn
SIjHaHqMl6h+MqM2Iteb6Ahe5WXWMi1EMuNVmF2zxyH5592a8riyPKVoJSYZRxzE
BVUrzxbvtMNTNZVE0lMLh6ROSR74H6i6X9eK5ZMHeDo1KTt34CRzApag8m71FWy5
5P0AFydytE+PLJops/9jU4CIsuxcTNUJrzpZ/prm/hBmmBZbra0LqRImI2gfxtgE
5loohmXvcgSexlXphGB8xZBrkgj37IPTlRKlbILgqNW99kk6cPsa7ougudNjUkrk
YpmZih2wvosbCwA3BGM9OK49t59lbmsA/FAS8NLMAsFEEmxnJ17KgF2UOYYO6TvC
ZLTMU9REA9ds0D/dWnMwO/A8RhtDhjPFve0x6jLbfda+4HyuttRYlUxpoKOIS6FB
LAJa+CdBsbmr6vxABA7oFv4AD3IpDPbZP+8yi+pC+e++3IEI2auoOiC2CBngBK37
NerqhaZG+jA7io3qCkt9ggFc92yygdCh3uX83WKWyIZbNnDIjBrYLuJWpuvURlZ4
ldA4esR7slWJRbT5NFBMpyyPxwxtuOiKpxCRAwT0oALJjtHvunV9yvltrGV+fwDU
ivqnnuWeQT95ixyopwmSd9l9xhhKchJN5RZzQ8aRdS1n89bE5lxQSpHIhgyghR39
ePQca+gj/RtC7HoM9Zm6HvljnXGvwrdHoCGU2sIKT2dGtiaU5zt22HNNUEmYmxTC
X3nWDmNlBFBCxQXM46YgXN7EDhm+ZTd4wCA8uGfiQ7Lej0j3UzTVPpeYetttszbV
otcWbTHsund0U435PdHTRDPBUfnAKQh7GfFX+YUwasPW9eQB0uuVDEegJxleRTB2
PCh9aE5iX3/h1HH92c0BsRYJSTc9r98VxmHVBboaZRkor6LsaVhbpVOaMWrxPO2u
BFVfXyC0n4JPpnCIg3Uk69+7BCMRCvaaRVLr990hAmd3s5GrMnRHCItcGYRNnsTM
3zmiAY+RLUOXyYzWCjhistu+Z0+nGet1oZgr8O9M7m6o96M5QVWflDdw2n8neTSU
TvSkjJhC1XL3m/dsM3YBfo0dbwirVcd4pV0UFczr11SMBAYM+/xNZQTVnupYw5Qz
eGjTWHrEjWUb+fRacWI6nBVMcQL8f/QQmT+q6s5Xr4fB/eE0dlc3NoBCFFtjfHR6
wpONVksOL353qqT7EOEduEAPM1aicj9J92vcL8eG7aj/zGXDI4atfBs+Brs9AFx9
fz+zQj4KyWfu+Ryx0uHTUbFzJa+k1a5Rzxz9wZRd5jjE9149CQ0n6bOx+xKOskoA
Zd5ETQqKULL7+mDxjQwgWoHBILUy4Im7u+1tBi2TkB3N7Sl1BR6zmbEtIPzBSKTn
+Z1d1FA9ANkToWpNzJ4QYyywqgbn/DRnrJK4Ic2WPcvitBWSqFK3ZUsc5ZDITvAT
jPklcfiKPxbj1eD1OAr8Xfj7VwXXj/vOIdJ9pqyDg/MOEFm2RGAy4g+Qb2JvHgcD
UZqTgPmbCYe0C+3ESEBefHh0P/ScuG38/mEeFG8VkQt1rWiA1e0sCPanOrEzgbzB
cYt8aX9Ly3Qm0/OfP32fODFFGxcBALoyPu3qU8Q2Tgdy2VTu74MEq2jajGbIGLFS
fyh1Os7kPsWavr59oIAyDzk4Vcq/Nb39Q3kX3EP2CtI0ku6tcD03GBsA8CHioLTP
XAxoviFSMWgEBxy+DNhYlykcWx93iAQ/cYr3SlleqPkfu5SgMFLDjLnQzN5CbPCw
kDxZ8IjXjy22IpERPbUD+NMegOmt0AnebfSkqLOgIZoRRbUaKlVl34kjY4JjGio4
dSizOyJwSPLxTDeHqNryKBOykzje1FNC43RjbBPCmxWX896Q11FT7XpjhkzolSkq
Cbtn6bycxKwmwL2EdJi4pjMd8I9zBSDbVgP24WhKJCD0R9q2Sb6A/PbWiK8whlCk
ct0ERV1y564QcM4ezeW1rXPbQN4BnnenxOq+YQfZApCifBNFBPMXcCvnA86Y9Bxw
vfuvliGb0LT4igyeD7DZZMTMxCiG4BXZLVJpJYI/l6Ywqlk9xR524flkfCbIncEy
76Gyi3FdzFwoYDuX3elN9Oz3J1YLQGoLPi+HXBpjPPHUtQhFT5QRxHRyaIdkEwBv
AptyTqqYPOkQAiiL1QSjdK2a9qnHyd9u6sE53SzPxakvCS9eI1+DL5fNiBRL29q7
Q7EZ83jI7Wjknr54PhkjfZZeeI2xC/+9D5kOC1wM28IcAp3Yyli71mw6AX9evWKq
/0SKL5EN22shZ5aNwTTUKk/2Yn4MIxaLjSLfZp7kYYhlLGJYhcBLC9kzjpni2ZiX
6QlDeCNZDBG3Pwi4j9dMY6Maq5U4CKnVkB5gBUwYUAAUGhbGDW6uI8jXEZRfvpYl
9xLo4emmjhZSC5vBjK2iLXcBJ43Po/ed89DsoJQxYayNlbFvq0OWB4QmYd0twfnM
eu6zn4GQ27tHb8NhWe+gKTWOblVjmEdwzBE9UwpRk6M75vHfW3zf6Yiv0xv9HI7j
AEeb3Neh2J0RKberKoY13fjxueHb97hZS6k1fVAr6EUsHp7TEGFkDs5loW7GhYNC
wCVRUThnVf+u5CnSyEz9Z7LeSGohpd4nrxVNov2OSXRC3CG+QRaMeYodqkJQeX6D
fJ62o83QSSR5+hJVyrRKto+j/8fNhcB1vuNcldPJlgbaKiYe2z9Pe1B2BQnU//sK
75iaS8sUi6qDrMo2s/44gHsX5XfZjtcJvQ9QH7wm7eWaZacwSon8iGFQkwgsCz5s
Bqf4ba4Llku46+Sjf5Ebx1BgKTYca/TLDeLE3AVHQF0WHoqBAE1qsLxVy07vgEqx
t0AQ8qTXY5fLRAyMr6NcIzHyobMjxz49urZqYFX69RpTRRONHDEYQmyFTpUUYIl7
Unr9c6V4aylwOspXon6IvvRx6e0XMKVrjPRc6QlKEO8SXyn/INQ9MS6dOjb1ynrX
Bn3iQg6xYFLycxpptVLqtJCncV2zY8GccMiZnQD8Gj2m1OWBxvEjIWByiE9504F0
1TZREJcbRxbglRHfw2K3Ir1X5RW6Pj1jEBZbWKfUBpys7H1ostXQn6jo5xlr3YOe
4gqxJ4CKhOtTQU5Vn0CPjavcGOI2RwLlhytrxshDKAAkTESh63fSzv4M4wLFvnlu
KlUps7INXiaNHcBFreDcWUymRooA6dDO8ZdKPFp+SD+FRt7TyAsqzY+LEab36mya
0bFi1if7tVElc5BRXqaT0UlbQVUOCE3XqD8WLznAMgA5Iq3Qks8RHGJnsSbeB0iR
c0hvfFSwTMEMycjcIz0Zkc8dAroACIeuiiuDPM+PV24RsYPLlflXCSM1Ed5kaJ1L
S/OsMdwU9OoYPABSlmr6fh6ZSzf3haT077PBVKQ1Hv6FfjvCcJxfgFC6Mv3Mn2H1
Ou6pCre43uDY6Bn4Ww2HitSKJk7fM5pSGPDkN5vsvDNPD6Zz8u86Pc7YU54eeowJ
4w1TcjTtkGSvUkpau5wZWrUhQ2FsEksQrhcj4IupykQJjNRp+LIgxUWq8OyC4VX4
wZVuEZppeMO4xHyENZaIrfi1zp+zq9XZDBacx3cgq8PiGTxzKI/hQSoTooElrOvN
n4xOoyr9Sfm+tKEe+jfstw9Ct+eDWIi9Smyv/83ilN/iS3Zjn9ySBwAX6A8qMPHd
DOK1h2AU/fzk7vzbKw5uu8YKuY3kchN5S02Ole2Rc4+AMzCqnG6whXMdtoYd01g8
jnGSli9oqhxROdV4R8pJGLTc0w+FTe53gcZWgZvEiwib2ex3G8J+I1zT3LBUBR9X
eTKjO68VH8TQnH/5IOD4LnguC0rlNVqz1iRsKLpKrXw6Sf6uAsXid1GgLzT/mOpu
ICExRr3QagEbPf0reJPQcdLQrwBuurozuX3Xf7k2ADzoqg5d2b1SMREemINAxTvc
5I1LDnELXetJnDQ9aUYir6jKZX6cx+4FxcSBPvTltLL2ftZ/HdxKW+k/I+h5ANr5
HgIgQv125af0UcEQcntIpBHHXEhmzUrGZQtymuq9/ccmn/x4rjKYgXA22a4iIlUl
Pl7ejznvZuVPWEVz+PexXGBlsaljKkUy2hOKcJTq0/JHoARYZkVXxEKz/obWTxpu
SRj/UeX91SoRghRw+a7YAn6VI4UlVK8XvvP/zSaZA02gEHtOlLNUFASKyjD8W0fI
scfJAU7WeaFPSHzthBOs5L5EjkTURpR0PFIC3H1HfOqIntZh+2c3Or4mEQ7XURAQ
6i3OKx7lpXdcX9l5i8kpmNeqN/gfI9grhlinicIC74KcvlXPLauuxswVJkBKwXFT
BA2b+Ns0bO/H4LILz+z7E33ca1//xSRMV77mhQBFL6bm65ZhO0TZlS9UEVwspsR8
6xLU+bKO5eS7PzM2hK2Ne4c6yGdPUiDAz3KfZNq7z4Ji64GMQT2+vionaoeiq0cT
+Rmp/XelJ1Qu0+HPg4wHoBN6/ubjEX0f1bXUPiZP3Gh0ndrV/086q52ybAOQ5X03
dCXHT5xj4cm5I3GYVpJpKxLW8iPmIwNbcPtTNph1nynlEOpNBbBscIb+vGAymSSu
FcnppqgMp1TUFtgjLlLw5nbE1KzV7GsFhcZH5bCrhfq0rTcVOqtCPs/qE6kd9WoJ
uoHDopDNfxl8f/AXJCClNg6EkL+H77B+Yf9J6um4ozw82O0Rjz5JAB6mkvJjLv7i
SaNAcXJWZjg9m0klisoWhdCpB31dza1RwsTGYzTXxIsodhqDTJggBjSY98rW4T0J
MVv761lqu8sczmQIH2WEQNyjPBMXbo++4v/iBduz1fObbyF/ZOk1+mdQGw1xLj5E
9PGFdZ4rkrk/ZlXYvC+eP2V6djANpyR1DbeOokVSfPqmAIAOVfe7jS6tOyIT3O4c
JfOcF/5tBCsoYCTBC74oplDcvuAWEWRG3fHhdGcsrZyaH62lIMV7sd8ewmjf2Djs
NP0j24o8+5NPZr8nF4nMBBtmgXjrcPeKN79biIwlN8SjUAaUwLoO6QYDNM/k+Pfm
qAr2rEmhcufYxNaNW1iONG0PbK0x5AT8iVYE1Xu7kByumosfdnhB+imuIJWdMAUM
ketF6ImwauO5pSykg3o7Pb/3/CYyXWJng/9j7BnndHEnUnsuDdcAJslA3CQskfyv
f6D/ugZyuOboWfXqWoF9ElCcFA/+CnHjYDalKmrlORQo/R9EyEXzY3jlTf2pZgwg
XZIr6MKoTt3LH1ZehEe2z9sPw6Sf6fN8F0kkwV/3TyJc4YF9NgOFUBdeXNld5G/S
NyF2Ic4cGpDPSEaWPjbq4dV47dVim9W1isSOiTq+gtrpbCO3E3zijzaBrQBWY4bP
wR4mcDcXbDwTpV8nbbce95YqEHYjWd+BZl+m74lPssR9x2zlThWSK6WdCqSeXDGJ
vwwLVLE6D3IAufhFXuEQQuRLCMaXbe9g8meV1Lr14CFwIJ3jDebojCQcGuY3Tfgl
/Ml4wHEvGGOVIO4E/RaSywX1GALVhXdyGVJw967PFUdiSxD1JRfrWC9FQJOMSIWl
d4Hu1q4YHMdMeWX7E+5zRGm3atEKfONleM7nSQt9ojD+dV7I6kf6AkP2/tk+yJDP
WtP3dr0DByrPWSOSD9yAw/jWVtHuRrgbFg6arhp56LwywatNyna+x+p+ZqdUm/4W
iVRZr1r+UZ1rxdemGwVFs6sEi0mJ9kuoVTjLShlZ4XsAEt+pTO6IRcjUQlsEBiJN
3r0Op70wOT+dCc7pVrYsanN0trDcbTZFESLZ62ArGN32CMWWyUjNAtiYPC+vwl0q
DQ4MLEGfiNlUVwz//zoHOJ/NXYYQDrCIusu/dl1elui2OCkif8QP883HPjCYqNnm
QRRRQZbin05mXgMVoup2UW5O8qa4f+YFOe3hEjlw1ltM1psSqWl8htednu4rmwSI
PlnJhNdlz8DIeLJxF8ed33BfYHTtr9ic1Vh6KiUNypZo0DOxZGR/o7WVrgNLEPxW
zshBcZxezc8dDm1+rXz5SNTBZDh9dCfhF3rxPlR3/t1Fj+0eJf3CLEoZh1kgJMQs
XsBdhz0dP6XSQH1KM1u1ZmtM+j7F1jbsj7inbob3rrBwvt8IFgIoHCHxje+IVd8a
bZCAg+enKge9OIFuxtIrtG/JAlWuGph8xjDFFSdnmMQS1sVIhAGhD85Z97orV5AY
bWReLg8IHX6iOxjUBjBDjgQ25/cmz7dWxQHivuXdsGungnEGqHfR0MllTkvXvT1C
8MEfePUDbCh6k4/bjdSxRWHfbNClktgG6ql3ydt5Bq48CftDh0SMpq094vOtG4WS
PtFSNcZrQ6Ifg69P7BXbcHB+psY/L5jROnAkCnV0qwQreMzL9gXuZeOf4Hw2Svgq
oZq5Roif52Z3RoQf3BU26YgNXmBcpkxjgwgjIuRubEuZJM0q6er6gaTHNRzSCwur
gOtgDWXfI4ypF8SO5GQ9inyGSWgtWxh0nFUC6F3pWDWmsxRWRZEGopCeIHJBCUbL
Nz8Sme55JcM2eiAt0IQCplR4UjVZEWO+e/qhln4MSQgiZKOTqtESj3Ld8A5ln5ER
jEitnIhHxjqyh0YfE2EmCG1TolulF5+L5ZCuGaWJFh2rDO9YsdYM3zxhgWmNR1Ks
JJ5bmYsebD/U4xEisgHDpLnB+0gNYHoRD25SZYDOOz30yH2Tt938/RvQKHHH4nMP
T6s6G4QOqEq4nWcTvy3Nixqk8XidBK71pGj7SAFyjl7L8MwkKpMV8+OWtdTjQeZY
29Fo2J613QEBbE789AZLG3om925HUogm8UBvBIa6YRjkRHVRc6OhQmwjaPYL62LP
HrH5MXxzcDD3qWhTWOQvwPoW83mytBp7f8gDVuC7SW1YzJFDjZgh1Kwg0m3Nr9Lx
qU7JEypSfyWCmOCEwPy1pnEqqoG0oIelfSHBThz7vpBi3G7lR+1q0xYRaUPinQt3
7j1uO9GDzTcE9I2i/hgSjviJrT7FpTziyf5h1ttsWWME3MFXbPuUQyeZKzpRIUzx
ftyk6/UNbyDcGAuegaGXVAuJ2GPr+zpSDQc561GHL1yoNXuLPEHyuSyG9v7lHG9v
pBV2utTE0npyOrx3L4YycYNM/7+GCGJ0xPH7J6eNc8xpJZPOmzcM7QwGhA5xQgxH
Nb5s8bBZyGP68ayUXZV/SuTICpfb9YJuZPAHX2XTmaAOAXWNzVHW/Usf6IhXTDta
JGIbui1F8xnxspcTqcTvJ+UiGkS4XkA6pcK4OxJu06NOk1l57NKu8/vpGqRSaTOC
+llg64E3ltVPZFYxBGCBMJ7hsV2EFklKAP0pNAyEQVn6sBTnZWwo2cXI15n6Oa9N
AIHe7QXXjpneis+pKsEnFMg8orh6uqton5AOdf9ZkH6f+H6d2fuuxtv2rVBhPON2
jOp5PeLRXdt02VfRw9pCdR6QjcTgnZP4+r+z88Y5EWTt5maJdKNUexjBWC1OTZ7y
aEdnMzACxby4F9/R2zXqHZbZcGe1Kir6GwCoZTyiPJsKswFAM4HiMvbsCYrKAH9V
B/UpfvskW1lza11sVg6KSca7JpsF7GBB8XzR5CAoHe3LcsVoilm6j/dGFAIjd09m
uNZMysYyOax07yKwIjnQq2+4EitOh426l3Y7uqmrHRg0W0ghjuwkszWeSPrUoCah
LPOi9/vNsZJOA7JNtKQLLJnOQF0HOmAsq+zWpI9oaBdndg3aqnZaWDc+wFsw8lSy
nsA3m63igJjzWSGuuMWwUP5mLKlDDAfMAfD5N6ki95a2MDtPkiR6iK/opV2nKEjY
siE8h3K/I71150zVzGZHvEP0Sq30SM9dzWZNYYzSW8hSSZLI1RvMug6l0BvP42Wc
7WaTzNPUXj+CoBwzhtZcGfASYIDhrVeaCdHJFa8irbC8tPzB40PRCnCSgF6CIzkw
J+4EoOBRfdJ27sTf1zIs9wvuGvsYhHzkLzmOUoKnveHUq9fud9YrP+3UD7cf6uk4
geQgF5BAFz87lqeKgjb8H4+QvhTC6cFouFCEbyFV7BXbIIWCylZW1+xywKG37twe
cQt4lltWF9gcxJ0bVVSxmBCIO0/d68p8G7Hwq3lEGNPj9Dm8CBesqajJW2j3V8xp
IppNyUpHSU/C24ANScMVejtOMRhhgoBv/vJDJTjxHqHgvMcVghJwd1jcpx2+EnV1
Lu/rQtPnYkhZutPOKdLUPElrtgJ8QBIsDgUC3i1rLthRAa5u1GEJsrKJEESfXRq/
O3ox7hRSgZDtJk73BIFInuKsJ9TVjPc2H0tN6vPPenMbYq5oa/VFVT9Sxs4mVevE
perIvqoCW/UuuVmgWJy4RJovAhi3dldiU+fkCUE2AXH5h4rLqS1R6tUvKH4mQQ8d
UWVm8AifM42PO2wNKdFmWy0886MBZf6Mgc1B63b6XKgeUzZm4wXwCvOZB+GAXebZ
qolUR7VT3tcGG6lU3J3P/AO9rGuGaAfAjysTibgMdH5KDi/hNBhk5zn4ons2G/I0
OY97P3MHY2tEvYZBhctqrws/yjIddvjQHTVKGXh5qVDAzGnVJLdjNWnasRHuJVCG
ZEGDRFN1zluzPQ1SsDr9puhBEEKhOIGRjPBsAod+wPZeN7zRHXuTzyQ9/MnWjF4q
WxHhceGgT6BOwS9e4KUEMCdgZtOD2aP7nx/ZMXrldXd+4UXlHfljRH7VxfjjQMbM
+GqxfdHMNDLclmo+1se3R41S4Ns++tIKkPST2GP6VZS7SkObchGTN5EYXT/eMQI+
gmhAxrQ9N3TMfY2MZ3Nc/BwrZatIWj7w1qrO4FkuZOv8GSl1P0tkPs82ZUOa2h4v
m2xGhep+B26W7uMY1LgN8k8J86n3PKvu/lza1fCuYqK3DIfofq8pNS2Hi2AhON61
+2Ao4HzjNJjSdAvkqpqPsYU5og7QZlY3+buvJm2d2Q1gJaj9AUoDv85fhc9OZlny
TdM5Rt5JKF3cvm/4JdvLnXdMtExbDt+v3GP/U0LMhcEniVM6fLQZPhH3B2H7dLz6
bFpieSzJIqvYVj3EYy3ED9NB+07SulHwE1W+eWZoe0BZ/ywirB5xKAd8b2k/6YLd
zpW6q7b/jy6khFaht8PJWvV9KIYYDS+wCYnnInSexnsrsv59QgIIbnXbLPxD8BE8
0p5H587FkYsomyRh3GRS2ERlxBLtzkj9slhhYWGgxVabTMKXMWqSrk+BG80vG5ur
Q/sYnnYVEjgtCn8TZfBgLs1lF30fxRLLVx3gFEkWVCSSvUxH3hHJvJ8K5SyybAxI
ORjl9JbtXfNywOjkVIqwDQfy490EHxuYGWVWi+aabogpfpK30fiH+40+5EXXx3+n
xVKMbt4RSJdSFtWucixZCW93TIIhJyKZgISjWVX+b2uXnAJN20jXXm74HhvIPUsO
mc8MT7u2Ok1IX5znqWBrHQa66LIleWJzwM3E4IGb5Zub1hPjCb47mKeCyGIpboc2
TFOtT0THkB261D6Twi3aUDX7hZNmVlY46YWFf0dQXIXdiAF0Tufedj7TYsTwb9aM
aWMeADpJIvmnHOukyX7YnA6W1bDi4SZVywYqPzOgBJ4Nj2AR0eGi/zeCq+SD0+nz
rYsc91kk2/b63uW+fm0QoL5IB5ec2y98hhhsfYfx8OIP30RRFfroL3QoOC+0B7tc
uuNMemxpc72ROD1oDTJGc76EnT9Y5x6SzamiVbYkRW3IV1Mh6owKQ0p0K+SGfpgO
XyI5PKfPVKAUu6xxbSARwNpUv0imFIOEpAYIdDOxPbcYoOLBdNRvR12eModysmgN
5L1xSwDhW879BD6Am/4POMMRAo5DR5Mi+RdV/WvrE8uX4e13o8s9T1rKMPY2Tczw
76sR9HcEoDeU/RUMxl0kxB/dLwS/NCqoevwdg7rxHa8I1iO38RoNkl199ooC8G55
Yl9m6YR9s8jM6vu03RA7ESnz3liIhmosyaDm3Bk3BL4puJ/m2QGSdPxDvN0DgSJn
wCuonlDgPS3xv0DF11+rHTLZGiE7Y/8fFJHA8ONnHeXQ8frYq3g0mlpDcr9F8lTS
JPLBjCSoLtEGWNcgx3k+5oSt2xLdC29CCsIfoNkE9WpqZg4KZaJKXCMBc130pHLm
YQGXWyw3lc8FtOIv+N4m2PDKO2nRzU+GnHF/kTxyD5bCjVe+dfU+zjZtSpmsIgeo
KLeifCBOtV0k37HKoE83lY+xC6SjadLD3J5ZU4z6wSaMAzm9bIchbuoBsGkoYI96
ME5SaztkUfwkpoQ1kszu/lpHZ5pEHgCVOwQHezD7v51vJNbOoeqsmeKPfL222q7G
lt6HbqZdvu3FIi56Z/hbTeVxAURYRcD322jUshvOdGAHdigXj79EGy1pCvdN1Bgm
MWAKyohKY/P3SAPvRq0TChmfMEl7tk3By7/5q6D8iePnoWd9I11/UShAmkFDhTl2
3eiBmtU2Skoj4eyj+RPu9SkS/69Dh8NpKuS+7j6NMucZqPk8yfnB1hmsXUtgnSHs
xxz8lr3Y63DITmdpjOjm4jKYUi3mbAwUf7EjsP/7T8JQFlVP7w2G8DWMR7JnmwUb
/uxFUBdpQ+x5t0YuvR7mbTNps39HVGsEAfM9/WdVxrySgAt8wRLs7kMXt46tfuMJ
RWbtaWFovwOEjE1A8G3P5yqDDHU7p9+bfnYPlutavM11ls99kn5EBxUor1fByXbG
YNpWTYkul/Y1znwuTcsNKpodHPaodU8MA7X42HmHd9VguFo/qp2h38HNCGDCzjv2
TE7Obt82QRFkNVZdeE6lpaxCt9CxbcnhY9D8QO7CLqCyRfS6ZTzjcveT7tSUJK0L
VICtydQAI/3okN4VcbjRFXp1o5G03n2XveNCNpVVdIPkbEWl+jXIjHeRRfYpg8Xc
RPJokwTBHgbFm1wFdve6ZxIYTJ0v4iur7IWeKBHGuwxj/B+VIh0lQvr+vclnJuhe
m4iCFvQJmJ7wJgEkm5GMrFDsGykgSGqB/4tcBi9784WUTEIz0qmOIQEfYkhOE3AW
i1nvFZ0edZeoYp4JAt/FhS51zzMuSFKw1Kv/gwUoFZqgRLBJk7vlH55o2H3+IynN
P8v81j/16yORXondsCPURYOSwdnB8aKDGUPuuTPj5lYNSFgmeOKfJ3G8p6aYrrBp
v3nCj4hbBecVYJFF8Dwj2iXj6KbjKQ6qMkkqGLAXbHMF2pJwfVgta4wB1dp7qKe8
l8WbOW9fyHU71saWSLYQVLUJF48sjOf2xX2dhoxZBKKBiPFa0YWyh/65tXEnpK9X
O+XQmuzEmuIg6hTnoFfSqNzB+RklIHfIJbMjlKCLMbTxIl+ZtNy13qEMRQGeghAU
rFn9Nt+GQcOwG+HMC8yXa8tY+uQvYN3IGeufcbmrsY7bDvu7FA7b/dz7J9fW3bq/
zEp/S1QUYEDvMqzcaE3RVMjPzP1CD8McHKcx6VkaRV26wOUlsWJ4fc0rgl2dYH5x
dVQLq41DseWJpG8Z58QTi+GZCNFdgD7AsgKhOdYT+lgYafrZJNl3uumvkQCWE4In
O58EE44o7LHCTuBjELekjo/yH5TAAK43nkiZz2aMWjlzsAGpl0S/FARx5YD4PzXk
GqinYA05aLw5teKOPwj/lGEkGSCywA2qkAbBA0OKKmvfgnwTxVMRkMZlHC0q0ERY
fCaZNEnjYrclohuUJi8XXX9/D4nJnExaeiNc3cVTax4ZlShwKwOqd/1QhOFFdkLw
9eFyZ9KxeySw9Bn5+bpaLcJmp+P7xB+IwEdFbXcBDLudi6s7So1KwSFcYvmA4qnv
E2TGdOqWdItdQk7RZ3hCRK1WFFfwMRahJ8KOWHSGGmn736ue+wCl0alPpcwGgnkU
y+rAh05AouVo/kYgo9B0l2NIV1a46ADOH7Yc3pNVy8M2Auavq77tkS1vF/Kw23qt
cseiAURc5oNwmqk5JJFGvkC0tp3QC4/Od+Qens+ljYmhXLwyWRP7XDj0XCjBEn2y
wyPq7jTkaBrujhXYgEYlK6qMIfMOHhNqKBWhpxIqLYpJHaBe22zqtceMpgeWIVmt
kOIRSDoidM9BTkOAcBKvpsu2h3Woc/evpyL4OLLEGbMBHdAXblPFGqhvJB8Nl6p7
UG42RjGC1EqHb+VH7WdrqzTirA07Cdc8ctVlqpH4m6nVg0HRZcdsMwZ5a+EP7MhI
pYChJ3i6VHQv0/u4XMhxGUb6z7+IHoWYBo3oIzVh6MR5iLaiYVhLfkRQeviBGbIJ
O1Dds/otgsQbrHr+Ez2vzxV3O9lMdm3qP/XjZ87bGd+Okm/uE+cVOL7Sz6Zjn21U
bxkN0W/b8yY82T4Zrs/1RyhRrW1m3WeO3P4Kbcv/unCpuTE/jhSl2XtwcYdPDjS6
D+yLPF0lmnCc5QiqawCWUf/6d2jiXemDwAQTMBVeWOZlFbNIkax//lP20X3TGfDy
8agqf24LcDlCya2UyD0tPcrCyawPWCaIXfIoXH+24q9T1exi7L4I/gfZ+neWglKX
PmMKgkj+ddjFMe7b9SXpzcPVMEVTuO9amI1PCDyj9ahS9bBf+vYzHMtpm9uOSgP6
M4As3/M/O884/GjfEPIYtyIw9LCX8TdEs1oH8wxnMewUMW09J0B0ZMYcIT1GMuym
IvFcIqX7M5ILXhdcHmoZay4ZcwbmfmuHN7KMPHB92sU+CJwEF9R4xI2+55k6XO6d
IG0oFwnTWgmR01AY5HNjeaXCUZUHPdnzjOCMYA0xuIxheYQGoH9RfoA1tQBjxpcX
hNVwJxsJFsrdIlvxlz88nO6y3WWn8+5oMZTuLwQgUrrCZKk301dKiryVT4UbKnXO
Mu/TkEKoaudoquGIxgFPXXClfL8mJqw83OXQyXaEGVEEbOCEqw6r4x0fGtOtGMD6
Oh4eTvpvAD/gmZHiq7O9z8JA4NDUF0R6M682P7+bYDcFLV7e0QtveLp1M6fctNfj
kaY44KfHtCb7Wechv5xXdN5KBfTC87O/2klw4jnzB5O76f7p9uT+TRQ1ZYIX1Mec
KJlAvSGQGfDTxYdePDRyPN+6zm2/2hWthU1J/XjfeBJfcVad5EfgtGKA5p7cH0V1
cBW29L/cmCi3ktyHmFpJzXsC8gZAmfS8KSSYby2/ihRCUVfiR77OETvJLuJAn+GN
RZHzvmChPxwRt2WC53W7lx4CLCDTxmFZ7apmU5gPrJMUyPqBpGbIf9X4QiQaD5jb
wcQYO4XbZqfLo3TDrfD+LKvCXnSSHlogCNuWyLBNIAOkLdEULVQo7SL4YWvETBcu
iqfUMYjH3ij+ypWHaL/pAhBksCjREtloJCbk/IVKOaPHOjzrdze12POAzVEYKUkM
7qjZ5Z7qXv+G2NPOEuqM2dLHBBtgHSKvFMdD8wirmnnPepNeYLfzwiIi+x3lLRjg
vfjXQWuXKw9bou7zRV6rBnRQkXcaZZSX0cDsKNvk1RT51gHVYPvNpW+XGM9+IH8f
5gBXA7T6o/rxsX7lythsA770ELVrKthKPpljiAmxJOk8sBwu9XGvCjyTWKSBX41n
VKBvhnV1tJQA5PgK3QTIqOKoASypecTVemd7PH3syel10lT4TAJeQ/7lNmQo7pLS
IAYIEFRXbEEQnAo+THD3xKgvghqjXIOrCp2mwQaxq44WeajlIkkdoJC0miENoZyt
pTBFCEi0OLQFjSxHDUXnzM0gSA8z9KL39t0tnq8abgZqDsPoS7n6+jrILIFUmi6R
C0WytZepdPKWiqugKhbnEJJoUni+Q8LLqZVyYX/vlmX4rTja3WzYFva7SGDnpDMJ
Z+A6Gql3Z/F64BQBNzXIaf2e0N1q/BF2tTVox12+8ZtYPl+bzcvX0pkoLJOGgQIW
cmUIQ9cicqSJdYGoEZ5XnpwSO6JFgOdPXedLhZjPh/twNmEL9U77K6w6q/VVcbt0
yACaEOdeQK/OF1FrEpozM5fswU2oFmpZKbu6AV/LI5AZO51mZiNcIrl3lGS3cYAt
l+cUxDWLpMrnD59rMhSbPQp/WUFN5z6r/2mJ58UFBE3BTMqGjMe9u8mrsbvRf2KJ
KLS9+zHhzImqS8FngAOmgjm8YdZxUwZ5ab+TJmQVHHnTkkNhYbVROuvDAIOGYQnG
LiTNPtoY6xyD+qTKZZs9jDoDyuIgchjOecLlxxKRHtw+wwV/7Z5ZRXYMOlx6rhFF
sfQHysPVMDqQV5v8qnbO8I5mifqG79GFzWqeJFCnrhbnkQJ4GOlsAjXkNGTJoxPJ
zK5Xga4+vO5tbL/vm+x4nQhZUKU2vftU2PLrDHx/Z42EGNg2wye8vwz7GZdm7Ddy
nITT98Qm8j1Sw3q18g4K8XTOOBiNh+eJEbrW+fRBmCcKPP03kYXEJ3EAWVmWbUi1
eX9QePFhKOc+VmjvoHA4Qy0SUzJvCBEoeNFoKjaXDs9+PTFTS8nJhHlveFxKzlV8
y9q10NS40+HrckC6R5EAdVvrEaRcIVbdgtPZjG5zC2fGlNIy2xtOplRDfn+w7GXW
6Hm8rmcA6mSGn0NwHzV4k6tF6jcadSU2USNkBI78AACVRMfw6zO1l4C2Ilz06Loy
qNTVj9Q+uY8WezUzJYkL386lbMO5Vjftrk5W/ognU6PXJ9gbRmy91Y2feSB8GHNJ
40D9jSzguBYv4I2tx2ROLW3MmzxHGa62b0J9Z2fY5sJoKhJX+wXmsVuYVuoBVU9/
iuupwAHlgVkTAHJ5PkxfiZSdMDgG/rsmujES1PxggNXil0CdWT4KFE8wfsVrSvrX
zwzJx0d84kdxY2PjNKSCOeJ3Cy0tr2XIReJ3A9yu4KIC52U1/q+cMXWBB3ZKZseP
B6g9q6CQO9hU24U6fR/MyXFXntNtZhg9ZACoXsHsV4HnWjxcTc/dauXfYI+SPMjV
C3T1Qx+Y6WtRuw4ZEXbECu9pzl0jkfiJA8OX+rEPmImKseJSNip48ureHQGHjmhl
+kR59W/qtKwlAsCR3LUDo4QfS04uzTEa7pvsk98A5dVyx/gIEUpFsxDp3uBobBkJ
S8SAuAjNE7IyaEHgzoKxdlSPuAFGDH/asLFiECBefTeY//AgvIhMVWVt2rbfaXWL
xXjU/WbfGHVC+VM+vFpJXKroi6MtaAjD3onQN6T2xLGpKpXnnugGqyozA4V01pVt
JCqAI5IhaxX/NXLAsATzVJnXXGUf9txWs2ciDOhcjchz9bVizd73bQJI/p9qJxDV
rr27h64xs+7n86M0refjV4I+2sD4LhBfaQdMBdzPHN5rivnKJGDWZSsYBKD8wYNa
wa6HSnWDsLStUh50TF8HIZuzCWch0dJMf4PT26qD92wRa7SlWSUXpw7yXREt0hWu
7f66YEVGDwDAMXdrY9Ldyn3cj5TwCgAJyyYZJgCrbFnxioFahh26CG4EwATzmOt2
Z6xe2iHV+vHF2nvqRVfmnWw8vlmRKJmaeZLmBm7GbRtbdDG5oF8icmgv1d5T2WDr
ZjHhH+xZC4tcRBFesEx0JVr2xzZ25lCc2JDwZU+cB7CNERQoy88O8Fhaup5VGg1C
4lVS74oXQT/QgJ7KYmigvA3B2DvJMWWU88dCEErp9PdeiJMNRWxpJFtreCvUAFJs
lKnmHdnwz3nbS9Ho7+GaEXF7wgAijH4JKINEKJIdpwTk+r0pm2wqCi3NQWsm67iA
pYKJwzTTS+1fZDupVUXw5lYPwO8J6brIZ4+tRG8M0T/3wnYuDF4KAXJ67TL79iQi
70QHB24TdBt3QGovQDNZfVOxeFCqEwwvKLi1N4u+hKk8C12GYuuDwaKmcwk9E3eK
YANZC1OBcttv6ZVMGAK2o8LTtcesSQZY+k2kIKcc/NFD8a1SaU3wPknxGz1m1+S+
hDRO/DcyUUpPLkLl8hIqvMdGyKyjGxE+OL1ADK1gyX1QZ3nCcZ2oEFFRs1FdS5sv
FxDtJwni15MJgkvo1a08bz99rSf9JltG7wjbpQXutrKB50T2dwmoX4KU5ouRniox
dJa0N3OihH/rGj9WViMlbxDet0Ii75yy5Dssxtkh+XQ8qz9fkC7qnB7BS7AYCdvp
YVEO/vGuC+nT2O+VDor46Q3fsc3BLY/uVSyo1lTqUyCNPYOYKvjuS0usnjUTzXwH
G5N7MgeFkL0QZd3WRXL9nQe9nZvZS2YnM4wACPEcrNjgogKql0KfjASd0BP5v/+U
w/snqY2XXDLm2AqCwjQFyyUTQKp0JC81PcZJcLynJaq9/TRk6UWMWZ8SsE8X485J
hjqfTzVIm3ohNf5eYUZ6hAZL5mi6otgdrBUA+BIln7dA0DlEPo/esI1RaqyJyJgj
x0kwl2RemvWKIApqtAg0w6Yb+AhVo6MsRQflKcYOMEcwlEJQAfnFW2UiXX6MXTe/
OKXxxSPQ5bHaRvfS09cbGY3U1gBG0S+hiNrzl5YF98xRV6p+jg/13HaBsmi1jdUx
su0jypqldtChDDUqo0Q5Wl6Oc6WEOGgg7rIZTw0t8WeeTNaezWHZQ/6O3zdphrur
PlzOlEUvaTzHPMTALRr0mJvTpCc0xfr6viH2INcJECnbwm5U86EyxdgPm+5dkSiQ
Y5Y47Ajc6jhH6wHXwO29d91NQXcLOulCGVRGwizgDVLQkwVdRA6Dzzeoy7AxTHgc
FOfF9V/OtlbEJ2dbLCdOHYd5jchwZe/UUk6q1oMQFyumODOvAuYd+kSyrMUyeoDl
TOmAmEngsgwk4yINbsv0DN3F/VCWfDgOuqlG6ltrM7g9BYLXFUZpRyk1CDtAl1ZT
ZNeiWA1m5BkQ0qhTxYAaqDWhf/AD2PJS5bMg7XW1O/nH8TlaEiDi3R5B57q3q8B2
rSl6/5+ex+UI5MK4q8bOfAmoIt9XOV2vlVcC7BJ/+ZQT+MCFMG60fpIrGzZBKf2a
VPC4n7X/ph3UIpWnKoDyjjyhtiK6kFbmnmH7qVU0qOHmbf1KNC+PqCSb+dbZtIgX
vdxfHIpApXe0zI28ss+yNiU+d9AiS+2A7imdYcbYKuwWP8gGcvmLdv3zK/eAwcQP
C/0ndsdUZA1sdrp+NnF10IU9bT0HCk9Kbg7PZgLMvKz79EJ4yESS6sfcsv5BzoAR
wMS4YeXQDVLnsb3peD1B0GhPdU9OQHsSKloj7HvEcir6kckOd6lkAG3WPctwWhoQ
Bs0BWdg7VUkCuC8HIcou8YNypGw1DTntdGYkoZ2PrHgRJ8RllRSywGLxu9MyxnV5
vr6FSysae2b3E0OjyVjuTELX+uHIog0BVp/jPdhw7/v+kHrRHeY0SpwcoK8SfOtT
Z9MtUhUzNpcBtu4OkQQQP+fUY2nOc//0RMRAAoKQdT23rOtmuedj3W6So1D3FV2a
X6wh/qr/sZGoxTJ6iLyowYQU2xD89ZRJCXzUed9DxdyiwfUoxbqbbkgJ6qycZxOE
Os/JMGSr5Gr2RpaUOYc5mBFxTK4UKO87SaDCAEYTujuynvvU/U5nZ9+EklHQA03W
PjLDneg+ujb1/Yn7RJeWGHBcurs9xlR47lxhtbfujwNyR/vlh10g1XOvUEzW7nex
p905CDJzVoyWaTIKPs1Dtkm9Jjxl+s+e9N7CvYUlz3BGpUO6yO4Tm/t4hQZkLSy3
wZUuSwkQJRjqVz06FgRKc+5fT/quFMJo2dIPCzwiZkstakilN/CGQ5/r+XcPUgsC
INtKp+AZfJ3teheaukjEtZFIuKxcaPHY9IUcMwldzGJ088Uhx4xus0TIs8I6R0Y+
CRcIJX5qaFJP2/xklfMzf4LT9aVknCbQKIOekzpDdmdR4rLzLmoo+liSSMKEEO65
bW8YquQh0Te+R7EB6vXsfoF6rCdDgCBN3S5hN/UJmjMsaG0BMLetVyLJu8Pe/AfD
Gh5Gsyt0SF4E+cJeKpq1TJv18Nkyq4QC25Mqpc9YLA62RzZ75jRQvYEAVZGwP9ZU
WkLvDo+aDTBOiFJuHkg6GZXXFdtHaRTGZ+vmz5LEvZvKLt9fzqSHmvAEhzkThxSH
jyCu5qSkGihqqjeKRkIDzea7tMMjoPu4f9xZ8Xxlbs96iPgBwirzVkROItlmNDUs
cmALAIH5qA+9FEYHnukUWPNicPUP/bSb56fy47iIP+mYvDUPgGFqbYAU14+qir5j
b2Cfidh7EqC+fXN5jw/PU/ewfBOlTEBSX8Adnjoka5cIPewa3xuBtdrBpok3RMHW
/GpiTcDsfNNwkTVDWNXv5EHjDEP75npPMotEfvrTJgRM572lZiU5UQAPGCcBj4EF
MHCYiFDJsA4X9oNQUC2cG4s7iEiUfBaZ88JLR/sqY/65tNSP869P9r9koKJR8hCy
KWuT6rP0qi+yssy8J1IGdIezvqUSiDo5oaFMNH5DiG36t6vCSVpKskIhuc566tGo
pXLo7Y4iCLXFxu0u64DmqoH8biBH+h2UghMgVdcIAq8HD6x0bjY9J+WGGWTGoTHX
xxlhds3divOuYY034dy1Bco4IDgthIAOrAsfDlEg6ERP1H+qjzvS5mB9thDHgboY
wA+iHtBjjngjLo/IIvIu0C6f7Gdu4vi51Eakla5Q6WbM6ysxuyj9vAtmUXhlqHN1
oNQ6f2VI2DX9kPmANsilq+PaAjbL6ABPdKgATgo6IlfW8THwV7FF+roWfhPt8pz5
S0tgKDOPpe31LpzzuVbTOXrxxh0OewnUToebqDuKi18Ltm/wpW5Kss4Mn01URFev
Ps8d936o6K9ZX5+h/w+AEfsplJ5inMd3ddtF8o5Fy585s/LyW7+nyFlr3fCqUUDA
9XQD3GX3ayeI7bGQQws9TrocbkHYuWKUOyviZ63AHJsyVNQf7LjrKxFvekL0AOaz
ilP+Fo7SQBE7kEhJo1dvD+rPFlCruWvKabqlH+VwjRii5qTpzOoCuyZKly/Yr4mr
VXEcd7AHJyz9py0KOkDQBqclub7mjrs00xbIdDNx296lKrx6kOe+cbZ53VaqgFSM
A54P8O72Q6+lomW0ywULgZ/fSOHqPtmNnvIrngE0O90MVw1wFoUXzGpegymUybJG
NYa9nbVeMcnyeiGhOFwQNwJur6YqBwdqxNH7IjqvkCzNVyTPBKoWEoVHzG+AUTCo
pTXiazlaI5rXBL/FNWxG/vM7P38jDUs2y3td7h0awpuxbk/+332yC6uz1p+2An/8
uhrW9R/M7nBnTmsNqKCySLd9qDmOZG57KhScolY57KgeEE25ofR3JqATGRthjKyu
w2j2X/50CV7AsfA2ijz0EEzmEvMYKAO8oP/ACkeyYOHq3PD58ZeFL4wsEko6M8N6
whE7WDZbyn7kWC9VSQYQffco7+tZRrt/efPa4npO8CLL0iH1KfCzXxrHEr8ZbULv
HC41Xv5c3W5Q7Wj9Yg6YMjT2kttCyKqOfYousXPGEO6Ri+rEHFqNCKrq2tXVkF4K
x5xOKL3iO6G3Cgc31/z2YHZGqABQukNbYbASqEEYDaSQTyN9CDUQwfcVMzfPeMTJ
WdW0T2GWLjFx0jfoFMz02QyS7AyNkjV+2wmklOR1+qVTYwd+lGASIag4XYFggl2Q
5YhaYxFIxw74odv6jlHF26148nyUcOyG3zG+qxm0upBUslTPrTpEtDBy7UWFG5Q8
wKbs2ZuGaoBE+FHuND2d/yc3pFA6P20XENkeCHPJej8NgEWPJkUJnrs9lppBoUFM
O7Rb+LKnKNVQVjEiwQiWzgIsYpqzuc0Xy+SM6Lv+4gxOuGZdsd2I3VfH0t/myeRo
QeGub5kXSc72ZTKUlQQd1qi8C8H52SkPLIAj1eGawsichwLMc3PS7zm3CB9OpyTN
BgM/gf3krwQ8wlf19Kjq3WgZF1gdEM36QjQ4b9xIQq8sJ6sDoynbSSMdvFL0Loij
MUE02IaTW++wKKw78hN/sEA+b4Vrz7mEAjEzl3YM6AOWHe95D34f6nKuSRBaxVIT
RhVNsvPOQRx1503PZdzwprlnQh2j1l7AvolquY/ONoDwS6NXpdxmGjCTHCKFJmRQ
7wgeRZrqTZEl4c2bDD/YizosD+OPcvfzlp1wlTPLlb0tWGN9H26R3bpqKZMLfc3d
ykIbT2/RRNUDdCeOlg5FKbYTaiVoxEuHfRfFsdtmZTKSxyE9cBUffREpNQMcxBKX
4eo6503T7wCyOYgIo+ATsocvNdGsaDoEzKG/gvml1JZxzeXyrCPKpOKsKUt6HVP7
785iP2PqIJaA/8cmpT2hRVEgUq1HPnnWyD5y8bNDIibOiqyQ2YEVFV1A3GY0TYR3
UF3LH9xw6oxeAbx8zSenRoh+eD61BNBpsjVblGdR5UcPXg0NJJQqy9Ux5kRM5oyZ
zfmApdBCETsja3EO6QuU2RAI7/vTkA0syBoeS4ux+HlppsUNERXJaKOvH3/pXs1h
ewf9aKUP86lY3ul0zawdgt+S2JhvYUashoNzmjnnWORn+9KWv4WjQDFv5sTTU+eQ
MZlnJq8c53Y2pvVbfH1WudJVbKopHzZprB0xJnx2+lWj7Md7a99I/BJTrr74adu7
bpUdzPnd8kwJn16M0hBcFYXjxRDpsLO6RMKpD9SGqcfwhFHqhz2p7HpjN+kvcd/z
mDih1MJFZSi4mIkp9797KMK0OW9kAiORpzBthIUYnTvdlrImkRl7IHHjLWCTrj4E
I0aiInJNoBZlBZZtW9Ka1nJk0ZSLyEZK+i/uCAp1YKbbrcL3jDve8ISJTeD4yW59
OYRUEcp/TWtmpq46kYl2bgv33Cqf0MwB7IIT/KicZUF3th45t22tIjLCY37DzBAp
/uYoqWJs/kj6iGobt5ZPOtM4cMAlsTUBgnsk2LfUZqAF7mVdz2iaaXFG1vkertuQ
uIElKY8ifuVhfW2mQ4MyIbQW2nJu4bIqc0xHSZRM7/Zqlca8c95CMdGL0sNcCMBd
5fiy2pYUnRvwUPvLxVy5FnF7wAE2XjTy+9Bv8SPNSXy7uJ71yTWvXgnsFugQGell
WkPDSM14dLlCEXveWFoYAnk7LG9LuSwQ/kTPg5/VqRHo80Dx14Rqh/89nUecOjyE
fhLnyfsQxuIz9qsGRjpz+I5/iayZhoArHzpUMkiir9wW2uN0W6hsI06od30jRdCJ
VBN4ulufc02FXyz7NBdRr/JvdngSeHBlyrifJXejeVFCEKHlQ/ZNoSGMDfIEi1dH
ONp4lRhbDeZoTtr4gJKqbQ7lzoG6p5ZWZe22m7ElFm0hBYYjqvwkip7eansG60aq
eMjiD+W68vgXKhSO1LaZzIEuRZX31duQdPWN7krc32C0vHfjOAzrZVShZ5cuw2qn
k3T5LTrGQ3yeqpri5b7WAPcl/nQGwMnXbuoXniqlXBpeGTKgc/Z6wBh6bJtv6+lq
dug6NuCMCOvK5ddyZnucQi85mmARSOCqrjfh6uRToMbj4N0rU5XYHCV6VOJR2Qom
7vGUPbl6aEfuftr+fKPkdxhUaAXcd5CtGY/AlMBobIZ31jHG5XzUGeM7Q85iGbxy
O0HY3dXhxvB4/P8pyRY/E9yX/+pZj0EF2Lg3Td1U4+5SIM6DGcMbkxhNxFCbMv4Q
oI0iMuDZQGVUDYER+B8ve12LvUyzfg23ht70ERQupKQEIM9vedBLcENb9jPZBJxB
KzxpwSMEF0AkModYCfzEMZM2tph+P3l43T9NVnboArXnXyzIsf1TPtg247LgLDjX
xxo155tWfIw5Vdp+oUPv1KdS8yZqNHctFrWAW+Jb3IQ4RULTUNVOmx75ih+SWTpv
zNX0TmpxPmZM4Yn5zx6DPgGr6gAQrbO5M62ZONK8uElKDKEthb3PMdf7nUEDcrvp
sYoWzrQaSxkzDjOr1pmTVT/klj4VokhCxIDxCARAekbrMmjbvD8gVJ06OrHrUFSn
zBCzneoyqA9GbcPSTX1eZwUtkUBunMkqPuy8kDABqIRiv+y68jgnpJMjJzT/qwDM
7gu2XEn7EVw5CV2QQ0QNO3gDk3sV5Uk+uLMRUMjSKIkYNy7NlKBihKAYKzmvsqqu
HgWa0XcXGMUbrAB5kDr0rFCJu+oZHNm0GpWhxh9nwIxRqfI8NYVeFJJ8FIKAayyy
PvXoG3CMQ1tGIfo5Ed2j3e4Yh+PCZUxAM5KlOeXbT0P0HEfuPW/3LTcPkFSzN465
Nx0k62JludvEBi9ah6yGc+AxYgltNmW8DVkUGKDrHKsmxQGL20cVxigb2/A41GnJ
BBL9VknVIrW6l9vxsP/+/HxWFT2hAn4oROxb/HpqmzCQHQrV27ObSihOVRpR6lzb
wejSK2j7cS1ozi4EyM+C0uzJxcOrmIOLfP356zUVpnzvFF8lD+0uak+/b/0qVZxg
sUNwxwCvBK7ecA85mmo5uonGAoMqV4JMMlHF3kUbsKszB5qM/0+0HypzhQ7GDTt2
JHWRTHmAUMhXuv7W1ZaWgmQ3hmVTk3fG9Qy6G/Q0GydkksM389zs3hCX30U7R2k/
8CWJF5o3EtV3pOJl4CJhi5Ty7HbyPVPIV0j/BsAonY+Mc1BGCLn4JxCxvDcOztwq
DHlRq1sUeQcymi4gYcRZWr9V0sUAjtued9jGL1byFnoO9V6tSVIISDfcxJ5Q+B+8
ktBupOqSHkWIScfmvfRuqroeWPYuB/F4qa36pzfdSoV9P/p0+yZb/AWqq+fSHRnm
SxW4W6sEIYuz1YbQvru8kA9nnl8+YnwQ2gutX1UqQN6fBu4WfWSR3Ws4FNpNfUNO
D3r4Pu3X29DVFX9xGbdT6oDTRhLczXb2yPnhOz0ORaA4MoNPLmL4wXbQB4yt/+Kw
5fCyfjO7B2kCDVZsZY45u2WNUpzSLLsWyepFASqkn19d6DJDT86pL7HVfP0GSgxE
1qHvHg/wiO/QhpDLujqVNJYtz05erbNTCWJd4+19h4LEOfPX13ZfsbVcQHrUtnpO
NZpnt0+AJc/ZhfO/0lpe+J1tuK0YAOws2ApRRBgENzmYXKZH0c1yny/2J38V5Gxo
mYGH2CS4UyCQlyd/t9GeRHNaTcgZU5py9CCy7QB5S70fW5wijh/2mNgNdKjLJ/Xz
cA5TgRhy0qAjAU72b9VF5/b+WVTbxFtLbmTOj8CeTYLKJgnN12dYSxrEfOIZnBne
D8ThvT8ViyCKhUkjPQWy9IgltquKhsD3X3UkU+SIM1AEa8LFx9RsvAOdRHhRI7bl
YP1lkwkIkh0PVB/w2tE0+VXoMLzR3jjVcd3F1fKeQPPXoTTn4yeG8zQFTQjeX9IL
631IDXyv8WH6OunGr9y5cWllE+LWyUEX9d6L9WBJcVyMn0vw8bdiEDCaPX1VND6S
Hxpq4yMAQf2pbfx4kd9uV9poe1FTLQYmHeXSTOgLWSNYHNUn3vNIduJRxk4KWE+e
5QpvosVfS5UaZBl0rwDRRXD5BqrdiOf7QtdnCmI82WOqwflLhsMmtsNZbH+tzBM9
piCiOf7Gh4aNflySIFGVIn732NFPhdznfW+4w3+MXH06BnAxypt9xPd2pRo0Leis
5f2STWuTOKc0zNSdZI46VxnPXKFRoM54Mze7UDwiOgGM12qH+Gxpd6T0VHUzxo0V
EVyKPCZfIg2qfxOO5QWY9lo0MyFFgnvUSm84FvMK9JLEAgnRqhcZSQ6JQVi9yJGI
oq2M1n9asgY0PnmeMk7mKxZnOdyRckMGV1sWCWbA1l96nToHk537Bw4a+tqTtxr4
RxHXjL+fIir0G+FPVXMQYVXs9kodJWlwRqJ9xH9W2eOz2iGblY0djsdGobT6KTAx
FFJn56/5Z1Y125OygrSoXbCPvoci2/+z1nXM5DjHbGZ/qjSnhIiSQ05qd/bPUpLf
GaPG+8ISL4vX4F8SXqAq//bn4WqKwiT2AvP8Gql42cJHBh1ZYWYB8YGB8pAOn1cK
pTd5XqQK4S48W6z7uWvoaEM6SoQhxrX2njwro+FsXJIUEVjZgz8z2eN6CTtO2hrZ
FtaNmoBJSqFF9QjWjQko2sQIrvsWhzANjki/fU3+DJG5D0vBW345sm82lHJpAOGR
3pDaHjCO0yraCL6rRPRcS2Dyt4EafPBw/TJtSowyWkrs2ux1OV8ICGgvLjFqB/Xy
oQZYAZ6/ImzgYCI6Q7VarMCR7SKp9N+MePmacaAxiclCImWqVcAckmT18eA4/fEe
yU/CQt3H5sCu/ldiySBV2MRQ/Gt51ak29fbpBgK/vb1UCF7mCWuQADG38OJTHFaV
+6DkANr6Z8LvYN9ahQzbykkd7tio/P1WWt57f8jgv40nEMYLxNYGujMbzbZ3zXE3
eUtiSadbo6BWT95YkXwJb+J5iGqK9ICvqI3qZYTv0rTRaAsMrsA5EucQlEulME8K
YptF6z46n0cvTEcV6RjRyeJGja8zC0QBRyT9MVhyorCxZ/DFUsnjTxfAf7X0cZUl
JLbwJvVYSHp5j4Qna6JvvkX39p+SqQ+cPenSiInDoPVOmGdZIJ14ffi3ADLnt0Dn
C/NiXbU9JHzHrf8OZMPQ0MuMkag50QOKknQI5qcIifQyU0qlwY4aHVcym7IWCJvF
+n4+t7ABeymS4Qek8QtOhfzvcH1yEYRVjsdc1aGBkF9y/ZIKJpx5rq11UQztdDe8
cCCL5Kk8ODzbvs92fwFDYc32j6XDi0yOvBqITLFU53ut5Q6bfOhJuyUnwLr+PVWh
bk2HpMyq+hYwJItxNqz2pu+yk6GjNHyJ179alKlFLjQ4rYtimn6W+E4UPPVsQ4R0
4n2gRXO8CnxoCAZQ6uk3vKRY1gcL3omUNwG+C+zVfn6i5V5WGsgabgvbSFvlgonH
3MDHz4Mc99NP+vIXf4E3MkkPJ/2PcIVqZbZiXczGdpy7CvwkGvHIJU9x1LJrjrmW
YRHJt5BDdUTDJFeF7ALzU0QLn0UzUt08aAF2K54MtYZnI+hpoGcxX5ZvRT7X8b04
M+2O4cSMbog91LrQjH/5tXWLk5Md+EBSeQtsn9dmCjt2zINow6lj7d3rPmtIkTbY
LKgVXGJrHEhT8vEMiHN6Zv5l6ulzUpAo6IB4dmic4A4VTDmgqHDOKCZ9qoVR96jO
pnwH6SN+EMA5OXnH7Ti4jL0Bi4iIDDujg40WKcJEo3QZmItGrWFQ/vrZq+kmPV0+
f8KVixJhxuKyNBoLu/YVSNt2SAUlPmm5z0LKKJ5Uv50+LGGxSFtLDm7iD5ln8G8f
wQXnd3Sw1dVLFhmtbS3QskLJozYf37HfkBscI7m0hABMsTwM27TZmbfYJNlbIAUo
k8VRfSu7Ybbiu9yfm80rPsg1QKFy3Ek0IX2RRDKb3N19o2VyNyL+xNWe6OYcFYT9
gJruPS0gRCdCgsd6QwbbT9Pd+8OLn+Pt8qqaKBwirBw5CbRq5K+K9qwo39+v0BZ7
PaMMKoZX2xq5KLOrYTm+6QgaWv2luOCI3l0uajHPb++U8nPvubRGiSaptVLCvXUY
yFtRTVFpwtxEPJQt7zWY4/WAmBpywk47VjE1JIe46isiMyokeBIRQyyP1U0aUoGo
lFo5Jg0zo3ibicicIyk14dpwXKW/5L8gVwIhdv/rxWG9J6aiRJuiKeVyZvkyFxIm
N/Txu9RL6+B9Aawhuv7wqs7dpXc1WZZdTQfrFeMlZ73u456Gvos7EklEpSE/XLE7
R3zZu++dh8h7uak9VLuXKTPoM1MMlfqaEmMPc3BS+V8nAyuWiuTXt0VRume31wlO
NlW3GWKlrBPjxnyeGlkxT5JcJquVzwwMQ/eqiS/8M4S3YbRng0dIDutMwS2mAYAv
QVYbvQZ7C22VdJD4ElhBHn91vq2VeiIeSBzq6moegmUqHy8TtEIeUVD24twjlRJZ
zekbzMfS3txAQSr5UUoBCpihLkafM5pLOt6irZWK8+hAHB4F+2w1IqpTDWLShTPC
pzrXEvE4Aua0glk8V0I4Fa1GlV8iJ13t5JRkpCUeYHwrE5LQ1bOUwUkXTwaRnFke
GrNn3LsugUICJmAjtf06GC8pfb+/BBzTQDGImJYveqSWUtJG9bcFSQ1C63TMs57F
2U0DBp4oym1fNom2SzJX85WueJB+HxeHXvK7MyCh0VpU4ow410FADvilfPZxplpq
SEO9JscueEhOPnxwX7D8HSQz7375HE30xQ+x5CucVjn6y3TfarkaBVsPLPyVNKOk
Q0d7T1TRAVCmgtzwY34M5CXqDbVfwXBHt+RV2Qzcb2FdilgA3btvQ39LFXWG4R31
374wbcVOJOmb1e/rZ2fNtIptNawzddi6tAh4ILAbl698zokjTLwCFqy8GjFMGNly
frISCIE8zK8C7XHJTWJQtrPERCqmAzWV5vwaubK337sLMvi+iqlAPrh1RG/Dt3c1
xQ5pTNl8wwGtwJkcFcztMoBhehu8uWFhfQK5WuM+qRw/M32nBmnqudRkPG3iTgzp
menEOp8/kxljkuaOamK0RQAYv1/mGwFGKw2YiWGIWM5QU7yGZI/Yc9WLmBssCtJK
vbWJsDQNbfWiJIixccu9JiBYJbRSUiE/3u8HDBf7rPxur5lf+S0o411wQgT4t/Vd
my0A4xSCDZy2fHwZ/4lVs2wyS8G3OZhrawjy3h7EJ+2qZfKPlVCBOLw3JzIZkcPz
uVeOYyc0dxfHMRIq7edCvuYkh9CzOqo6j4cdt3Wvd4Us7JloiqRRZhbhnzL7Dlt0
+5nH/orVvny1barYRPK+wr9CAwFtmLML3oEC47aqUV2NjGVd+C/G/pWmxBlkZ1n1
TQeda6P4mI+7fdjnR9bnyPfHnPpCvcbwnHtP6ryp2T1LvxIZBI6w03G1H0qDfhCs
e9sAyGpM1YLbD7hNyym+CqyiZ1Uj51vp88+o0keSSNQl1AbBSNWE6291ynn3gPgi
hDS+xxAaXOS0xvGkUz4QK2sdQTRpHX328DBMiuknyLkTovoUI05BPLlnM2LfKD54
IHAUEgQs+fF9CVrQ0Vlje1O/bJQsxgSEfYnOAPLSneiSFhBwJuCNhIShZIdBzKMf
0xhz0mZlyndW8wBj3VCTlZmHroJXW4ybllWCFoGNI1AorDLpqhJFZtDX4VB25mXy
zSjf6/5RoQEbwmNFl7fFc0VgNe1D0nBeoX3rZM5OYHt02DSgXdXZfAcvKe4qu+qg
q7rrm0oWq/m5C7ZIzFpqubxDQzWgsFTo+t3LfU5jI+kSkSzsuN2zJyO8+RUsGhWy
J0ws5hgGcMo+kLpI4SAZTB46FZd4dHAw291c4dM1hVnDBsxkReP+EptsESBwpylF
4pLIAT7zO59pkaXBjnAddaTybf15aaQdwG91k3zPpidfX61stcHE/NOr6MQopCvt
cQDxKDg9k6WDMOvtiUymuSiHLOO7YxIpgGiH4QFRHnaTxR/VgAOQo40/sbsAzjv5
2jh2Rcsc6QzGyMqjpDWeUO7ct25pGix0n8W8g6nGg7dvSGTaseJPaWMNVnijbgAS
h9o80ZsBg0EV5kN8oawmLnUU+SjyJJ7M82r9QZi34Sm5S3BqmVSV4FXR1oo1ODbO
CrMLLPMqLj7mnfSg8VahmoJW3VtBbsE4luNEb70VinNuMzglFESq2DI/t01Tt38w
gdwiFUS95tLu2WYxGfhzhcOoaWu9RI86RD94KhtRciCAzm32O16KaEuGSJb1kmOh
zFpEwonyStpg3TapW5mX5Vlhf2tuLBJ9r0pdtSjyjxLVJF1kCnAcC31IHr2Hlnqt
FoQtaJ2s3RbpfOtwUPXfoxFwlz835dV22gluBcQitKLf33GPacJGd66DS6P7cxV+
xiNSB5CpKbhsc3b7PKNgvxgmmJGwZy787BvCsEUnj7uGLkt6+90ZactH8LIrH2uN
r/AThncpJnw1NXEOvsL6JGO//An7BDH6Vl6NwKIhKTmq7coykH+0hVX1UGR0AAj1
AGAG5KRqKoiakYBXQrTPfk26/eRCIuSM2xJhiwURqx7PvN6/bcNR+KH8PurW5uFI
xpxQh6Oq0MxYLcILlEYkGfZmbHjC3VQ+2XWovtA9ZB2ILpAHsetqTa8BQQeMxEnk
HeDNLDCQ8R2LAa4xQxE+p/NPWdl9BXrvzmOxaKIj3NzZ3FyfLzi0KwmZQv51ttfA
VHcbHFgGWsWUeFMK/AJo7PecFIaTVXSgERAeEqCeaToRMAsR3MTvMDGRltbp+vrC
QMvDeRizolfdE3oqsTdIm4nDIz/JMXhoaNhf9FgQla88PyAzEUvIwW4htXZNuDFe
0cFn/VEUlxNQ9K49TDApDkkBx7YE08p1XfEUNCy31SCttNw+NfYnU5bDIRocrbkG
jC0PrDV4NTmPUU5vJcL3xXaJte7yjNUC4lqtTGXAHCPtNJN/AmzIF0hbYOu15wFz
++2BYorJ2eNQvYDbH4Rp61gRKlpubq5s2VSYP1EwoA2Fc+VDcLxde9uX2SwD9NJL
9A1UUHH+bQzRzkB/M69fmTox8MCwynvzN3l+jQPge3xbn2vzn/pVhhmaO2iwtZuc
J2AxVtum08ZjUAKE/OUFXHCtqQiI0a8aF96jcG/uz0+H0eslSjy2ereKNWHgOMZC
Wj5jWqO7WYTFrysRabyLyrgZS7u71yjzAvcUjmzPkqLGfieyHmSzCv61GiFpcTR3
x1RFAzrg6gQtLkcJqq3SnCuXTvw+VsVoPztvkZGwv/+AL9jJEUnZVmKb3lXicVEq
DYA97vmRkGpwIQGTJPPmqs2E5HkJb2j6F1akvac8vJVlkQblBbTsG6A1+viT964Q
zRU9bJIKANYkmWtY9ndCHdcX2SK0s/15f/NcJ9hXz/IJkztIN5DPg8kF4EBJLl1/
jtBZQPUAhVf0lWeLjNqM6WJjpyl6hfu8iD7iME2Bx9vhRFsqiuaOPs/Loh6Ih0Oc
mdTMSPJ0D0Qa0POMfxix/FIkfo+MwhWe7SDumnIIk+BwGFbwGIUWV5GddZncXXeB
dXA5bATrONUI0Q5s3gFzx9I8F2Sr0xw7juieT4pVw4kIgRmhuNEu2UrX8tNIWVxe
qbMPNJFelPRsURoPGyGr407VhXhuk9RIbi+UQTZPk7prPkww4q/ClrFx+mxTP1pP
T89X9rzMA7xRivwB+QElr5uFLD86AQd/hM3tut9KHWwJRZMIvxAuWbxMK9HKJnDr
C5wUgxcxSVk4R3YE4RZURTGd6t/pTex6TMwErxodLzzdVAEO5PlYDfyZV029bhi1
TCKTJgxDeDIwtmdcS4UxBsLVhUDbcLPfQPAbcErg0y9XNZo/EG2mi82OuN6B3OYB
Bsnx8zBUaJ0kpmOJxere/pCS9dlQkbcXRTZ9TjKe0c2vdMptIzs2Ea9gZbncLoph
SPHuHOYwyeVGUH2kzf1ZFFDB3Z3HHUwZ6it4vTrHH4LxNDZGQbsnoRl+jBuzUESa
uBZzYlYLpnTynL/9nGHjXu8y7Dc6PjCWf3Yf0WcXWmRGjfP2nzNAr2105G4p3XNM
DY/rZzxH2TDRSwGxjxobqTY9URZoLFaHdoyjNeD1H6iOGCO8QU86NWafUja1tm6y
ZarSWJCkGuvxG5iKXU59naZF/2Kpf3/OFBnMEQWsvwKWkxVj6P1H7fWyowtTasT7
GwiELtvSqWGD7bSmBTU4hgnW5oxn9WFagnDyXQAvm3WAHuMA0d3+OI9rQt7Brn62
WRRTi9X9hcx4jayl9NDgD4YGz9k0lQ9el5j8lrKu4wxy8p6xXz6mf4kuDi0WarmP
iB4Ed07uGGd7FctnozAMT0PZvqzYpmHYiAaBsQAD2RgTr/EkuXkc6aMmcEJhYBss
+qkyqcuEFsnvbksyn1iwwsJYYusHGFNcsxNCroaq3dFpW5TjuLPUpkvavdnxz0In
CtzebTzRsyJZQo40yja7x07PiEIGYhZnxNnlEVpE2845TwqodpHH238odJI5z6dO
Eq44WcXY9CKBcOhxkhhLst2IHY+7ZiJ1s3UJEwEYc3iAsD/KS3WSNG9gnJRRomwL
sz/fXXzRXmBewtZ3HIddyACMajHwxE3Jlv/ilkqtJ2MLuMo0K9hYa55eVGyRjDrU
ZHLF5Rv1ck+DDGkG2rlS0ixisGxGvywSoGTeuTZGBNnclcjQwMeIZVeO5LnO36+E
w1bRyoZ8DHmxX5t9p3bmb9mdpxa4YiyMhzhnrJ/ut29BaUWz2YgmqWnZpMzXqQUJ
CTFGmTXF03YCSmgLdi+tigZuTQvvgWOflzIfOx/5IzOtSZ0VLt4QiTDmIINQa405
xOFwUiPpRVqmqFLIy8w7ooSJNEtLDKfaUwyFs2KUMpi3JoGw1ToaEfZqsb/SiCkd
Bdnn3D683CUr2kLiUPPI6jWg1GqXOgoxk5A3zkH4z/FcvDg3dM8p69/OvhnUw/S0
HdJWuGnw+F6lh0DCXsC9SeVptBzucioWW8CU77pdkGDa6LYH9R993ikHVQCYrHe1
BC/yngdO3F5Ywsdo7/oARiQG98FdRt9xyNgIEZH6nh84UhxyecFqyK79kJ7Azqfz
kI/EYQcr0QaptbysoKiNtyO+xrLmUDPpBOxIImi2MhOd1B8n1z+atZkN9alW719P
C3qQ3IVeqd41Mfa+cGPPGS6Jm6Oug+XWbMfYwPnehDFXPv1I94GKnBXLU6pDuNYp
RqkjwmViM1zI8BEMsNI5xxhoafUG1iJ4XqmoLN4e+7ax2BOox7Q8JxtF/OkTtXda
txeeTkT80/25O/kaRzXxAbZBGUNtVjfL9gHJ8U7QOarnKJkytgW/lv4lco64egXh
1Wqz9twegbm6WAfNl4ijkqOgSCcsJqg1HU9b14BCbJdMDyo7ZHEnsJu68btktWXl
vCnpMz2YpT7UenTHMJP3pmK/UavF+cgn3Qo3KWCWLds4prXZFBtvY+RYGUbjRWDN
YmFOLjVgwGBGatFHdxjePaUip3TBAY6g/FHPJX7qXiJqLKNTWo8o0Z+lSXdXXfcN
/4jRk/p0WOGrzZ94dL70xNf94mKGrL7lUQQcZgoXLIESDXk5o5fJaIIsxBsQIO/u
npgvu9KwASIeQDR2O8PMPqPpOigUUfHWiHGPerq9JgY/PANWjuuN1QANBzt+HYux
xC92jibveRI1tGQTHn6SN2X6eTmgHHSHUNKBm8xEqAkOBepJQ08bOlOTOMgW7nNS
MEpHwc5vgMUKyYeO5jLzFqqASSDaSGy7ICdSm4W9wJBMiTOOenWqni62d4D+kzmJ
iBoj098LLnZ1etOymoNO8PT1rmcGyZ1Klpx6lrV5bWtamvspgXUT1epo5SODcwTP
0LakaDKxzKqfYeeSue6QdrsMqaNAniGJO0GubmSQaRYalUko04laf9zunrGeKx3U
+Wq+8iNAh/OL+5zxGcLd+m5mdlIk9/ZVGOXOBp24TY0cTV5iGyhQi2IWmWJU3vtP
nO8kaw2hsTx+rqvAQPMIXAxaFL010OeqT6mIsTngFXfi15fOKBoK3o25C0NQbOSo
s1UlgUAOhNxFLgbbS+2+Uxgty89JhlQG2gSDHkVQ6HRr/LSQfa6AVlptNRvAF9nq
oyA/6eMBLo5UCNMyogqJTssDEAxCiU/NbKBE0oRfhLdhepFZJeCntnksE41CZlHH
3DDa99Y9t0NxOyDXDZzxWWQyRV4m6TqIVk7OKWx9en+bfRqccnPwnzfhz9qjZ5Hs
gLz3oKx2nE5duI/keJsnQ6wqPeiMKJ+eDLu1LHPzq53w7/jNGSqGkmiNmJ3B2U0W
LL8U0uLrPkCF6slVksL++NpwoPWP920cfDzdnk5YdefCNF2qJK5UxFhhmg8p39nT
mAW/SIpjX6VKoNskR0wVd2YLBpZuoEgbt/1gDXooBLC02GkEu2rTRETFAJv4LYXT
Aogh8b2A0/5qliKa+FTvX6rYjsH8DNCy3bGvmsUKoDc2EFMGT2yyIwLkmojZqh+m
hJthMWLx5PhVcvl7zVm4Qgq4x2/+RkPR/P9hMhnUdCGKl+Z1qhwbF5Ubw7xDjJJ4
Jv8M2g8hfJt/joJJU3e/HPYPg0MvxjIxfHIUjF839ezDOMsUUb6rUb0Ru+TkCvGG
XWpRy2fgpH7Xpz0woFKQrHSSYMiJoFsYOaMNtkvLkNGUvXfAgskiqG9YgOOvXH3R
E48u5q439e9GRfmDvsdhVcHHmsj9gNu741bpGks0qgItRhMH1cMxri6dj/hdC5LF
bYMaBtgw1Us5+RKpP8E8KuMjhNiwYdGstVKm3OaGeOv4OMXuqY15GTGUzJkjFtBD
/DKDo88ryDvYzGWxxLQFsbb7DUD/N3KS4cPjLLwdmn/ZT05ZO27tS2L4ljYnK8Kw
iQ916RvhmgKB2ND4A284IO20o/Wb44itnmKbV2iK5JXUgRl3m1lfmIPYUAANE5So
fZFXcCGPzDWoBuQfUGJcyHztVA0E46rMTG+dzX3WVumxv6LGCna0F/+u/R46A/zW
zjoITAmueyWl46/pZxVnB2o8++Pf6IkQhQa9gTD2NmGf0UKC6+nrolNYQWkbCD7A
ASwOh0qFhJzxI+oiCmfvqMStnEbkOYlrNO0cyDUFao4e1pyP78QeGjigJNksfJxU
sIliRldEINX8NoiZVLmEfsH+m6QgmiGRKwvso3fTpv1nCBI84DfOe++1k2QT6aw5
4qQW3RWYv37clxh6/lP8MEN/JHAW3yq81+CTkzNL0wqW3aoAs9MT4XpMl6g31v8w
pnAVvaqFHw0YZyBjkFfgZhsoava4QNN/TQEagLJv09iH8FW13EN92HlTjUlLLBNH
AIaUMbtE5kNL++LXZVQepxWiB8CrEPSMJeQH07Z3xzOg1hD2E0UyzBHmlBpJaORa
pTLEbYfUwcyaJNQUoY+HVpc1J1B0+hUtDrkcGfwctANQcSGJLpNRKQh6g2OlCHsC
ip2eEr/DcXmaXr2bZb0NxIix8J1nlf8sUDm22bcXt5BDb0//vL692btDHVCIwrOL
trB3k8c3p5fCsKH8t7K50mRxbtqLMuX+MlQrCWRXZyb3m624ca/3o1i0ooTqK4xF
pbitqR9iLSFHEF7iVCYbSBoYBDfD6t+gVaBeyp0u3hYqANy+owU5GoFJW9XkbfKg
vo2dmlJhJO9jwdWgGOXa3jpes7USI6AObrXW3Se00czkO7/qB7bffvJx7U8gElVd
kiDWNZPbXCsef0qk3nEzsYimuFB5KDlRuon924DPy83nzo+szqByepEp9KTh6wlO
6SDHDcqyLwpvfuBwdehLSQQ2ECeyO9XmWMaX3geG+qca8xr4IUbfCy08J4jPKCZb
pkT6hISzYbQKsxHgrV2m17d6VXUCubOu0hKpoBZNvLdwHu2cG4mEHn/TlUPWke2q
otsCEzy/n0Snc6D/VSQ8+yeYxsqvSxc3pFvgumerguBShj0dAALIDZ8yr2pGLMzi
PAVj6wBPYsI1Jp2+sdFBnWaATxU65InHJvV25A6JFMLNJ8dmWcShHVJrhA3i05Wq
GDIR4m6weoFXzD9wf82qz/UFGQKMgXU6tRtV0LLrLT+sVpSdb5wG2CWMLlrAQxPE
RrCSJBXaXrO/nNYtve7qPAEVyD+pGBKez+oDrA0O/Y5tQpvN3nmLAeER57fz9hZv
7fdW3elKYnwG7ndG2gO5cdQr63DpZlC8eqwgajjojkIdcMfX3++qj1RlZAufU4l/
9V9Nujprbsr+rhLmdAva9v5wem7S3sqCWLm2q47zUVUVvA8cra3cGbRNJgXzotKj
Bz3zCezSDbWIt4cTiLwVW9pSAVJLb2sIiSW6ALLpvUnLIYFpm4GqemA4GLTqW+Gl
LkZloPCg1bNvENAKA1J2lzI6IcO4oGkuDzDmlDvUCEFxs+PZ2gy3+4nw+2cjLPWx
4TwrOI6sDMlIaxKVqP3/jVhUckWiPefUKM1euNexh5WK2nqMNGaF9Rulpyetid2T
E/5Em1RmkDnizrSAeSUjGFE7Mqk9D1uw9BY1Mcvsjl1ghDj+3woD9ABWQu+iGCuW
pA7JIj673G2trRqF/fVakq8xnHTSbImp1FO+VMinfZRbd2s7GAnyVwp3JpqsgTro
jY5+Wlfq7fTeyW2I/hhxXxGlOmMzpwj0vK9bh1jgRF1Y+bWzx+iZ0UU6MYyqChNf
KrgcYAvqTt8Z2QEboxKrz2ACPqUlNEbITb5wy04Pxuj1i63YcRECPT16FRNZ9Vfi
ZKyNmTPOsd5EaIj8NNQaLY6VVZgYeTtseoF3CKEF/FvMDvtYZUU8C+/KYMXg0iXu
2RZQCqkJelhCar2Pq7W4e33dMyRF88+Kln2dTBEoEFQlcF8x5bgGyTCWJqNb3Kuz
6ZOflP5ITcIwNzsZ+CIFjvMiVcGkEdSQJD1Kulr8WLCjSZ/2TDrc5sXmNaivstIQ
hrF/0tRKghZ1F0RSbtM2qmQjoq4vrBqzkjmpiTijHDQDnySzrbPti/qAExD2jy2I
Ia46v34BE5B7ufhxjW/Gj9RVH3Y5BMG/rS1MpvE0LdAdvL9DIQJnPIo0bsOQAHl8
gfPNeRpdR5lyWl6nnCHEVTuC9ijKp8+66W3cGTHewLt3o/7gj2sgfqk41Vg2jiYP
H0ijKV+Wm/9NimA1uNkbYmDjh7oTcWc3oMWGhHOA/mgT4HCYI0qwBOXV3v3GfBdC
WsrdwUxKvb6qjz7U1y2n+SGfvusjHimjqCg0E1pPhRjHF27o8yrEDyMWWSGjone0
dwqFZdaSg+DVRVbhVWOdAkfNoEAdcMMAmJorcGXJTjVI7sohQ3l+Ru7sbKt4UigN
Qhyu5ccr8nzjshmXkvR4pV91UWIFJ67xEvsCm15YjDXMiHXpfaJ3H256BtxKJHe3
dVd4c/OAzh9HZ2UeYZhXLk2tmCFIdDshm7o7cNusfsbUezGLYWL+qHnVKCTSAD28
E5WFkpdjkl6xG+g4BuRD4GQzt/srmCsH4veatJrKbnJ0vmo2wWxhBlBtox28H087
NqkHAAdGYpSj82qYxZQkHBm06MbKlbkSw+3LL+8VMYHb0yOJkV0N/GGyPGhLtnhH
vH9fJdKeyPwbK3XQ+rhrz4p+QDRG9O+j/FSZMTAJ9oxSkNkaR6+CBeAq18aFUMay
6ku9+3m3t4zI/u0G2OMReGZCkGSqc2o3rsqUl/9nhSetFY0F+Mmrpj2UkORo4wao
wxbn7ojabgDvcu0l2vThDNhISwMjnltSSdcyLURUy7oGbO9A+ivDwooYiWZjMwUv
zGLhpZv4/U509aDi8+JRkpBcSuP8vD3BrUQu7zROGOAUYpuKJyvM8Hus2abKYhHK
k0YKoFPiHQhmoEj0MaYl686WfrPO3B7Uh/lAFFnoXTwQ+yMtv1kzGL9Su6uvGoZ6
8xtiIUdxOpHFAQ50DnogkByi+l8myQ22gW3o7o9Y3WSy3kpgMBgzPsESISFPJLlg
scOEV2oEkWnL0xwQ4jYaWKsNtzw2gTmv6UvnEV1oTCqMlpBKE7hCeZTpfpURXQG/
Ntr2Iu8bLSSz82gCeTvX4CYt6qFLlNdOZDt8k308y9roMg5GmU84n4cSRGEb/L1d
RR0ZxiZukpWPhHwMvhQwLgWAqeTXxHgM2l+9olRo5aWcCdyJzV5gX9ztlsWj4R+y
dwW0QpVA9LYG9McwoQJCqNo5m6cQfu95ILn0/bFcaZxd5aFabbZMK2xx7VkKRxeJ
LTxj/FANczqQ1ZN8jVM5QjuHnHzhHeOdJu5axhpVL4Na2q/V4uLOvmOsFv1Ck0GR
0+MgFPiJ2TqOFupcTSGqJmCWzJ6jeUMszdfsR4XAAQ1oENFPcCqux2sZ9b5gdSyK
OhRr5nVIzkLJVHSktheJefijA4ETVoo0pnWESvUAzKOPreQJJYNMw3twujj8QQal
7e02jraM4s3jYw9lhGUirz1Zfv6kNdshVEfQLQ01QDtp9s3hRpz15F0a1gwFnfkf
x7rY6tg/lhpteBAFiCZgZg4eldR9lww/3v+15Nngxkan4aGyyTK98d8dFiGo9+Ac
2gD954/ZryGzqSU/jgS1rOsqD4nCxR662+WdmK7lXAoJaaEXI/LlZkVq5IzAh0mv
Iu61KFg2Y+j6DYPn3kHHQ6WQoWk3JBYvoEkuRBKztyg6c9kwOOCdb/H2XFGweAji
hhs69753IbqyH3N9fwGII28E+K6hneEBaPtbkxoESAf989HW68wg2p6lLiBETd7J
ycwYPssxjOqjClj8f2PHb7V6cG2l/XV21+4hhXyKrKeXK4aqEKlUAN3ztIV3hBfo
Tu+k30sclNNQxpmpXYmkh2OHcSE8YSTUzr2pxN9Djh2kttuR6pb7QTLxVaoNki4O
lzaCtQBJTjrxoTXBH2aSwi66iUoGcO+fXFYlpptuj4sgLQLap+K2BKYytbBumD1M
espReJ7zFBeZdrRz3ADNkFolUK6v0ODHCJuG1kquSAbGlgm6AJ1dcmzXZYHW9aEH
rZaedRLqjsHOYMkLp/BA+sZlf20r0ao/gNUjhdXBPsg/+lUdtUhslUfX1BkzzCv/
erzzYzXQWC+yQ8Tns4d5LomTDIj+Zyn7DCEdpLlRyCRTnGlXCCVzdvG12nk+5Rbu
gjH6/H5OxBLSJajRNHyY/JtTTFjII8VCv8L0QElOfn0wm4V2B6MHbP2slxv6YEGS
2I4IWK4NT7au0bfOkq+Qrr8u5PsbpqPjJTicR5pkcfadZYpMAgIW15UApUvHYD7r
ADwwnPq95hf7NC2XrdtGUNQ7LKGbJlVwtci6bBQCeuF8BdKEy1LCGRpUwhyCTqiu
jd7pkC9ahEAdQXd0mFDoltcpXvLZmnhbzTcV1C9dnYJdWNLv0e06NgRrcYGAsWIH
I3WVzObggNI0BK/I6TuGZv63JblPLT2JnT2pvu2/x4DfN18Tyq8bFAb8+pzxC8U/
WYK4ZkbetZqNJ2a6XsgmbVxAcgCt/AV+nTFwnR9wzJdJzi4YlzQbKLbDPpznPeKk
YGduvOHoqota66myBqEkdl9UfmA9u/zo2iD1Kwuy0gBMkZ7+GEE1YOC5xkzYAytX
5r6pNPnYbgo/+7IewfO3vpdIqIIdcxqy5Kseptog6AL6VObe+5888ZXedJoCwyRm
+Iv1NrFtTH422ne7faW6q+gecvnZwyhT24gcLMzP91KyVaZ0tLfdaKp6VJxgdV7T
c6nGIB3DVTo5CCKK5N8hf4uwVfwNP9XXnZ0x0ZFC7+CQf1f04CKdgVaARsaLLiit
fCjWS4ngZcbdr54rwlMxG27Zh0ER2vVzH6LaLQAfu2mNW/b24YM8xK9Oz++eT2Uo
VXJCPiNRAJNwkfxwAMaN/cYebkSTqzu5yP40W6AfXnOVtQdOM8M5ABxfL1DypUvm
qwJf36PzpV/fDwUxu3ix2xuFkcl1u4Ug0rLmd8g0eheciuF7D2gAOENVj04BmaYd
d0Se1APnoKCGidk6K8E8sn3GyvEBXcciEPLN8038OR4/D9ZnAK2vpzD8vZ8zuh6o
G065K5dH455DI0CBpvL9K2D5P3lJXufcLG7PUiZoG81zxnL+pvB0bWOJUF8zWnZO
MheF3V1awrQXFFhZFBctnKAEUdU4CIAR0OVbSuDJqqPoUV4U1wPd5zgW2XuhEJa0
B/gdwVhEdjl2Mgt1ABW1uW7gajZWLZ3D8WdFeerWHApVJVry7gLKDJTmtrkC7VIh
ORBC5qOKp+pgSH8eqTzWkvgqxQ+hVBryT3xos2KkUWi6Yoh6HOVaDyzJhZioiAJs
NOeCgSwkKOL6Uk7yww+fYKSRuqSIzaH/jiJFwEYvRSwS2+uuq+Z5BM81GF9mFu6y
vBrNuQONubUymtQTzBv58iBdp+p+8LVHeCEuyGe6klyM7mHUALduVIad8JjcTJzV
gzdoDw7BjASOH7+aX8yz6Q7OlYZZJP8AB7BTVGEZEFUZYMzO2EPb7xIJ2lUopF6a
Pf9bNiJGtO6ASa3AN7/uf/vEkS0yGRmWVCvagEs2EpQh/qKTX+yxZFoVNfY1tXOd
H3hvelVXKxrWTQi7PbbwSxD35jgwuIzahakzjSeZ6LsKRkgR+JcF1Jr5Vobqw63u
u1c0pBLqQw9PFnnXVmX/MY5fiDnD1nS9TelFYERSeudwtgBPztFV+EqudbzbmizH
mWZfEzdYALpRri9bdE6ePqe1rRDHxDGSCzIjxjsVJXdYbMzBiF9X6OBYlFwQkdya
9HBwfFEaYHpgqCVOWLaLDtltUTAwa1Vr6JGW1EX3Z1MNcjgKn90vT1tuiLU9A7+o
3OFsbjZq3McBMTX8NKUq64kmowKOR4WjyMuGNakI3RO3kThTV25ED0FyRxLY6Uay
AqaK+Eksttyz7unWs+w/5Unz5Cub0rNlU/y1hDS/C/c+sUgteKyGTX/pZuvn0OSq
H1IoVGBTpWaQp4ve8V+W+/LvLJDCWUwg5RPVD51yQ61iqbGp8a144Ib3Aae316Qg
8gei/uWlVa99Yf46yRPIVXu8YIrlV56EYJsjU2ErYF7JO3sB7MPFjNtciWKCVEI1
gUTCdlgvsChU/CCXDkCGTXd+UPFQBIzUrcmFhsQCidPpPc1i40yQpIe/0Lm/0ZWc
5SUBr2T01COADsJTbAnyKknPgrOPgUUDYgXijqxkTssGNGm5NaAypCwUi5TW1XZ0
PZqP/6ldLmr2O2LjfgSOWB6fKgPZynPLP+fyomZh65giq3oCZsrEvMxcRtu4yvl7
NF7MgBjm4HOwVvOTaioB4KfSA6xdckInyXXPi+H6MT5XSdj8DXzUYrSPeFv2H32T
FTEkKbcHOxkHtTd8maEguGKr03O9q3bBArKoV380wCbmz+9lF0gQhYnuOqYyKQ5F
AWaGioNEzIS7pbWLV+Vvn1JwQUsnHoKvxF1FdTgeKoONbJ91jTjnOGzfDXXoSK8k
P1LeBjBLrGZHSshN6X2iGysl6W+BUBf25ylQFrlamgLX15y9yoIARdCEbwLV2NPv
q20SCXwDINEaZ4wIL/8XDfvrN2ljd7bjwrqtFtiy2ATBtfcwR+OACGVL41luIUsK
4/WLUK4CByUV7QGgtGDBQda3oeVqsyoGwldnVnG6d/JHBG1yirnFxY4E8wk0zXfQ
afJ3FbEffz/vRWO860QBYKl1mNAC/dy8dJSB4EW2tLjOqG0+015jNjfMtuvFfum5
YhAxVhP+DL0hIv0sN4lF8HhYMkChPnhbV7rRzME+AajbgLsQbGb0ZwUIt6XvSstm
By1n0qjXmyGsIeUdNeBiQbvhiS0liYq6rk83nZD9SnmHxmZ7+i7mfit6HjlxKIQG
MmjafZrWddLQ/Fdxvt+2wvHVry3Pzbt/FF4Ih7DejBxuab3w5iInl1rSz+Eo0zYR
NpFShGFZtIxWt3izFQWQmuCKICGOpvCrRKowAwBm5EbVqUvH5msZONel2dL6R8FO
QmphqOavs0uOjEA6RervSbCGpBiHzbuoBidhLtC4MrGr1QBcAjYOZIsmxck8sZRX
Xd0FlKyCl45iwL2s24abhlSB4lwgXEIduSs6JZThv7+ZRpqTlO0oFiAmBpMOVO8Z
EGE8/+6KnwopmEMWNylEF655FocdK+F00g3znN8v+nequCfw+H8rUhHCOs35WcDw
a+oovryCuABG4OFZ7mBWFfVAHXq2UkYr5V3feXIva9SwrnT7y1PQq/ItMGvF7oKn
m5RYrNIdzOLWuJhmC79FBwUBqSruiFM9zz3fady+Uhf2BXJLerQHsg7qKNe8HPdM
cqWdg0V9AB/VDvNdr75Vj6RuxwCBEMWhZltTHGJ9j0XJkElyA85jpvJnt9Sc2lWI
o5Uf/pk7YIkkvXcsjq+qeBbi/OTLl+fffJVLmtUxuvCAPWm6zHAIcbaH5YTwXTXg
lJcGsr+ozas/21b6sEbCVTtuYW8rhfN4fozEnVRmteeZDGERbFDD+awHw2ZmKu3R
UO+QjTxfrg6edybTsLCuHnEnKuGcxEvNR0IZYpiT5NSC0/MVSdadCf3Na+gRY0oa
iJgEbvg/GYQJVgtXAQG7h39eNWjSxag/CASzcvETw8IUGYgSEpndxENnRhdVUB9z
uAWjuAVNnkVhIMXX2SBiOh0y0bxOQSKK8Vd4L8N35VaYI7kg2cUKjM72B/vuXSad
GrTgnk/cWykgXF+EgCeEPoP/gIRhShx3N8XsRXLpHRKjTUTqB7kNVZtAAT3mQE+/
fRjq6ZY2Fp6cmQ4n/v3lURALXbwL/vh9ZEU4N64lys5/qprUf27mpGCb8vv1Mcy3
8i76YwPJsgM1iMokYilAz0Ual913XN/74UBLtPMqcCM19AJus/sp3tmVJ5ptBUmZ
bTpQSfIB5vmjJTjG/snfqfS6wqoopExRtTsfAAz4/PidDue+I9trsuhXo+PmNSyu
a/Efa6fRppO2yDXYaOJS/4m6JjhKvgo8p9roPKB9nqYqlg8OyqM4E6z4L/pk9qUz
jvaX+vOKIDN2ad75bdXNwVWazL1NT7DLKAnmKn2Ls+Bv89YfXbmuM6pR0TdByAMS
Olt6jiQ7SpASJziZtHuNVGTJUs1Q5PfI8bNCdtLlSFWsmYzWID5RUftg5s3DntF6
8QkIQM9y4vSSLa9i0RhUW9332R5t6sDT7xDrsXGR/NxvASvuwbqHBntdQNUNKM/C
65WMJvjyp++aqw8Cvb6kKDHGSjATAPTijUUIC0UBwz6itNPMEKrrekx0O9+6VD8H
TIyA05mG8cbdZh19N2MkccmzhNFRoZKn2rmg9W5pc4EcJJBBhtdviKg3M1YZ48am
I3Y8xahVN6uNJxdHX/wKaE61PhJ0w3dy3impRxB6M+ZMd3Bgb20nJ9fMnz9m7B9u
16ZNmg7TSgcE3xr3b60/LWbWvYIHcbeJgFSrrl9zfwSqNU34NWPfi7DZ6J5KLTTw
3BH4X+UHS9m8WZiV5GviGNaeZ49/KGD/9yAB5qBwhe4ph2sJXWRO3dm60P0ncIbQ
iqiF2H2fIYMmXvvjkfRpo1xE/+xXFg9/jgTDb8xuTFvwlBW+YGcxc8cOdmCztsgB
DfZPl8QRP7ZA6W1kEblkRk6sUuXvqDd00Te9s7xez+Ht6iNnASh/u+hJ1oqfxP7b
L7qvxo4PFw/ij1QLV6F9u8+KGhEK2uYQGc57UT9eR/gHlRuR8F2XIUTdCcNPI2R2
xsyLOrQqJQ08h1Iy5Q9q0H7rCjb4hjB4d5o7lZ+1Ob+73p6j6YYFd5adkKzLbkuQ
ezaMMof1f9+D25NSCp5zN/fLWJs3VESrnAK7uFfqpLGPLgXMiWDnQuKRWk320z4i
V+GQse6RpfP708O+8UFgwmLtoVjBeKFEd+Pl8vSu6SKFzOdSWMrRASD0TBiy+BKd
smp4eFsg0v2hddTZ1Zq2Ph2y7BgVAYkVseQTRASslwn5LRjAtVUu/eBJ/CDWK7Ti
VRg7lqLBcHAwnhUuLS6NhL7YSZfE3BUk15n9/XDyk88ka4Rc9B8MH2FE1OuPyooF
KwUZw1GTLoV5DzJ+qPAODIcopDfBoKLyoLeexxsGQ0MOT/HQ12IXBKxGDRK330w6
C3j2mBXZhs6PDmkA+6+HInBDbNzduCdx8fbNl3MOgFDb/LkrVjhd8wGOJbTxdkIU
8Qr014M4EYBqvFui+HMNKI8QHbpThKfPvhtwyOFqUsY8ZcXGVMtSDMXwS2sNMswA
sp6hfxzbRGRsQYiXMeWTZfCf8HpQKP3DLYPeLDhh5K4Sl8LQ7lF/B0Th98O+yRVt
11LT4D/zU1qFjtIczzY6rBTfJM05fkb4CRfwU/vYpyMlYksy5CnEzzDaqrhz35FU
fGRZ7AxaGQJwqAB+jvFn1ErAs6jE9ghwOUSgucjt9JuMylkcnZkdb4ocaPIaOrc+
yh/4RM2N4ocfqQFCQccsfoH6lBHswxpsMogWZRyV+cUmGtiVKtwmiTSUnd628sQx
+XZNPOr+VnJde8mwDmW+JQaGz2dFUwyUlFCHDucADO+zLBezfPwZmzgWFtu14dHB
kSypp/YC9KEefOlp2kR1o1Clp435jKSxiOWtm9hh538j3+SMqK5+6qxvHmQSnmnw
k1vcWek167NxKbqwd21pbSJ/z541fP7ybxlRY2+3i0CDagUhYnkgRK3wfP4dsml2
Jm59BYSOpugFBuSy6W/G+JuxLBoNHvsW8UgjGmlfimcLTz+6aFpjjlPsinLkTOlP
BcAG2gzomxC7r2OqNp58V9AyIO7iclN4bz3EZFXvkAfy0oPDW2mvaq5moUQh8c4G
ZIu9jzddIoa10caHC3edRLxn09rvG8QKRlP3TkqgbhExSrBgkmApLMs82fBJWaoc
F9p8ajMuqfewzQ3xAP2EVw/dFlHMQibPHIWBtjOV6ME0t1V1FRHLOb6vZnnATn6L
WKWwFexqyNOqMXVHcoQ/UkMfdN1e38veW3DIYdjZk7To5stwWzUSPht3CFSmABb0
x9clmyjoE9IF3wkBokykjM2QTmPi5JFvzRMPCCK99OPE2Ip8jx9sroSrs82VTlmG
yOHkU76wc0p1j5BbbkdAEaUgzOqnB8OvxGjs4Xf0o2xZoMKcK5v8ShAU3z73amnm
qICdVY3H0cPOGg2H01NGWtKEFqPXKpyWQPiazCMtacgAugZ9qlYR8EwzSXaVtxqm
vlfKwd58r65zHy4lpvrAK3iY6moWUonjjZO36FBM/TSuVENvK/+A9+X264lnaOpR
6v3m9kMhCzC/lGwLi2I/envQyZ6j7RVjiCfuoaO40V/Jr0vzko5tZx2DyZ/OScSX
NAlpjEVtbWvrtOivvHFCL6liXdOWfSl6M8BCpJcWEIFilTySMaV4oRXL7JjkQnyP
KIXNb8juY1BGE9MlVhJ1on55yjd5utn9YpcKLpo64jNnkNusEbUa72pkcDwXv+oQ
uXkgCZK7OL7MrVqqyxxKbXW7sV1cD7CSQmrFeCF8FMyvW1H0EmK75GD1/0cPqSKG
ACcRhxVWIpCG7nZLz1ZJzdeYu6AfN8BVCcGktNOHdKy53fhtQGwSChrYjo/CS9s3
vi7lGEULzLxRxdrUfiioH+N+4pfJHrC49LEwRg/Zrr5jXOytIUgujetXLCfyaTiM
EtowKPRiJvX9AXPNpOiuM5tNwOftsEtHI9JWUmtmTd08baKcVTnBZp2p01dKAT1j
woTNVKHuDUPNT6O2hz7A/nPWs0PRfUCsx/D3JpaHMBgretMGiimN3gjSjCJqbKjB
/yW5j96zOh+oMSfa/qKFWXw5FITEeF0qTpdFDEKQygxNxLbQsKORA2Obv3HyIumE
/tC/6kgXc8IpgjmggNQcU6zvNOLs7lmBurD8Olu+6Ab3W/Wj+wxmQ92n0JfxJv9X
JP/cixRPtBVA0OYKLjKUfdVTUZcaxQ3jU4mCkxzf6iH1+xmXgaMXSUoQcLKYtPzh
hBDvOdrMupr9eAUXWlwlo+wyhLTxBkyvYLs7aw2+b1k41Zox/Xka8h40d2tD/gW5
38lUKmzCtje1qehKKMU7+JYHjXClhQmgdKAwKp8Lb0hk0COLfrjt0KvwuHLXHj6e
UGcUqtz2YJw86tIepxGw6zQAG+CvFsXIwwUrZ0LH9/dVP48NXJKKOKVF6yv6PUqL
WENocl5QkpZC2yHslgmL6EZvIufZexInG+laM0ufIzKHpPBvRxXZUs/IHPHGlUQJ
hutt6A+sy5KOCYeOjibzwXum/naQwSy7WCidnSCcLHGdypv7ialYBFV57SrW5OTQ
cKQwxJS5K0Iv0O4nB23BbfrDlgVYjaJBU0jZ5KJnkJhXYz9zX2PfyIuQDZVRaZpA
AQrVhHL0Aw7qZ/VpQiL79DXlisUiGMHrH9ZxTdGGWLbu+YN5EBUvS7rv5IuOOOKF
bDT70n3gmt5j33tzx3ygtSv+zmOEKsCNOyLLwej74Jx+OcWQsWe4+XFfU3QoBUm2
MRnUhF3AcdSnW6xlttYiXZeaeL6HUUlISzM1aCyRJBRF09jiX1pvvYF+aeE3d4hQ
MpwhXQEYlHAzUJhuAc1HqEum3MQr0UsIkBPhH0O3dur0ouelulUOmMe1NecQbkZR
UF/d5BwzZFIAaAlEICCyi9ZCfYMC/1+Y4GVDm1UgEvFDOvhEPg6ND44P7PrvkChB
RQo5IAJ2iq7WuZWCafd0q2Y2R2IDXG0mxnJu6wtBFHCC7GhxpnfVQZtbOsdmPblI
P7HxdlpLSLHE+MTahzAYVz544YCAEkcLCubCBBV2yoZ/AWzjwkk2sgz4Y3fnA+FF
VQzyY8gOBn0b5GuuUKSFXT+d1gRci6xZp9cvlgAfq26vdMfAsGoat+LzZ/80fJp4
FMAv19y7DS1Ikhqt+JV2lP9C6YdMS5hwiLwq+0q+l745BVKqJCPsw6AkDPe1mgbY
XLByb/JfU4Wsa/bpyqaPQHaydTL9BpecYhrcs6dz1rcM54aqQ2xUBhl6CXPXDFT6
appbfAiNjKSaTdJjRIaD/W/okiXiMyJZj6C+/9XeHcj/V8Kf3u6OhwLCUbiECyau
smbem22IexhkuFuFG6gsZyux82lWf66bttZzA0PfpGNh2gQEo9eoFuvdyBZF8mRk
mzrAxaQw/g7AqY4AvdGbuCUgPEArBD4wJrN0w6YkEZHOU43blmOjve3Jn2sy1oG8
m6Je9T3wznhPrVqEHj9K+NalDXNjle1TNCyIrEa49UC/OmiiCC1eUtLolnwLMlzs
I6qbme6D+VnlgZxePopR19ModMAaoqHkc8pCTq7sWni/G5yuxmfa2olRv3DaLNeX
rcWJzMfzmQTJkaXN0n887aF0+Qo/zCoM4Mez4FoO77TWvBLBFAdP4VHox0fTBRKv
cEgJZcs+CcztRHJa76nZQkqWBmwv550TmQBK72TZLQQYvgxfEvC80DUcBxx9t2PA
eKQs+T86wpdg4Ktvq5YgpaP90WOskrg1ox9NfDdgSzMGTI6fOtqUaZLUtmo+MQuH
5caONW8J7lNTAwAwcvSWCRp4oGFATeJ11uf0mMDdvBByn/nhWhfj3bYi1+BhQLmT
b+Sq62+6+6focbgySYRo8ILpKn1rG2IB8ofWoT0Rb9wLGD881TTdqnrxQ/eIWXSX
Qk+sm0epm//AkB1UKPpSM+q2Lhd1ehNvXCQbq5/DhxfOOqlrFU+OGT91N17niyVr
RYvrZjbgWhy3bAUC69bjQGmR85NJ81eGIBon+CgGU7GocgHsNGyqFAjfnD7TnAZV
AXFd3me2o+yHKQUVNO29di9/cmYnKKmPpCLBXgmERm6TagmyrFhoELvTl+0JYx5a
F+/VORZ6TYIvaDzWCxBewazsl5QYirs8wriM9UWBnwZg7ysHWDnRir2hHZT6uoPG
mbiy2NYQhkbnEGYnIq4Cz3YZrJh8guUF7RHwjMIbWDAXgklxEBYSw+6wg61rpMVZ
7jp5iV7d/nXqKm1nom4qbHgHm9XUsaVCrNwwGYcyOMs4xaPI42c5Qnd6lOVf2lJa
jLM9bh6hNZ2Q/Z1Xpl2/ZAIkiwiQsJznrpqXIEeC8Xl9wHYg4AMBk9dEr8FA/rpu
JtgkBZw2eecgD0W+Lwv/Cl36P30Op3hXv8lutcbKl2ZvaOfDt5IVQPjFV0DkDmq/
ra/jVlTUx3N/Ei/VpepYGE5bIX+BFqMblFJ3CD9aT4cXigBCAuBj7y/rDDDu0eM2
jcqbnaSU9DNbyT67qg/UfqESxx7EpkH6/Bg6VaTInXbEeMihXpECfm9Bu6lUPtLB
6KPFaFBJvZrm+hP5tprodoVMLGlcMU505JZeUPLzFiDOAArap/qmHa7LAXL2yDWn
eVY9IREdA1EQEViPLDLgKWrLV5Z8OgL3echKgr1qwH7UzO39vD/dTT0Wc7s3dOKL
VmztwnzkCvScSxEX8VwNBnienTwtx8MwdeiOxh0CAIdy2/AETSHHbg7uV/DkeY4D
63qmBTlYarfTYI5H5q6H33n4BcyQSMpfn6wzw/Y/rE6GQ0VsBOuPldhooiWwNYiW
bAx7XPV1rD83uWI/wzVBQCvRJkPRXPmUzjKEbAVAR3Z1fN7NeclnfAtjS4MSzW9a
/hXqLotmQFUL4iueM23nRaT4Jg5cKQda9yPRn9BbXhzFu9KT3lhoSC0JDvWlYYOy
zPG1Ylk2ZmoMZo4QH1rViPn8/49SXoEPQ3mcq42BIVPXknNbCNo+DV9J6c9ssVXl
1uae6PsSV6lqthCKqq6R9Xu2JzIQd3bUS3+E49GNFaJBn7HHreG0vhrJcgz2lVCP
5FXH7DameFjHXaJHd3bNs7usCa752mUozmfHR4YNxCd0kQMw9AAb3pMm6N8grPAU
+djAICZ86kmWyZHEKc+4LsMJl6/r7FgY5IbUvk7/LKel6gxmZmvljbMRTv+YU9I3
611SZnedR3z6OSieT9zTi/PMEgGHn7kUAlDDe6QLjqDeVvqeMufUJY6FK2PG17Gn
UYOLRFoUAC015thcVv7niFDlglW/SUGyBgVeWkgJDBlHwrXn7Tm0HF/Wb11feIwp
9wkkPcvqJgbVJ8dKhO8pAht2opIl0Sgus6/sW1TLbLQxF0PpcWcitja0c4bRhl8e
jyBER6WgDCeRqpuaZvOnJta7UNDKMrIr2KbPVk+YHY/KvuNe0QT6HgVwEDCfJGPd
reERhM/nEuheLY1q6Gw8NIxfRFdfYcdzZMcKYcURV0Nd67VebYpVs4nye/FrAQD4
Bb6YZcrLGR683CqdXRBdjwnxKjgR92NHy0Xfbb3gpivAOT8wziJccoeI8Ip9oRCe
I43IkeAoh/tCQffsJ8ahowe3+xogFcyBTDcTBnCGWd7Ne1qJzTZhtBlR6IHEQi3b
ZltLiHiNIY/oqopMEC1/lcM6+KkX4hY75mOMSqBacAkbpZEtFR61AMjDeCy5JMTL
BfZR6tjv/EeHIHcFLQ8OSSSdRtxc6A2XBr0eNUPpy4gnZXv2vJy2+LOFtGSJiddW
Hq/UNf2DkrrDcBVh0KgWb4cJ+kIYUfcXTSXxDCe8SuLW7aPlqG5mPzI7a9Pkd0P4
AfJ5NyJplZPveVlmLbtO9xshskPNYTJf2A2J8ZUkL//ZQRqCD42Fz+MI8nHtgTI3
lkdl4Xaj+lbmnh6ozQto6THKUtcoQA/m4Ax0Og8nA5ukONlHXkJxYZ7LA6vtzjCA
wZGMinwJH5UgA7D5vtKwIaOySOnSo2X818vIPtur2V4m7aI0BX0zVw7O3Zf910Eh
VK9knQy5CWrsGd6R3meIMtucM3Yu45yybVNUICXGFaH9AlH46sLy/SEz/rTIbG/6
JKWXRK6Eh6U5TVa3mi5xSyelbTC9Nf3jqABfQ4/WC3ioJ66QatfLeJhcQ6Jsf7Hu
57KyE7Pl9sBFJug9MyJHMDme8wIZOzrh3A4Mm4brJXXBXieE6ixPWNQbLf4Kq9Z4
p0kAimDe7QhMciEO/zK+MeOzwfFGO/HuYKQ5coTKTdPGiv+Pdc4L0aKGvbwx8PJW
rgbMs2Eud1W5IC7jw600BpxjtQrnGmZo+CqVu8pb7uEB0pIuuDo2ZbhKFOiwfwpT
uwwtWAqmCDb+Nz4yPGNHbP4CJWioHVlYE9cIh27bcrMX95p6GsBy8t3vPgr9QjpR
EiCz0MHi4h44pfFSlNcX9HkJ9kK70LuPnF1UNYqVlu6/tKfP0W3hQRULAyj3LSoS
Hh9Iy/MVFkNWpf8SvB+kVzObNUpqJ1vtxvFCAl/ZqsxZ7kkzppqCzTMnzxAMH1Mw
nDPXtzS6B5IZGb4/ty3qOORVWeXQzGmVIka3xNoR17QBCpJylE+KgLzxeaJWVGhk
em91f/ztf5mMZGFUicUrITlHk/m1iGApRT6ZH+CQpYKKLVlUnJDt82DZNtSQI/gW
qtKdQOxulJ1Hb4SppgI0Jxlxd92UuzNq1BWkabdYom9387kXuTFkpaq2QdrvDutT
Xryv5fm60wDz8wRSi1xVDkPt9/MjsQMx8x31vygMhpGlsHeXlpgsv03Ya8/eBfPn
i7sepZNBSU0scnHi+NXi4FMKnx+POKYWsnLoVixhwcBamqKIiMAshGVRhoDJpi10
OxP42hzzDX+bSVQXCA2EmbOeXdaYFKZFS2IPrQxeQe6/Wkg8h++UN0s3x3Gg3Svf
iWFHhCV21l9CsgR2jR4bsmoVNq6pzGTJ8F7cTaYtN8UAg2d7n/a2I3UVvWUV0t2t
u7ZH2rp+vE4Aqyjfrr93vWZtdqTXwI6LrU1tsGnG3D+0k6qMTV1npwSGMcr+1Ugr
EkAgqC34vtPF3+pU955iJofNoptiDi8/SivUWpltMaV/0pbG9UhkWXcSAjQRbOCR
IQn3nqW/nfItsQxEiv733ymRIdbqaHKehir1VbUrkG7YL0hZCKlVEcgoAhygl4EZ
F2HEBNEvJy6fwMSPS+eJyzN727VcHfCt95ncV8PFNChQMV6yUDQ767M73S00R/Ym
XPwVRdQdNLGCwTrz8ozY7RUHezLAnyDyPs+fINWSK/CPWaYU6Beodmfl5sO+g+yK
DDvuilTiyrWnAlcB1UQcC/HUWPrX8xEeVISAWn5uTIP0yl9c8JHiM7d9ei1qeaXd
RbWH8UO68RzkvJai6APQkXgPp0akdZwIyfLlrLXyMUq8HmtcHwEQpdgXO/t0ryP/
41idY3PAUo2XKgzeRbyYl1nuH/PGrf3XMoPE+7npt68vQGiUg+rIXRgz5PqmXuMY
I6NV3IJVeey2DuZX/eOCmVwtRBhgJXQuDfKUNqLR1bCWlXUPjKFEOLxOODPv2ac0
/q9mr8+duXgZAs8ENY3a7oaGDLax5crtAzjI5Dq5DXK2olHDxp0F7RiQlP2BLbtL
FGO+6ERzKa1fsG1flHEnODPrCSVbpcGV0MfXa11FVcDIVECqf2b+ICXVEtRIlBi/
+6LlBWNPV4FNcQ6u8TA+hrMOeLyvXisyywBjo8p0QCl6nJV5uuNm9JOiFh0LXNcn
8QnnbZlxl3rIdX8az61BHwAB/8lPsBGu/LXk2RMF7U7lTb7fiWrgm3cpgliFn/cT
sW5wsa+OjXkQw1faaMr+x4x6n/YSFN6pbLV/osA+sFLzOrWP9Wm9JE6iE8bCU0ri
23HHusSpKPdGOS0REF2yaCM3KK31HnvYsum5/NFflnCN01jV1RQpkwdySvYOo9W8
dmulqE1+rFo0wCS2vbi37WREiKoa14dKOdU62LdaOUYOcgBQcjnvP2MquRVTWibL
pOTPte7Ezzwjp9Xi1R6PCbGC+GeCx4dueIrM4gRBR+9LSPESSacu2XDFbHvGbWN0
SEqiL/Z8kcRHchY6Dl0GOdLF8Cz+9gtDMIf4+6PQ/B6zkv+J4o2c0+wBlhrN+Mm3
ep1M9mfdtlzUojKpt3A3EOTBeGnYYgHWolzHU2eBrhSKOkUOnxpbcliKHfaclLLP
j6Yn95/lr8A8wr+SFcjjIFuaJgLKjMZdYMvzkeezpjdFRbd7LZ84kgeJJMuIDowd
91EAkmHcMvZtE9VffjLmcah/zhtRWLp4zOhMrXBP1h+2Dt8PPn5wu/8HPbB7C7Vl
PB7XWO0OzkktOoGdgc8S/Q2y1+MKVsY4oKdXmuyCMexEsnIawg8jYH7u6uuKxin3
mEdxb2fyvAVonRXVm11wprVu/XxqRxL+DKlhJZmqMyuuCMormy8fI9RRQ1oADyVt
hZJKwK7flhhV0uPZWHiBk5TuGgq93Ji6yiDS4JIButg3IHfVfWVPOrRyq+fUhXY/
Fofs5/k/ke5MGiK5AuTRGaTMR/N3Pur7oDQLYqPcTud9DnzKIAbxLmsRmairKTJh
e9LCrpL6SkPb8VGirzurInp/WS6PY+GlDJcF9VWaeBg5PbMIrwYy5yu9u8CLNqJ3
4zrq5O5vN9GDyfPFi1jqPQRCft1zHuqxouPT2TE7g3NSXLNYQKLjZnuGZo9C61rX
WhOn9L2Vf3TKWK51Mv6tyj0Qz2scSL/5EyevzGZC3F50ptjcecH5s+6HaFz3FksQ
e4Y/6OL2WLHA8+6vTZmKVbhpGaVbIT84aqXgIN6bhK4p+4DM2j+prxMCy+IOt7q/
+MgkL3NYHPxuNPIPQo+M23168Agl1HT5e2EjQH7ketRkLAWmuXjpL2gEQ8UkfGjN
Kyl5g/Wyjzj2VDbqgpuOaKTbzlvpdFMT9M6vK2rZOBV5B7lHyDADYN/p+SI0QNvC
rOe4dw5S7uF2m/AwbUD/SuBEtRLVuXW0cqi3w83xfuhdmlK2CUJRI7FymSpSL7c2
pBbzlElpYToWkENR9LLOJC8TjsOh9B9xTTQTLcYrk/CpiXibvHlnvjAsBP0oPKIY
xFleMtalJJ+J9u4OLFwfiPa5q33I0bboQiFxSJxojvt3P9POYdNhAcwJ6Tc2Lzmi
gsd6/S4Je3U4evwQnS17yBpiuFs8V69pyW4CMADVhDqV3xkG5A1iUOiwHmMDeIrA
K1DXw53HioJNxkP76lnykPrKcrMdQXWptUHNipfrPgd96/fqd79WyrhUyjRWprRJ
ZewMWiOwbyZVX5MhfTWE86kyNvZHluK4OEIwowNaSDbHAp2lSquQrJfryf6AEr0D
MV8n/tYR47rsNhLZU/XhujOqbFVW+qXtiQGbmq7bgYqFzeguWG+Q07M3COMuzGeN
djAZobUADxcTw71gS5Cm1jO+ktmyDhTTWkr0SzjLatfpf8H42fiewwRFnyGSVUTb
I6qvSu9WLheu6iWaiRRj1DC1o0kt+W53M73KBvHCfxpOW4are8kMmLg+BK2XxEy9
HHleYkajFfklNyoAq6EGXj+/1EwHYh8FvgsZQ9xa9Hj8Bf/lYVCCj78+kSRD6szF
4mbe8VPYG66m1VLkf9UVXSbz37tcJjsacm67gthOR5l3NWKA9x8s7GoZ02mWisey
DFJzH+madQ8ZSjlhNiHu0U7xfiVIxQpHVj2WrspoNR8C+BAmNkgwot2tj5WqlIW9
HNGEK/vyb4lrvWhYctGlgrB66ORyHxdl7fx9EBYOPftOAEAemngX8P5nuRqvK9U5
iLMVCDpac05CJrzZq+FsVrRtUULcfqRO3gcG1qNYc9dIoIvQA2mL9Eif8JmCxoRV
Kw+/BK64xEEhuBrs+G1H2FLoCT/tC1qsRL3AD+NqlPk7gCvlemmCWJ6X6PlLFpDz
uwUhDvya+18OK+qJgBI1bRVGtP2q/2FiDTpk6KaWJb0veCBF6gIwCX5Q4rw/0/I0
Du9R0gDdbfZW6+bJPCYP6O2d9O4SERPlsAQhWbvG9p9Q/AQHiDUqUdgeDXpVdP2h
tKG+AvhXLORs0wXOqRarqWWqz8xeX3+OGi+4/30EVmm98VyXNjKo0FVOfRiHQewG
QUqN6djC511TfonhzSFWaCWOKLuiwBa5VMfntMUo2ptz3Xi+VKMrAnW56mGA0gQS
24BiORLsVVCZ74o9EO3DEZaWjA6bIzQgM67FHtH2/JLmWf2WTiykkjJ0+KXcZH0t
1DI6tvZ4nQn9BWgc+AECLILIuOCfVmx8c8ndKYusYFsR9NEhW/8vwrQRLIw+PQqk
aWE5uTVX7xIqIj5pvh5ETUfp2KKP3RYjMwGKdzkBn8jearsvLNJMZ7/sIFeLYV9f
c7DXKv9b2y6wFWs+I2bOzVHZMZGiO91tJJR45tJ8SeWtphXaXdtFkOAqdGBSiwrW
vADAtWFQWQE+0BiBPd/OOpmO82MLRwnNYvdPv0fH6jKbhyuGb8EWrVAjQIbjgZ7O
H/ke3IfRfVF0DP3/Ib5pnbdOQUrEmSRIu86m+Lj5bMfoHz7n4cTL0HafdOQjQTl8
cp3SQci9D7KSSWScibfgRd2ubtocz75ePf78FVCvOX2thUVE25w1rQMpcPi3aNy3
Fs+Obv8885CqrypZw7SRziP0ARuKlRvmSe3qkG9RPg49sYiMjHzo0Uujnl+iWrKY
TqlTbx4wZwExdFM2+vlVcz+8yUGl4QTO9TKlpMZ6hjPFJOrWLS3V1vk3mPsUWDxI
/oC0DeFrKjCD7Xw2saX0YzwoaAlDHnncuuggFG5eRp2vh/ivuEGKGOLIF6s1gcdT
eo+7JYiGTnfy3mST6QlT43Q++6Y3OH699t6htQMjV1nxnrulvBW+ff++bdJCCRkN
BmYKZAO2EwjHn3FBQQtN7KaU3KwaV69f5+SKgU+GIk/y5xPYBN4hXPs6HPI9Roh7
0dXrSJEAIxwv43qUacJ84JbtbaqL3kJGC0ldLNF6YBDZkm/BjP5Ie6XMnAKI6cPr
L728Olp1LjW3bQT4OiXYIpVxcdZHonx51W5XbIzGU3XDdzc7LnbvJHxbLORVANMU
cv0xtnl7zF54lnECWb+zYQWARPNljFIBwx+uxQ2nc8MbDNT7bmqlACJKNTcsTKSb
mc8cUluAjd6nDc0Hkgub1ZSMK/bHsnlSUkNFL+mhgC+N4qf94jIWiuPodfliPCPq
kmCQP46LB48FAGphRC2JWQAWzIqVdOHhriOdGXWsAGrwR6jX5eh5ZjDachht1kCZ
7XgWR8IG4dgt1q9G+JGEAbo/xQSA3loY0lGRNa4F0UHfajIy+aSmxSLFoBX6gTbZ
pfJ/3R4UY5DTLSerlWerYiFhuLrxHWoYwTcGLD+7j3ri9WE6y6ewqxTAtQKO+o1V
cBtTW+Lt8CkvHM5+YBXciA0xs0zrgHfYLNq2jruWwgHF5KGEiJjH3I4rxrhPQ1g5
WUDvAncyGaEBtiXnXFpVuVjnIW8VosVuOWLHbb4dZC+0Cj/uAQYIwga+i33Cqzal
zua225Pk9EhHzBHHYYU1ObzD6/4wzF8fzHhNuePx36BiG8jmS62gkIyDdHa4AMLd
w2ViJ9tw+qF4DnUff4jUqa3vG3JBw/KMsEjjCkJv1rLyOH0flYJHSq++xM1F+9+b
7VKIsG2FysUDd7Axqrf5IAHgLwvY+jKPCHMBIQDKC4Zam62ZHrt8PqEt2ENBKOAu
zBGd0dA70BrmlLRdJDQvJ2AWbZEqxmoqJOUx65n5B/GEXabImo2XRPQC1khFnpNE
7m0lgePnMst8k66gCgXwzF03E4IJx1teoTcU/uAZnXz9ADRfo55gkkZK4oo/XkvN
ZWYi9M/5/Rt2FDIquw5nN3iclOekJ2AxT46TCsT6viMKd6sJTIjP/7RmhHQql6+4
HLaGFQ637xaQel35vspi46JCWkuEKgGKyxR2TwYpuvc4Gggw/Mc98llA/jlTaJS5
A8YBj0rsFb4fiTUw/oqEabaKOVDbGYj5GQ+ZeHgQSsk19ZTjFIhAcLNo7SBRRUCD
tFFz+64Cjo2l+xCTRuSJcMJsiLjeNRmMqCOcJ9vHewYg4VFgZserPgPkiLfOyTzx
wJd1tJlH5mSFZmRkGmB39Ch0+DwRaIq/ATiOYle6VUKpcImpIEw5x827Td5tJnAs
gmJcXbD22b/4rOL9JYfkiGpV12e4hWJF/IccgHypD2jHb+6chlsXtDiZJ3pJs6PR
UF8a/fP9cUD2zXYMtrIcQ8DynMYwweSTU9C5QuAEYcpwfw89tj0WPcBupue2mJMu
qk2tVrFc4UolBnNDHlp4U8SbcJg8RaV46E0MFf7kG+BK757BUPMLHKPA7z8oYQH8
gb3LGPNIJQp6fNaIblyZ2I4aJ9qJhbztYxBTDONApE6XkrgzH0YwH0Qkep2DsO7x
Xc3PSFUnVJhFOTS7i68LdVUjgKClXrQN+jY0os7HKpl3neSG/759z23u/8tIlytx
OpMHzU6vvn+jO2RKNBW1EdclnQndVHC0dzS2U/6TEmNBZlZM0XlAp9/gNqqSiPAT
FQsZBOTW0fKjLONrWGIHgXxtELnqBGugZS/DYekuNvF5eyPkozX/DnoXaQifqRBo
DUrG9A0YWkIAOLR9lhj3RsaOlercZJ3t/ZkVPyFC6qentacWYb+qXamuRV3trn/C
UZYkgjamwaLi4uXUib/rnhPsg5LMOo8+Qs1fZ6ml8l0zJK8H1biOswICPixgM0aP
oQKpkFJjwKSJRhCADYPsv5/DK3xEX4dI6/OlwIfa3HS/wfhtiZTYj+muexzvCu7v
YwKyHcSZklm8WR9KAyfZNGH60d3kYBpzGSxV7ToqZU5fE/4AGjDP+SQ96roNjSam
RXFuzd2U6qHUr0v8k5hIcCZOhMEvrBSHY9rC+9Ie8oBQC0ByvCQkVZRhuAcVc5Ne
cSo846bkCwB2XxwalbOm6K589UgFCZfdwjjxzZccXgUxeiem5/haaYiib0Ad2yQK
Z1bEyIzhVMr6IR+sjcAkIeSnttRRwKdFOcLUJa+ZtpvR/fCJWx1MqbgAmJWVWwOh
9ph1MFqobCiOGv3V9b9tM6ai4W+aKu0Is4hVIN4vTJwLClFo2/p6+KLRhw0TLHUo
dvcUzk0CXRvB0Y6JtPnt6rLdCygDUq+fcoshQHSnJkmqZhavqdy6nBZiFanyqgRn
5w7f8CrpynhkVXHRp7sNaBGkY+JYWK1qGtBTXUt1OzA/FxbjGc41PUlykYEgjnfQ
4gkTzUI36erlymNr32JYJsAGK7ZSH/Hh7bnsc+ZRAdR09NQMrEI2ncQAE5o4XNuY
by0D0kbPCkYbI0g9hh5fKl3d7gROicp6S3UlOSBq+MEdU5tJOxAy7F+b5S4h1M9p
qQESoGdj5j4aMFuecC12rFbznK1sqFV3tQeNx/E5G0ScyseezCAVHZ8LbD8+VWDq
v92XW+eFZOo8CXxiKSds0GZxalPfkKEedFfDIiPAjs+JF1TTRunqlytpYeNUiLkB
I1pp1bNNalrwiHCM/Vxh+1Q55ZrnAOT7MQPi+8xDehVzT2bmhLcBEgx9BuApdAMW
hPVbmLG+aYAw8Nz8V8WOG8ZxBuIUKpkOq6uN8rS6OVaNI7Lj2fATJ0yu4yy4s/Lc
Xi4bvvj/tW/nOpiaiy9WdH+pam5c2iUP0tO6NGoClEzvlH19DTO0YWxtG9AcUKxg
I17PIEApUJWEARwf/MlGbnQCadLblpfC1Lsjm1vOY3EJeMekR4XX6V0WXaSq0q01
kH5lyh2tT7HEsZ8+piWrEbFfssRnR4JCgIyYjA7ziCPkUCPB5VEa8u5VmjFksw2V
j4vb8tXbud1hkg8k23oRaR6wDIEPb2LBOeUxS2tJoa1Du+OhbzXjoiTKPO82BKav
mHSTV+NE7CILQIbWhQEmaWCk+5AoH9QuKF+F6XEU+SQJHrlBES0hFiBGu6yh/oIG
LVxLDbkkJFFSlvSAgXlSyhiByPlyTXp4GtCbJjiuwv7emkW7ifDW7r1CQhzKJZMZ
AAgYNsb3I02dlgnr4fzfI0DgPA6Rvv0+lAptQpokDtJq1s2kDkkQQ1pdUBqKQoR4
HUa45FBg4NMxovv97jaMGnnB9Z4lbwiunTPX/HLN4hGtxS+N73UxfvONkrAEp3Tx
wRe47NdphZMZ70AaEvWHLkkg63pXesuw69YgKGNHZ5kFEzKTtWGlThDNLPcwWH3E
yARbODiE7YyRiB7nC3D6CjeJrIw71P1TfZHI65wt3tcZgCkCkSJODlDysGJt5pbJ
cWa3yh8BH/OwdbhFDqk7lnir50vgmi7DAHKD/u0FoJ0PuCKj2XZSajWX6GPuxj49
Pvcw3+QSNMiaskLNfpbKJN4uDUdJPUYvddtN2EP6Hxne79RDtKvotHDqXyGjpqsv
s+a5OSi8cgIeCrXDEYP3ZcTFhPKX+xDxAUy/4imWxlu5g7SOJWY6WRfWi48QLdsO
ejMVmn+YZzM44ck4Vmta0t05whlVR0qD25ccfDhuTDgei02jy6Fq8PmPznsVYmYl
vb82E9TugXRiWwIxs8bRLvdqMetjee4poEnoEMGBpbgiRmsg8cr3ogd3NjHMLZuJ
bEB5okrXtC0jtFmTahyG4Mq6CInMTCSA+QyVLN2Iq1xfjx0ihjX6Cp0LRl8M//N7
NTF910zLOIgsr+qL584JERjBnrCjcWwx+gARg7YcPYM5cn1PbxAeqARZnj0Ej6nS
aChzPuyJY3EPAJeg7DdbDEjozs9QsbUZqEvdsMl8EnDgK+OYm+lxWZ/KciiChELv
rGGUzen3zaAyHueJtoPBREP2IbZpjpIwDddodMEz72qu7u+7UwXlj++G+SOeAXSo
nwv0B7e+ofVZEW2w1ecXoyg0ouwoZ8zVa77HxnKoZjhdz9QtBnhtcUaaZ85fqPzR
DzmvKOCmrU1VkTVXVW12+cayQO6CZqX0eMZP0H2bCxpXI4/eL9iMk+xH6y7YZa5B
tRjl7McxDK1rM/TLAtkFAOME0l5jisX1aK9HVgbV7FZqEBtg2Syt3FQyhbb7EaKb
j1A4wQCLzMG/VFBsynO6Nh00Ms8VPeVS+4/Wx13bNewNF956PiEbPzxpVSyJ6pLu
jpDGHR7/iAq+ZcFus3G6IvQGjEyvxEcctwD5488Y11d+mjOpY9RNyl4Vz9hU+MmB
cAtUZeiljg1Z5WuzaLSeQVBbNxBUC12GoFaGnK6/g3T/tJvNhhz9cRM9+wMuvyA4
J9NcZrTwFhCpuwmqkJCQk2JyU8nh3+n87nBoIE66XVs3o3RJoztA8XngGO4gxnVn
CaiRdJznwq+Di8FHoAPP3fBBzcNyPRmNmPmWYU/5mM0UZmW78MCCIKKYp700De5O
O08hYvN1+ssInFTIjWuMfemXlVdl7aJchNCt2gGvD2KwNKOjOPYaBwyEiqUyzJv2
nufi7JY35OjvSQisHWjC+y8fEOO+OXTkHNNuGVeIBoGguWhf6g58NkINt/2Ap1/k
DAPpoFHFWywp2idbaUtgOS+QARypOP1ERbMSIadhd2h/w2VxClBbz5KsVvxdDbnz
TTClu910clkZ3/OHDrdXFG8fEIbwMKiDFG4M2JbCIjtMeu42rym49Q0S410Fe9cD
ZxE6GlZD4+/43smFHXxkBjRAk2F8cV1I55BqQ0ou4FgP/BPy8wbFttYp1FVgvt9m
aQHDGQku/aWzqI1OwGRsqH8bEMAg/C1u2YBbFN8a5EA0BZEkKdNwU5WGjuCCuih4
G73kL9Qd4YA4jMhwlM8Bubf0YN51VlL5ktaMi/QImuv3yNfwOg+kPVlehZyRfZ5H
B0sviKW+iOLe6fcKrsPunQIAxjbrYz3+H4lzURh7M7ZeVHiwzvmKrl4ih7emtSfZ
YHE+avaIZuUV13uPIAj0h95CZrABGylCI7AOOTYvPaTocIuF0dugQkPcmM/9p/q+
KhUM/s5WJP6bD0/6BVHiiH1icFMJyTvuzCoxI832qtUvKN1c0+yFzqozRiJFH2vI
sUtPlaXyv3gq7/bGgHFpwh5RFY+S++QpHdA2GF3UDpBoG93uzCI13V8qe/KnhuY1
BzOeje0lnHNlmC2mHl5u2onPFQz3TuLZB2RIxityEZwupPxituNJ45f+6Xo2BRMf
UHO2gg939kvSLa00UVdidWWHy7xqEBQ+DQ7qFnyX8PJw8j/ZiyRsQ7suWpXCMYLj
FyXYiHwtp05wK/Lj9NV6QstTDF7TaoJZgRl1raWqP05BbWWDA3tTFMch1S+ZlH47
RbbMlDVQJVSECE0Y24NTljF5b8AceGmYD6eP9g8r6YpOfQ24cW8QcJ1QMAwJVW9/
sqX1MXAMD5GinNw7khdhJA8SVRYxOb/Qbeo9TX+cPpZNM3o9bsPQTDCeQUqgBKfG
NQmT6d+KLVg/Sd3vUI2uhp43kh08JF4VBSiHhyJ1u7VmU6b0+/RE2YhCdqx0PE3u
OPPBhDFR5bOvfebDkaSRdSzy5/GAvN5ztNTiN9OEBrNCjXlHNLhQbvjhta68G9jK
3NJ12QrJjLzvEoJUqoGFyH+ZzbJ469rp+i8lknN2r13Qr+Wdeq0ehSdvp8Kdxb9R
FRJWk3qeWCavVjPc0ucFlmN80UpJ1nObk6ICUplw3jbgBdk8Kst45kVbgIPXvBVq
/X9XYr6IN9vlQA3UOnRn0NzHTaBYNwqd+XZSjVQPMhxVl6ohEOejG7mHdEAOBGBg
J13+TQmTEElhuGxDNdztG1IXVKxfDVImsRMEUStXR8kvv5LeLGZImFns6oI76vi8
zL53NTLP9HWwVgOlG1RIErtmljQtCqJ/f5VOlxosTlcPHDm/dLxjBalC89Ug/ASC
RQq5ywNy5oshgijVl2jy3pI6dTHUyOFA6ZrEGlleUCzXWtPyLOyNjXov9HaDfhYe
5LvwICHgbVRMYuFtal1VW0GDiLzVZKmsbdT6Zw2pAE4GxpfXvaJ4JDy+iP1JV3Yc
MQ15S/oR75b3ZdkN2alDxBnrC1RLRo3zfKLF1XBf6BLTZPkVstLbJjw6otRn8Um6
77u0xOJ+EWZX/CfyqNtXABNXcBwEBAW/d/M2AtsrV3/SgmJMXo9yIFZ7kVDNvy6q
mHmWrT4YAvlu6RqEXschgdI5FL982CABiBplwxZRnHrilej6wau51RICaOqfFjDg
/TMDrEhFn2PtgiT+ePxkMWfCJxqxIfYBtPnPcITSVPNd5PO7sH+l/zlYaJXzuRTM
2bRxJRg4R66Fjxw2ZUsMJlEgxPwxCPY7bcur5qK/SNTSNxsdvNnZQyEFCw7uFVoM
QLB8oUEXa5lhQTSLoVeDL8WUxZtXx7Xje6xZxLNUllCh9ODG/ZCSFgsVtmv9Uzt5
m/yzVswyMAwODA9MMRiJe1X8FppR+4NzmMF0cbnyNay2aY76VUpcy9uPUiQG8VpG
dm8Rvoa32V9xg7ae1SM2qR+5EXoHdl93E63mXGygsIg+s4Y5x8PRqXJL6FES8G7T
Y18kgcAn408dwk8CW9jTvoPcfMxzA0Osc1RBTXOUcmSCKCZ76rk9kEE+M4nwpKe4
om8Nu/OJD8FCVnXjLT6Me9IpQJc9mebL5QqH3PXwnT4Dy0P/1LnImkeFVqYef/lh
mL24UIm6SHEJDUGpiJmRrm6aGN5mY6UBaRZnnSfigM5n0fLkvlba7A3QojeZYVC5
S2R2cd5B55j1hcGGsIy9UyFy3D7zHS3RkeQLH08NG3pQ6ZnsI4P2D7T+SLhur3Vs
oDNN+VyXja3W2Kp3UCmlAqpj0wKWCQFgoJgcZ2z6dCWo06Xk2Fr3ycS8MxWkx3d9
nAIGDXpnPa/Qp17XTurAa8ZgWCqgyhORpRGM8qs2/SoeG9UxUpGstVNtpW6BtsQS
7+fSdM9lnT9zUzcoPpWxWbrC74ZqYXsLdQNcx3KdEgJb9WJzBNSAYDSqBD1jcQxo
0vB3AOSgqfy9NiC+vV6Q6bUKkhI1pD8PKRntpSQacKOLiZa28SWgqhJCRRkLE+Wz
8uYBTDY5bnkwL/sfgxJqkB/2dV4QK5539eXLRxXdMKtc+rSRmERpHpq4F9w4isk5
B6kC4a9wI/5rywFBnZt6of12vptM7PS4NuZz+ThZAkXxqPWXSrq/OgwLoRE1DHga
eoZtSnBQ4L1WJczChCS/gbU577sKrxQFePaYSJr51gRjMfouTnRtgQU13lXb3zyO
M4W5zJhs8N3RnPYDzw8JaB4GCefcG62KBB9W4YAGvBTU+C+PXpA91Fb1OcVHtT2T
ZczV9fgAMGm2ZYE2izLd6/k064fWLBErcpqiTyqa1vsj9BcfLGKaCCXNKszWO4d9
zHufr8Ce4umb00XpHZYmdvSoN2gbZEFZPaViOazwfP6x3Q01c9nv9OrAeTEzaGXB
KFdVPdEZkc4p+54I6fi4+2TDfpLFlPWIEyQ1MZa/4PLGMxDu5xdNsrJ+dltnCCos
6KKZy7iT7sioOX8wpx10sdmmxYD3QmicPHolDCzywG5jgFojkl318K0QuwqGAhPt
BVWYhpGACJHSCR51clAWqaQub1AIigKJ7Fd0WwSTrb0AcE8xdBdgirFlSYjlqxgg
8FXKzAjw0REk0jyCVocNRU4Frz4eZOQBhR6Fwz04+GnMtJaMzmxJJonVkepLOoB2
6WOQz9zGhVurASfy42EO93+hNfmyNr0sS0DwynOj2IgZ5E8A/gLQ6UVMKGTtWkOX
pfpp7k/0S4g8Iyb1eOE46jTDgpZgPi+vX1nwKTgXcFAQ+lDYHmcI063iN/Q/kli/
b1Pt5bbOX+SXfZj/Xa4Gqz5Dxh6ajEMaOZ9BQaYkIK6FlpCw1zKSGoP8t8YkfZXG
xXgjCgFMeT45Aw1Ef6JZp/7c7bBFygcj3dvvtN1zRdvhyWtU6Mx31JEbQvGvHThO
kqkgIfXYEOLLaSp/u8J+EBi7ttIp9F7T3PTPj1lqcSZgGcL9ZdLhevN+kmi4sXDc
fw+FNbzBtS88UiYvp2AcAmzlaMcC7IglZslRGWsPq/1yk4xOih34YJqG0tBqXTjH
gXAL3SBZf3xrx9Df/JhfYvdqCNJu6JzXWtkLPu1jbK5Y69+oH1d7sbJIBNZF2eBO
Hbl0M1vGs2W7QLX+UcSeWpvt70VJCixV/RXEME8N2pUHbgssdN6k2PnfeP4DSoXD
D+Rv+LUMNr4U2MYwfNUV+mkXIsmvOWtIz0Nr5UJEz6wZSb15S+CE5iy3MmdCLs1z
WitrIwNVqNxRIEm9Vy+ENWpbt2LZRaQ9fN5K7W0OzJZ4lmLINsZQVr5E3dmOJ36S
9GMpPIysFhjAeeCkOipIvmi9k1gF7WpOYY4XP5NjPg0+n3kkHpOm/FXMla/mTtbr
97ugTMdO22rajdlnxbIxVSlHHq17wsN94flojgov5Cx/nWipTGPdNRaIrTcKzgIU
KCCcchpd5+8fox8pWTBUQPg46sfdA4RwDEg8duhIUaWOeFzzPqUiyHTOLXdwUC6R
Mt/vgo6BEiK/p8yfqCwPyNMoz2hbrKnuaVJ/zAPM3ludcZ38WXed7nPTB/HLI13X
MtRbc3q+/vEPXmNzhVJVRlvOPtbgyKTG6jeb1Zf4kPZ6U709g4I+TLuUo1CY1qwi
7jfr/D6M8EP82loVbVgmPoHuBPUbv2ULgdPVRfTaEfeQw8HKW1ueXd361oY9eSaW
nJGKO/5h8pYt+I32jv66wZ9L01+vbRn5xaFU2a7bWog0wHAIh6WIKsnpnYuCJ6lZ
/YF06lmyGGQeDy+QEHxKay/RIGfvfWZrpW0RtnVijqRYDfDQnNq6OaAlkUv6ctDK
FLAqby7XuPfGMbZAvpdMe90B596ZZ00jXp4Q0Q1oS4t7AIBlFNXBaLKTl6TzzwcL
K0Q4xLjKk3SdL+dBrnevQmzNjX9mOp6VVu1346YCGHuEKfYSvTk2XoNYn2T8uzJe
AV4D3TKDRy4Iq1K8ywROdaxivXWax60gH3BkKc0TlUBtygEaXW1Wb2mu93VnksNA
bOqVT4jOVow2YSTCjjH0fjZ5fKIFOQYNwU0Ndzw0lirTLYMkyY1sCwHI6+cxI6c4
4Voa62Ve6pHUaPX2Bqxjs9UIUJn/QViZWJvnfsvskFU0xEbdEnh2WPCeZ0k5Jefp
BwcSq4Zt4fdADQotGTPWz0hyQh5XBWPHU2qRKE5VW3WwVmag1U8SSUkSOTSRTNE5
m7u4Qu3cjapt73kZMnRGdl8gIpwEecFreikhsfogb2mK0+PQWn+FPOhKB+GK89ux
tj5mXpRRGHQG1ZRwXantrS74Oue+13mQbMRQSxzDYc7Q0JdrQ2CJ6P/i3BnGy8hI
Br9Sjm1i/WUpR0m7mKGVTeo6CWRARBc9xIS6K9ZWBPc0HuYrQ/uS26xnm/KMyVv4
PmTDNMeA5HRYUxOSURyCoIJcIayNJ+8uU+WNBDBaQrjO1pUbuhN33+It+A9LfirE
O57JGIMDTtC1eu8ZujsFipVZGtR67bZ1FscZfSrwgXzhCOVEeHmxlxnLOgLCy1vI
zqzPamS7Jou6d+mu572BgKQDVPdQa7nLfuz1kJpjdjU9sircCbTZisQofLvm0JbS
SnRUKvioeNd/LpLvT4p1ZjSskS9ZNeAuyEhsoEg6GiWiP0FigWBOAfyS+YodU2Y9
gPrGZ65p9AvnLwiH45kvHy/hx5EYjPeDgSsZYVloEVcjQKBHWa7RFmI67KsdkXPc
thpi8XLA4IGL9mhe1k9Zm5y8v9uvV3fM19RdXyAhwshqtRcuEz0UiwPlc3F/lV6X
V3aA24razzFh4FfsOnh2z23Z5Pf3LkTrrGtVIGnRNbQl2oqhhe1rtLykZIJINJMq
pE33ORbCKd5XbCiasZvJRjZpTIhVFQY4uqMWRpgwm4Wht4Ob0fvXLB8gAhFbRIIh
UXNOOtGfeFv7FIkbar1HaKyrhJhKO7OUMOg0WVjU/U6Cqz1thqQNsvMtD4pfzI0S
gQPy/ahm2dvSf84lF/S/IpGSe2168EKEb6K5ccIIHp+vpsep/FYOjJld4ZbxmTBY
IkVvvOSUDYJipeqh52nQ8qdnQNYokAVvo4t/YAIvxNfiOPdpSF8YBUNKBpspbF3H
9+5z+/qSQlq97ZJvhU6ut1u/nrtLDXGVecm3M833/BX9z8wY+a+hsTnAxhY0mMYT
9wMIayC4aSp6Z44j9kk4nIpYGcGHCLYPVMPnHF9XCW4lgLwK+5RohjNqOgHC+0YZ
mjHe1fzcE2QjsUfWf0u1g07i11oEC91jvQEf/gR5+8eut60Yt2nrwD5DB9cgAEBc
GbKdx7FXDzxPvpp9+WxteEjtdFnzbszADMv6FMbMVrqEtXudIqN1hhWbD0/UU1Lb
hgAM8ZRJFsF4mn4CIguqqp5Y6qH1KQ6oypcVCajpfnaHLwV33nxtg0pRQjvM1/7r
kEJw8IYwucn37eZuqjlidVtM7T0JAaBI6uRs9qnA4CuUGAaw1Mj8m7eTjzQKlRlk
ckDv5onRaRdyrkW8n81+4Uf5WJY+Uw8LRfsCeKik7bgxspPI9YWKRtAe07shgi3Z
3bD9p9hxePVt6EWySZgzQ7fZgy8xUoE+V7QmhIjSklaqoPpgaPAB/SBuYyLQNw2B
oNyiBP2UyfWH9IHKCvKADokmFA348Amnf0um/pnPpzEsz36NsyaXqnewmyXCW9fH
JWdgKWXFNNu7hlZ5BAXW4jrXUSJSFY0dyiMteW346CZ8htX+aDyIfoXiDgE6uhAT
G1wEqdzGyjywlhz5CXhE1+HHyHOcZu24j+R0bSdUV+XjqG7MthQy1HO44rC3kkSx
5lM4QJdbtg0WuxMqHIO3nPXbIU9i8ehxCkaZq532Id0ujl6rxZcCWVTeF8Xd3U7z
RWCgcy3AJGQkvI7dY70aGZZ8z8j1b3vdaXAIGTimfTDsCy3QLMBx1VhOjsR5fvI0
TWVd8TEIkrjooWd5UkMPYYEdwFE8BV7QsRjBLhb6n3vk28nHGVtxonz2ppz0u5+R
ve5OLUPA0rHYtz2Bz0sRs0B1mitxuSV8lC+Hifh25+GtcnILSJqq/WGh8djFbdnu
g5deOU3Yt8gaZpwHFpdPVgWywz+MTVaStUhgci39m2Q3B4Fjo+I1U++mHibUvuk5
r9k9z4s+Ul4mJNfME07AGjTadOxUSHE3162QtlvpLmeo8ynGCXlxCTOqlw8TZ6de
2/d8OS4G/VR5Tj9r9CkKL07d4waCXxR0rJZIcz2uSOIPRHSGILgdNKis3a3QaeLp
dL0geeW8L36Jp62vF777AzC1idNTui2GDRseuzSc1BZot+OFDarwetBM/2swN82E
ORPeP5kM4I0/wSERdvf1WYinQW9LNkOiyjZ2csY8zDUAWqyfxuztqg+qvzE+smra
RWErh4NLWqu2JmSPameRPcYuaJLARiQT35k0hfg3hiHeGcFUy41md4MVVgGUX8mF
+utywrybg1yB/STKFDqU1TM0RqC0fS2Ktvm6wQQdI5nAwSj7AqDwMEdg/IK7vzew
q8YjMFOA835XcPatNx5SFzOkZPS9ARdGRAeoOAS9ZZHbkMpsizIahMf14SCdF56U
D0scTcAYiqasMEvjk0Jj974Kc0JxXw6kfpFMtKL0ELBJgRJn90bTGB7KXod6kH2R
KuvzAv/PTXcdzWzoehry3xnLm52jRNYA6MkQPfRGPzX6ueQzmUoMXC0MzYZmNIeG
upNSdxlcyDrRBvJ/IIJypbm6cRGBgTBW+S+5Vfg53kMer+wqKGdujFiprd1Cw8Ke
I2m42QvUT1UFKIOXK9XuQF5rk0UT9GpoGGUSeGencwrDUS17v8VoAQ+NDd2j3H4t
RIH3ZDbgoe0H4g2OF0yCI0wgjZWqK5hMf82KZ5Kdxsz2EjOTmz/6kr3aYf3hIizJ
Vct6LVmBWdx/UJNoxXfUrgeXAh+/yHvEKI56OtYYO9oDgn6s8iydur+uSZ5/sW90
MH+/tk0wXO7fHU/XwBM9LFkaqNwROG48elo8twl8VWBTQ6ofdZ4zAKK8RbQm733C
Jpnlw05IeXK67mPlJsdvyz5Rin8NyMeYMuMFRkz6ZBp4cfiTt7ZgPLLy9e9VSfcE
skV7mxaz1Q0ZFy94AYCeT0yzzMc1vk2UXvICRIDAO21S9Vri246Y3osfADQCAXtN
eCrGLJLmF9A1Kha3cycVxlMGt9AYfgKv7ybLzvp4ZhAwuIUoPIX5y6ZE+ppCaJA1
Se5qspDRvp3k8H8KtqGR0ei7Sua+8wI5pUJcg5uomuHmuqKcmKpohL+bxUqdAK7p
qLH5rkSCwYnFXIpkywdlxhI+O8/J/5w993VX27cBeKvF7kY0DvpwyD6Sqrj9SwKR
mjHf7xlJhCq5X+IJcLsILJX6lqJrRbJoPsViq4GvVAhEHXtFTeRH8ta+ROCCZLzr
DkGEgBXgrPwlxciG1REcCxVN8FK/OxtYTlXhkNX6s42OE1IkLiIyQ8WZ+tTKYpfM
I7zDU+bCU4cdntPRiB62IQ1d76C8gGWlPHftkQ8kOuNYwb3753xL+bl95ostD3c2
sDFxr75K6Xnx/rqkysdTZWpVhDwO9CAtqRTOzn1gcI9IQEmg7FASSkvg+evLCOVD
5jFEm+AOB0eQrUX+zpN9Kk7aP/JCodenLrSQBL+t3i41zMDCdAsrnoRjPcw9QJfS
EWsvWBJPKT3oMhoPn9E6GlTq/LS6LyZ7mTGnAY79ytacLOjCHFslm+IM1Cm5mRQT
KfnSl3ND3KX9Dr/2SzRIJxEmnEKIQ1252UI9DqLPmB8jt5OdBoxKBeMnb54x7avd
2d4J0sbJYK4/WQ5WyyuHK/jbNnLgKDmJEF/CJT/H+0fY+kqxxYKCZoJQDjfV36jv
qzpaWA2sk7yhM5nXDNebhTry2YWqPIc108lK0WDOaevdRJoAyaXfS0KkH9ubyR13
gibwYKgKRKDseRxNl4C4Ae/IDX80Cc6WcCtgrYuk4KbR8eEpX6U3lQhEvt5Ec0LB
s+CGZlOMqnjw7IqzPRxs2UZdfSZO43PK02VGHP/+KzF/NpQEIHqkvv8eXihY+YzD
zIFALb+aWZ1K6NQT7fNadFzoNMqH4cDfY9P1OVwfFx+eMv3kLcUyQ3DceZhJhx6R
+P09HPMkizEr02rT6xtzbJVkQiKydRyzkUQWB6bod89AATKBZGKbkCo/Rycbf7rC
2RgE77Awdhofm/fUAjhw+4yMvVWs5viwqhPvvFmRZMhgaVUUz10urCYMZgSe1/FT
N6l7D/cws3K+yqKs7hNDhoW6lCsyAAYnWfSmniAARwuqX+j72dLEpNV0+CXoNs7s
SajYGdB2FacJvjWg2pOjTbGM2TXBgU9wCktNZKr0yoJBsX3xR5h6u+q8tblLQCRG
9QaKeky2CT0dvIQbJEooy3V8dtG4kuwvLwXLS8EXf9EVYDgYxnrLO26gySoDKDSF
OlkB75GdXMNne52OQJcF35UDYDdv5No7QFg65OIeoPlGHfL7h58g2Hs4Dc71ANGh
gUxEBcK5frMp9Jj4dvMMOKEAlM2WBZN+fwj1KFTQLeKTsz6IyKRd8oaxAlLXweLt
gUTB4kJZ8stnMkICJE0/JnLk78k6Bw8Gywp56SLmmf8++y3hjdZVga406+TaWf+c
I78RnYQLfo6eM8D/GA9JPlyb0I2E61nb7MFf5cSQCBJ3t5ui8kRAIbHWUt1du9ir
UjzEK0DZz/rtN7EbKqMQid54S322bHF0ii8mt1Sb981Gb/SWV+khZvOslS6GrIph
/dIeQ68Z8dnpMCqXp+17FqQWohiMljcH8wwuTzr9e32oDr7nz0k0EQIOj+US9cNG
UP4994ooceyfiXM/GWp9Q5MGZasc0CrBmJT9lx37xalrnOEHMTdVLI7RENf7i3vk
yy75Ym/xF6Pt2MyCQ0Ns0XobYHJGjiG2Vru7aHlsmzw7Wvr0w8++tW9z/98jDqgr
lodOduBfzeiCpqAmSi+Cld17aq/H5cpVvB1X2BwwVwsc453ZZttTBx7oJuYS5Cry
NxLVl3GUQ2915rLQj4YVerUUMrLUsjVGRcOFLxkkb8mYsXnJkPL2GWUY3lVM434R
+m/g5u4jS16KiVSnZa2EANo773Td24Ou+YGiDjlmG4LDKd7LPOb4mNsjMD35+iwg
gkDzJ6YovMKrWjHMoW73nVtnnD4J4kMM/nM41HPf5I68IWaHivsBqWBtYBXraTQY
d+d9HID1eefZzgMpMCBHzowhxbcKc+6ZqXP58iDkRRd6hZmXXgoy3fHtMYBoZEMU
DQCAtG4cZLpQieSmBXO/bQrwYO5ZpZe1H2fi+7V118/pFxhrmrlZELU5FzOGYwRx
IH3FVb7HuaeFaRk0DTkq3zK3Z2EN6DUo4HKOfQFydWRMiPnIjDUR9cIVSs6bSu73
bhuC+G183amAUcvzk2ZrWmjEb4fjYED0hkMYtR8bRknZdU+9q23Rw5iqRVQ7w9WH
fv+aZ2+50RIOc+JCNmgsNgukQn3BX/RbkqPz1HT7lJxmVZrV2EhL/nTqksLlhj/7
XC5jO0RVvqYpV6Bn9u/UWG0rw3SrOZh5vM7Lz6pn2EwLMH4+i8EzSburn4/+zuiX
AeaMlDjOvMv9T64tEmRrs6J91hW6IkJsLGdDm+ut6UOeUGtYFE32h+Qv/ypmxhRg
V5o4JAh+1e1OXQZTzerFz3bXWO1tV8kB9CVVY/csp/IPtZ0Xz3GRGdOG1//deGMC
eqzQMonmCduY9TjnwaxaS0lb8KejdxUIPI1yfrKDcXRWqF5MK94B0k+WuamMrz0c
q0pAklvZr4/90iz1OO/p3JP6NGB8Ut+HPVlNwkEmbzL6eHR5kjp2nGC4FLxgLsBA
AUsLjDlhW6w+r1rsNbaRxICtAryEkeTLvOvaDBVkBGHgylPLySjk0hmhiEKM+YsL
PC27onKaerwjIW3IDDos8k5REuqP7BHJMCYoOvKmM3qAbbkZmxcU46pkRoN7WdJd
ycEFDM6ZI47MRofpsyNwI73VTgvlfT2KyRAwGYa/0sqyPuxHmuYzG8zo4/Ia47pO
NPbVLD8xrXTj/wblncXHcCJF34UgX8uV6G93AmHtBvxZBrD0sulo+J1kFRJ8WfzK
dq1bWuZke3tmgVmLcA+orSkAMwssy2f+WY1rw8ImPzASp4wTQHRqio3GVLrKOrp7
nK58OeI+rjbfLCOQTsGdN8nh5DzdEjeKiMXz6nud/91RpEQUWzvHxcMD2XrMQYod
pmawEn/gOonanThDe0zUNwxfpn/kyHCcqWHM+XMeSuNPx+NTtrrkR2MRyQpxVYkQ
IxoUhM4VXrAf6LHLGZw5ZgYQdx3wKX2pYI1wZO9od7JDK+C8iyqESdqXla8612bG
6oBLhVKIMPD0HECyE5DCrCl/00Nf2zWOh+G0mxkvosSNv9aDGBNhXrUCCjDEWflr
HVshpt0qcr5iDlG9eUU+kWR66dBwI05ca0ZDnv2h13AJyDYkrDyUS9aZB7D4+wN0
KngeErLEl6I4vFDBOisaQsDv/8TQ409+I4WxcPIGgZUCSAGvF4z9Rg23Ak2LosvO
ZCuN4skUgecdHWzGmOjPKKOOoZqd9E0n2v9akx6uicYySg2ctkQLGQCU75CowJPR
6u8jeAuk+Fy0TTuQQ7i3RreT1I6oxCCNsGlDvgHaYkm297q76JqGsgOn6CSUNplS
xoEQ41DhkgMNvhxsy18Sxpd0dPu/rD8iy/bT4G6OT201NgXYE4skW4GB8p2jRUWH
7Jo7JgJw7vkVSE0OzCgUAyGPYEyUtHVXli9NXis3qv6olxgkAyYDubAx6jq/qbqM
ZKHoSzw1VTatHDKwhRHy2Qh1yXLPbzbRoHSyiJzC/i8nbkGegFh80tUbLPkNsa5Y
zdJ5DHzWu+M5/OjtNSNIS0yCIDqmc8XX/Ip9f3XLVx7wJXBPOsHC62pVnpfj2hpK
gEJMZeYF0ecFRbKiR2muaTi4SEhJarKAlmE0skOUHTzj+hrnJ4lbc0Pqs8fZL6ku
qlPh1QOAYQun4E1FZNl8NKLjpBIXPIsikOido94lPRsCAu95IFfx/MNA1w/nOup0
MeiSvQlkr1G3Hs8+AnVxfrKLKuF+1VoD4dXhnsNQeaRn+06HTGafsQ/EMFw06+aq
eJ19ETe6mZUKLhrpH/h53y9Pyeaui8C1ZBvc2oq4MgKuR+fwPx6PLiZhek2xhXZl
V9nhhaF2sPGBzWBVt619PgXiFs2YLI0/o3b2dy4KDTw9wofs1oOnW1VzUgd19Ad8
wxb3MtPsFx9PqC59QNI5YJQxEbz01fI5LuOKAgV7AUjILd09seTI/tUmddlWU4CX
c5nax83MO3swYy3XP65rWetwg2MIDcq1XsUGnEJ8n9TqiX7cOO6o7VNYsVuzOb7h
CystOO47oK8y54BK+CZLk/BToOMNrv370YqrTNWNUJLK7TN1Cd3bdn+xssiTlQU+
baohj0FVWts7GF2nj4iFyR4L9940AsKQguAj8h+3320662zo2q/WT1HnFSAYEGsf
bG6loXaHF+p3b4KrGafka/zaGBSkbTGYlOEbrgkdMSxF9ypbGx2lJntJglTOjqGF
1uaTH2S1x8E+vtW5K1YtlkosXNJVOKJAGNIfMzYgC6IGCzgqYn62nRiHJthovT0B
7D5fw/zCx/NsQUb4ysPj0qP2vdnc7kTWawZSUvHaJDVFkrsYW92brA5lCS9nVX6G
6IvoElPVEOGnj1pmFeLd5vUHNbYn7iATwLa/Z0jV0SL721hvvvGwFcunvq6Y0gTf
hiuBoDWVlr3EaBofejjHVWVDh0JMcHIKdVmFjamvLQFGwfa7tKEBeQ/XCPZ9d8y9
tDoSraBRi3huWfqYSw6WDiBAQkW4CrthC7wnpDf/stu9aChgBaHhu60owhLlcud7
Xwwrl7TIkUfNHLc87VLZRdQvMbPP4uduRpXBcknxy5VlJfhtQBUGXow+T/GNVqfB
L8hFqAXPSb1Ij4UZ7zOpqhXjLJsBCMkUY2Ysh4hM7Z99VZd/waaIZpwAtLirvCxH
V6FLVqW9ApXoGMQtC9V+3hY5AJ1gU+EQARnawqfLAaVyhLL5JKCxs8pmGmAh4GIZ
gnj7fGSv5DnXR0YS8AEDOWKBvkNs38Q0YIp26z+UwCXlaReYceBqc6+bDhxosIJS
7Ge6qZA5r6Xdq8uLNBCs9auNhQ74tJpSAx0jQMyBZIqSDoHrGZ29ha7kihA786QS
2ISIQoUyPpjOp0/rxuQckvQYDMTQt/p0x7dMSqcXsI2L/jBQwQF89pWpNjME6w65
mh2/vhvytWNOJpuoFQUTPJudLmPrsCYtgY1PAkSLca2VzaFX6/ZCZIqdQg6DbNiL
sLMfwlWblCwszvgS9fMyphOBK6UgsBgfkuR4OBFycA75MS5CkYKBNJtFrkqpkWol
KQGYUaJKVx4yU6BWfSAHlaDaqwZnC8o7uaj+r3yyxIe4qygfESf+jTw1gfl+JvM7
/mrPY9EocACEusDFQ0sZrB3lpn+sehsg9HL8G0IMCh9Moprbphk9fH4qpfetPpYY
ymAMzoFrcLjrnp4944yXKiH7KNwA+N2+bxyOEp5P0mXTbxWGWXjHceb6YCyk+hZ8
WLI4GHZkT1QMxGsWRR/1RQz4Fo/3jcx7Gmj539zy7nGCuSvAIkZeE3MhBy6Ovf1i
RSpynclo80hkTx/B9iIgmfeNTc1dKeklNjaX5azeZMIyTKCKNhRLk/N7zbpszvIT
m6DT4HBPEw/y4BuLpaAEdfSNZ2PkruXtN1D9CIWlReTgZDBN/pcFPGn89Zeao2H8
5A6vlxuupcGEH4lvhJ0yqGESgmUoB4jf0sXb02uRNlUnJuSDeQ94+t5BwriWdtCl
ybjnOoKWHXw6Rf7FT/+bC6XzCNJ9bNAhv1xGVSCOdITRZMRG2AtRiNI1aIklSiX3
Rml74E0OYS7FrukwHASyyfJj3fBgu5sZ8BVrgZtMS8BkXWBRVIGqALSK79aDpsYS
5u0kVeN8QUjBO8BqJNtKYzp8+eqiceQMKHFa3G3z6mYF6jiQmAyjE+/4tORzlx6f
wGOCkHLlQvNjUFXuEaGYtAsvgCKrkOH5Ia+uzmVOsc7wIKwXiKlHIaj+bLyXocpX
w7j8bqNrLKEOycDIZlfGunOMxuFpYqNAiQ9y0JmBVUzdFGNGHqiTw0T+6QDcDl5m
mY/2XIEGt2wBUEU12jr87OYDd5dhvWdTC3Fv2ZQHxCps5V3tfFNWkeZOsuuDnObY
VonD631JPP/URnEGvO3514xpLHHn4sDUDZpT/xaf/8qbPxAtHBwrQ9KPaPeq1lCe
D/LW4FVirjUghYHoipqkgr/ymQtUp0RoYP3vhm1U9Hv7mNcDvoKRn4IzC8I0nicF
mKGxl4omBq+zpa8bjdIwQux3fFUF3vr5+9LVTf9158an3+agaGw/XhgkRhUYgKYv
iHdhaCcV7G18yc10KTP/eM4ufMEDw/2durNeRoTBo8OoBAbOOR21QKc9bN3b0UWl
+2TjSg5ncBmYi6VlUQbmzz8Y95mdQcA/qZZTtbITjqW7wQ71TAFxtp/bSHKnsvAn
k6hy92FGlLOTirRlqZ+zOL4wcs//TBae1TPA5tRu5PCZ4dZ76eDpAW/hcKO2pGS4
PlnhF/Dd4D8JgOJWgg+HFXHI9NiWev/dXIW+9ebAHjdI+ANd2AfRV/sUOtKNsXDH
yyYRk1dUp8O5RCy1fH6/Hr1jcwWguxJ+1/XKz7WQTZHMiW+BVWeRskWaGXMvc9ik
VAMWCAOKeBUOMNB5RszzuGcbCAu+WTUDmSCwOAPayuVMz5imiG74KeaJSNeTU2th
CW+MVWla7reBa8Igd8/ELno6NEQyKUv3L89sNZS/h7BOnYfpOJ3STfEQi7oKw9xa
34PIjfzhbzDjZOBNjbOLzPINFmpDaSzuUxD9gocpuS88GMHqi+Zd8FtVWaErLMvY
8uajtgKI4wlvwWLHWD+QYhPl7mNMXbYsZSK6rYYAGA21BaR4jEnqmuYV6rQitr6H
8rQHw7xh8K5k3O2yTLFcAhwrcNMA9rJ6wkh7X/Rv5kCuOQ6Cd2kDXikUgBuqpGtV
5AxtsxORInaeZfBfrSQQfJay5vlWc5BSXP/+9S9f8hFljXrGL0WiHU9O4Osop6j/
BlwuAuu71K5RiItVg8frIW4rgDbsr2yMb1flNgtddC51VVCFOwtYZr9gdVceLodB
IPTSO77W2UUM14lBR0tIia/PHWAvPkJSFjcVsn9UijUQkDN3lfH7CBYpuhZ73l6n
Ou0Pw4G4CdEbXJ2d6FeX/ZKhpUJHhXnMo5WGZuUKMmaNUwQ9tZUxKcOwB5yb0qyP
OOdmTjYHSNSg4GhNfSVN/aM5ive4+YIyYcsbqZrTGtFFXHqL4oTKgkzmGONY46ZK
tzQkUAyRxn0gwIlHTo7FgqtG8UH2eIttX4jigQ+JgbZKBjWNrrZzIlQFxOo++/hj
FEXSeaHg9LiTSEPJF2ig5DI7mK72O0hxPznMhC1nXcCnFep/44dWvMT0XEoGsc+a
TfwGVh8GTMdWLcSNLvCQvB3olhy36+iVjB0TQpX2gTrknaxtZxvnAXOKDzNaeBzZ
7bM94CAZV2NcT/h5sqXRxhJGz73TI1omA9CdNuA6Jcadq4L6ZZNo1gZ10eFmvhEq
JutQ1S65oadF0thSJ52oq71d+o2cRtaUK6bzD5ghaan4i0Q3bcFTGi/0u86s+Xw1
U/9wlpUqf0JAbQ1sapgRYFvJZH6PQ3DByF9/efIP/Gwd2B3OEkxM/+LJtX8gRUGY
qGRYoqoeh6FR5jwP9h8gKXNNKYGRDTu1Xvtiy+G+2yJqGTR/pcjWpsh38qwXG5Y1
UC4wOEAeLz6rtl5a5WfMqUry9PT3p6BW6ckAS5zZINQbuy07WjWvt3Ta4Or1+2Px
zH2UYXlsXyugGeJZpw/TI9/yrTRpa0VgZvrEu3PDQ9b8qwJiv4MkBfXjrueiLMKD
uyGwIsc/f+eR0f+HnFX1qB0jci+JIvogiCDrRAEbZh/mA4izaiwxuYMwylybURpV
aDA40TQdlNpdt5XiNpVktOVSG2VHNshgwtWxiRXbZREF2bl0jdndnj9qlSbXTZPN
3xYlUNEb5yUJci50mjGfiAhIt9Ofow/N5fQjJDoMJocbfzHPBatcD59nMApimv+i
05JaS1xTYHEd/BL+Ysn6drxY84oveVTjGWPsy8ZUwhP/utY/LANEGjnWFHzgbjR+
x30UXVtvcXcC4iiP/jNvNrQIEdE9cPArsyU9KXEvatZ0EM4QJTaL9qWSYyZyG2vz
469o+gBQxJY6/QUYU0S2JTZ8TgtvthGNinj96P3UVO8DMTn9EmDULmihqQ/zW4n9
aCfqldrgvZJkRhl8z5qBQif4jJDqmaqgUZzNxMzD7rsiUl4W+fd0gq1peSEORtKI
B3h4FEEuFa1p5gzs8yqKFjgd9hGasRARixiGrhGLpHBOlULX0XgazgJfbTbWUaJG
RKN7HTFlEwlON5SVM7dSDsfu8YwMJkQBkEe47VxN+tsPHUs9rG/A2swWtQ9SOKQB
GFIBxdR0l3yQkPsoTG7V0XLUsBs7N32xEXk9wcVmrXUIkAf9r2CdYE83IjlD4vnR
8T70sliLzuRx/KJV4WMO6pmHiKyy0RrbgN31FwjgcFE2DPy352quoOXYstHQy2jC
3qEtOjwH1CE96TBvJ1ADjHc0i98u4aquecgnZHWnV6iVg+z+58uX9jgHSbzQbSZy
V0qtwg331yuPVFmfbwtJ++3MkasTIAHOE7A0PCdtFRrjIcg9XNdDLwnfTjrXkgBR
Q1V3/88n1oIomlTW7TESsbbkMLIKyidz9D50XZPuX3zk07DZRJX6tzX+3Ad0dEPQ
Pql0Vg6DVB26Zo/h6g0WCP7bAX1dnMX2KaD0FF31IPe5arGdICXPOTWVlht5AaiX
ZVJqIrjeuJdWctNV3tHp5xh8pr/1F2M0ZSPX2qUX5JpGN2QHmLGDBng/ZNhCyYSF
LSRaGTVHWN+miKMvS9um/Edj2Sfgg05XjQ7LjV/j+3dV/RDenC5hmw1feJuQXDjM
jc53xWSgql1m7u5yVweN57acONyk1yOB3erhl8g8BYz/pAYzHVZ0XQC7NxpMwY6H
kJwwxkkjRu96k/W7/9d3/wMpq4trgHVvkGZpDM/Xf+8u7GL888uTivdWm+lwhnwL
EaEpvnr6VFQUhUn2gNeg1atRobREl2lDnc0IjZX0KqWbiGAcYJv+IIGFrQTcYqq8
B/dU4RFdjCS9BWkE+Bvk9WMEbFcjKSDPIMXvibkZ0iNeFxI2EAqcu0OXD1RF4Rm9
ElcGpIXa56La04xl+iXVqTAAuvMnJAQo8iZsW4+k7wnReMGC6ncNDcszyJHuOn7V
hzqVoGbTwQTbmfdJVhGAOPaoK9x6qfni7wmrFcfe7XYFJ+9RPw4Ol+YrVKl9UdLt
MiPHsNLVZr+96hICLfSwDBQYZujmLxad8lx2CqNLJt0k7UMMLmKjsS6rBmpU4IF2
XCq4CYIld6todb+KrxhWrpX7ETQpjZa+5zXtGlYVTSj3mbiJiWkyGh3BeuB3BC00
f2zcjgzhQOFP3bDI1nlb95jeP1A3/8TF3SMydVSaGczxNfFJ8iOCgmLFiRutPQTq
tUl9+Jh8yeist9kA6bHkyGXdmab68gsmZuVenR2lK1xsS8GkPsMs2ZYgGf6ssYT1
tZ8uEsvN6UOeImYQzNM9/0Nv+XkkPy0VOx6TfK9mdByB6TBqT5cWiJ/AdkSVu8Q/
lrNY06h4ypm2s9Rwmy0xl769TiZX6lO2+x30FL4PeV2QBlIGJo/NdywpEeMSTv4i
nAy/nDTwG1AaJ8mZHekAFlIPW67FBEPMBESiKPIjCyd5YZ2kgqg4MjL344UQHzMr
3SFid/DKxdmZD6xwBTPxXb0Ty9B8sqHAAgv9VSxAuVd+xItzWt7BZOrun2pAovia
NG5DVW138XTHP1yU2GMEpzyAV1yDJ/bfgVCA3JP4R+yErsRGDoMJRb38+KxPD90C
/SYSq5gVQBBvKbok/C06nx8SmAzLjC62Ybig3iH4rO9qBMRuAUywSuo+0ISURjwq
7MiZC+tb74W9LvUuwsex196HXZm3ia3PQA2Bs5WcHCXVuN7IEn+rw7b8TO1b5N/U
huJQE1KRGq7L95icBLjVu7ROMmE3UfV0uis0FrCuZIp+613OOqJEqNCSMkP1aMT2
b10y1WJdhl1Noyjb7PBGj1zf3lZDE/BY5mpYx1WA3CIfYZLT9zK4XHqg97U92blk
XqbCrGTcIrQyje26fQXrJldgdqehATp43O+8S2rIvdwcayLAlxAmyh38HYEffN+j
PB8qTXUAmtEeNupY/V7TARiNbc7+Ydbqa/UHpQqRVRx32shAU0g3q3Gsbt25t9QT
quAeCJKqhcCrx52/krdSZGOI+KoESLmUKFP6cdAxkjNGEkepBuJvoGfK8eHDhJOd
aTrv9nHTQWFyHntoN0B/76mz48aiWjpRe5i5PXuF+Q7t1veh0Zq+hIhmMY6rVxdq
XauY3UbVdO6krJYummO9iBnOPYXWl0O/ZIPjsMYrgxdCQUDpUwwwNqDCIj9PpEww
faQkw29xElvXGjtS4X4dJpCF4UqcpODcoDTvrhB1RXVTksz0YJnVewGRDZMHsiWP
PIb2/j9thGUfRGoinKYkRlB11w2Y5piFKwPwS2XZYNwAlNQZYZSwnX+2SL7dQyJO
WcX0iArcD93Z8Dgoy3QoJtjBhgjLxxDrE/E+Y/NS94GhbQ2Hv81Xpx+rMhUO7UKL
merzwW6ats18yakBucoDK+m6rMyBBRlw8tA8puRNo33ba+J6n2FCTFoMLHthq7l+
Isg+FLeonl/qXNaKdrP6+svEkYUM1VPp6FphWF5ygGOv7vymjK+NSVNXW8MZuY06
trDHLsvQKnTYgwlzxzHX/GJNkPTsClMCgiq7+t/Fd12ljEiwvnvrUmMsS07EBfUS
g4tY9t5ZV4LqsZVkJqa261FlEuhwDvXSrZyKODd2pAW2QfaVGGzy7aBZLs+KV867
fkDOEoCtJiRKvE6AOaEzGYWpaD9CoBOdmgnvUz9gsbYRvxLttTNQs5Ga4CQuOsvc
NJfpNqN0RbaNTNpjIWbg4vMYqEY14qxdrVu7kBRv7xXFsGIN2baj+xpV2DVaYHzc
qzGllfw0VZfZ9kL+s4hTgl83OJsqW5+xFSuHgH1pP3wKkkTwySR8HZ6f9xwLkGUY
Nx0jD/85RIfJ8+DoLnf3YG5ZGCeLh0OzVui311BS7tr5dJ+vS3nZJgZ6QaUlsvCh
RS5ql78/vdoJpfMlX7TOzuu8zzgh5wh1E6kFJ4mfR3u4814f/qFozperalQYgCX0
NFLGK+Bc8ECibg4qnNvHRXubv4zAcfK+cpYbbca2zEO0iVVGXEEJXefJb0Fshz8u
HPaLrcgq1glsCMr5DZPUcYdenKM4V1pIS5zoW7KLALl9Up0Uj1P4ChjJ7ecNv3mG
2XXWuwd7fw3W5y2mAZvGxcQQah1hD2mVKOkY/7a599okZ6rCytmHVuda3+TWbBHb
eSpnZGY+RiQE0N3GfZxxUQGgyyZ2wePyHxEW88B5MiSMaSigVo+Z9a/JR38ghesk
T0JzcsD7mnNl61W7nKT3Jk1lS03fRfjATD/zLl03/OMvXwsq2Zm6GsZoG5vDqDZ+
4rJPrDONH/GbNYT67FLeRNPjh+0n8AAF7S4cDt4f04XaQcPWB1jKho02iYN6IL2L
sUfvTm2ceIG4ddxRf5QtZsAnhgar0TtT/J6hQz1wE5EzwOlBh3wGScXZyesnd8FQ
+9NLVY2yB/17kG//hTzrwaDVXOJo2eSijquteTX2fY8tlcisH6/5JHPUqgOs8TQb
s/nkAa1Vc+sYEKjicz91SoQ8P4LFbW+ZVL6GN9WQg7Vug7W6aOKdMFqGzclPfgMj
j/dmkdHyJHAU8INueJzSc5g6CTxq4g9NNjkDp5HAumzrZ3zk5Po2tNyWHquqeRnA
haIdRBeVStFAkVE4LrBe7wl/QmF1MvAFN746CqSjBNiExBMK+5WkeS3sB6oBhrPZ
acau2Lvd2V7/VE82E7WP6CM4YX1zTdPHdfWUtSQzGiMDDng8VkSPPzGJH4oPJ7Z8
TnSpbZDeSV+1aS2Bdbs34FjG8WpUz6VcTA8bsPDrgY23tskycBo4sNdl2k9hUHvD
z1XWyovu4HRFT8jEaiDfuagk9fw6ShgyiBZRY5QhKTq5eEy4/pgto3kpfFFT2Req
q7S6jXMIxpflqRGljT7f/xdk28XbzDN9+x3xbQT4t3Gw0rTqMmWuFWgFiram8Yo3
umyo7hl2jpzOh+Ro0RHDrSFJRRhFmyh8zQS94Rp2NFHjQsZ2DBeYc4DU9FQSmlTb
3mB9R9VH+eM72NV8RlGPJF+k+e5U+kjxVxeHYByMY04/UDpKjFh89EO2vIl9lIME
8TsHRZURTQAyDE/sz4Ddm8xooRnmfXTdgppkfrSyB7ztlD6NtmlOaVRC/4NBGVG5
4n32wzXLRYYIzS5za375O0r1AsEZHoMoMJspoMVJtOZxd8HVjaVe6YZ+tmMGLY8H
I1K2sqvCevfAmDduDW8iNG9HrLBlwbVE7KRT8xRChvhkaYYEyQc8Ii0ltX5Lx892
P/0y21jVoec8Xp9u7yPWrrN0of0htEq4iBBQfQ76tHzsUQP3NBNxUi3jKjJiYu4s
wj0bW4OUZBXR3zmZ/6SJ2KIeo2C8JZL1MVjKCLFzIB0duxWufJT292DbAO3Pk76f
mu9mYf6vmhyhyJwNZG5CVSWyxIdJXtPwkPndhRbdHqjIPODQJ3KANIoBkfHV38fO
3Uy2kg2tVcvcNOpd9BU5idLCkE7D86D4x9T33ULGUkPeLVWpb4f44GPwdCfyxYQf
TPSSshJWeLdb3FEaqn7NLaPG0RLdDRC9v8XidL/42ZqV1jQlxsNGsvpoYVlMNSOd
3RBPDsFyZQ/ASkA02WVDl+LLySHPAOwwNx957KQC01/DbJkFLFSpkMPQDk42JXNB
/5mULv7p5a3OJaTcqIzsmlzAxTcbSvP+6vJBd0a7YRTMZnbjqjDe4lgi+kHvTxZ5
EZgN8UrRttAipLTEL3ghIBUG/Vj4lu+YdQBF1CrdId0mE4GpmShzfhn1lOud3YBe
Uu18qXdHeq5vA+vBjBX8NlJPEQsEW10RHvMp1H1P64sAViw+yW7bv416wTG7taHJ
n0KfJZo1HXefbIM2hN+nalbnGcBQDVcZFJYHoa773yw3H8hdqQQp2IL1wVDKKq1C
PR7Ni+0YeDc3Lm3RTthNCzzr8MNjIodjq5ztW4KYd/dHyUmigmnrfmJa+PXCsJ/L
jyO9WCs/ziI/tnCez5zTCTskxH57+7HlTq2+SjFLEexQzw5jl8BcDW5/+D7aAy/L
ckSa/C7pdE/IYhfoEExepMIK9ix3mN5mtQYJKi+KNedaQYNo6jvboLeRHpnqqfK0
nkeilg2tWLm3qFSNCRuUke/vysZP+9wCSVa9z/9PANdyo8S49DBksOg7QRguM1hb
23uww308Wo0IXJFoQJYXkzA5TbnjQH2xI6Hc0BhAoiZAis3/6MCJ3PgT2+wlgquw
wouaE6aRebd+8Yk8asFagYE6y9/n6nNCuyDbFX1a8qcxYgvEVtKq626K6jC7zyWb
RZxcokMmFfDh2DbKkSWZJ0Hn+vuDixnIszPI9Ur5Ygi7wTWTz101yV4eC/gThqy/
gG2HCm/G/gBXxemx91GnA71KPVystE6SXFuZ7A+dxKn1TeEAa23VE1d8+nwLeCvg
Vm7tmizYCrKZosK+h9zHFTD8nlG2oIRp+Hxkg5wiP1GW/7YcqItARH4synb3kYsE
Oo2nc1LKLJLmwRrMqcd/n18WH8Hh5VtyhRVgz6yXU4AV4/hnndfioplpRmAycaYv
uGwDLxCuc16t8ZA+sYoLop0hmO2hHS98Trt2ATnndaho4Lm5VBfeTfJZOCBY9387
FKgy8g9JoRZ2BCZT9IckEZk/ojqpNOMaS4+xw79npLsq0mrsLFGcous4J+ZerTx4
zo9fqDRSrkMr1D5qdc7IPaDvT/AdCFVBOhnpgRnoEMG8LDln+m3J7tGr3rY6XT1F
GLn+8OnXSkDdaPDjC85PwbbbOAehssoRKvVe93l/RLMWkN0CotED3w2iGdinyKmQ
9cyQAdlQgpR6sbNHFViDK6O/fECN33dVDx+FtXnYDhiKSLqdpXp7dsMoVDRx4ac1
24FqSYBE6MdYA3ZHHMSu5iw6Mvb4JBsshQ0i0orJut196jOqobNtzys1e8xmWipe
8VBgL/ay5iHoq377YjtMhQDD1dj9zbmI+eP2xD/Okz4MFmOumdqNiVMsZGNgJHhC
kBzxM7voak9mGFZs670mEkrP/nV9qOXL8fwZlTZGNz8hhng4Rb0zFvdhov6sUp0u
dbXYFxj8pcmDRTcA7w/xX/QF7nbnnbPiFdhIjD6YtnRh1HeWlc7fgoqxq+vah+Fb
GCBh105C/Y8D3m0LOL+wMGJVQOk7HRtFYle48B0tR7nFbmDYZJ3SHM5CnK18QNHu
uyp5mrucxlD9/HnO9Uc7Mr5L04I/GmYQVw4gsDM12U80BGBFm5q43rIM1j6pfrSP
Xv23bPutsQNpjRbKoELErkX+f10OcMyeU0i8awPdRMFBYtbute79KC1pla/B6cno
Fj4Z0wV+VEoHpr87N9iz+UeuVDPJBb9dhlZQbuSmPEn9PL3vh5T86KcWTHMwTJZ9
Rdu5NyjSdJWY3odlc3cuZ9wFuP1gu+dz+oFWoxcza+8EeB+n6JbuU7QdSOSBkdyP
VeHJ0Qn2cTMPN07D30KEiYyFTInW0HDmgpVA7MUWzWKLUeyCvEAfbzfuiOAt8tRP
T5qhc/zT0qKWvsTn5rbwPXouoAxPAMzedPm6Tk/sFNmE32+gEpJYdZm/XhscbOza
C5frKCF7x21PEfw3w+D1naj5WDWQjBQOBLmKBS4rnGmwK+BLym/QLTZUfDIZqyVg
8ZnI7cvq4jZMTMypyPYXlRVocq7TBFgnc8IpsjJuHAZ/ZRe1TqfRkJcigqJL2E9U
2Xrbs0sSeH9WRjWfZ6QFhBurm3kliE4VE1uGjIA4lcFlwqnHzGX+NRebcX8z7cyT
MZsZPkAx1LvoHyLrtJuuerYcpeBve4AqLuo2b+nZNbq/KPt+tMsJ7DHCqjbXuadU
CtnFncyfjCph8BA1jfKc/HDI/vr9sKPAQKOC5/z0sEGOFf11MCd0MgePpaPdOFlt
XlqKpYiGm4x48ypXSasFlDkMWoVNOB6OM1rNNq+FuhxiRmIcfWf/fKSs0BnqR2kD
LsgBZyeV9Vnc9Ycn6azjEWo/1mJfdUURwsjCsDfJ7iafjW7oy9R7E2VKEdU9ucGX
lmn2R1NKq5IpUpeYUr10yPaY90gCVwGjRMDsmdCZsJNNIAaxrgnu/tnaJ5BjVf7t
Z5M7hxMY0i/PfNQKLR1vjR0+hFEYEhw1zVgIpFfHnHe2xeJ7PUb34o0u+5MkMTDN
YH6VXE8eka65yvg69N27hq8lRl9VxPMjAfPMAcZgnef/dpDbgUCrR6MAr684DOU3
GAGx/LCrRgjVl5uyOTTvat1J8zTJfvuoWnjYqtYsqJmkiz34AT50H/xSqPCN610U
TZ4HjemwwxsyvXUCBo98scyL3Rxu/g2FQv+EGLsARhTvMkTj7N9GExVzgblIaXXl
0Uu3ktMyYp9p5HQtW3Ym9vVpZTTO0l5M6DVQQ6al7UllMidxGDe7ie3rDVGMFZoI
PcYG1O6MS8oUBlo3xLJe9rEtYO+oVh+9v6N9j6/pkr3jBhaKTN6onzSJc6AGPcZb
mKF4sNNiRx8UtiRKiK5OlDK6irA1N1vdD+w/PqE5SiUzDpXwILmoGggRoM5dfqSb
Q52Lou2LQRavEY8vQeuP5ntY97yLvC4VuYPx9w6yMaHYXbaNAGt2LDCJPUUzE2dm
Uk3snakfW3DqId9olzRPUr+ZbAZ217tVGi4YoIJmveRvWufmBXGlWBHgpKzZWpws
ob9CLu33rxGKcJsKw4TZhIhxGYTmMwuYwljD9QrD5d564OlWfqNnPG1AhIYlWzm7
SApRzhbLyKBiGaCpEOvbcrmfUreQ98TmZrXdpE9IoAbtr7GtgzSAhap9WSktmlHQ
JqVc7YsJ7m6SGWKG3M2wJflYsedpDIqmdZ5TBBgpAfiQeVrOuK3hkpDDiZX8f2J3
Lzh+Vupb3CQ4gCm7ZlztR4w4uliuSXwFeIPcgZsGXMEqNaDmkzkljvcOZERM6PEK
uMahXDCgm4MVqGb5ul57UnA8LcnynN58QyExjA5hxbqIofJF9oUjsMog1ury/0Wu
/K8ocsTuWfbTGRqiKSSQ/cEK8dI1bwSUNUKZ+Jmyy2xIj5cTY8tM9fEM1zLBTRas
3brW86//BAiq8SeTOejz1e+qzRJILufplNhR/LN+CXcBkZN3mUp4r7Fd/hG7c0TG
xHArp104YFuQdmQxNpf/+WvdR1aasqfKB9mJCBdrSNFdH/PWeJlX8Qoo7EqgVaJq
ydYEnTWq1sA9l8UAsmINkISP4/C+62G/Ddd59LR4YZds6K0I0ZdqEn03ZSo7y0yX
/V9oXreylDHbBeLtH4fN0+lG61hheTvy1NOCgCUzUiSlGfbjrSxfViF7ZuiQNjdM
kYSmHh3dBrEuoKLG/J5gHzzdk6nTuaF0y172vaTBuyOo9AHNvs/cw1kHyc0QaGQN
PHvXycZSum6N+YB5LXLCL9+w981Dv9bNKY9u5Dq5gq0nJHWRQnLQZQkYrWfMjjBq
7vLRldxihvTvhn5wG2IjkmHyYsRK2QKa2VtUQo+HtXWQxpWl4rYt5ovg5/+753/n
mBsN4t2myzswRCK+SXAb2IQBG3yUaesVVkmhqZA25xKL+SdWoz+N8iyuEDv5WnQ+
M2NhcW1w4tpydxxLuErlB6lx4cpQbHx6zLChhq/p7eSsz6ofx3XoCuZtFGmaxlkp
YoMIfWywvPpMfpJmyUjPI6pWbZIQWXYvA5Z25e6kstKTRvMa+hyaZI/ce0sCzt/H
SkYGrJhh/Kszam6rVVe8c2ygk1LsHhXQ6loMA891rKOjydEXe5SdLooISjE/tysc
Av3ahqdHoMfI7iFKD/r1vy35NmCOiFSio7dh2qh7UYBbmcoL8tqWwDuyF8Vudj78
8ayNkcX1RM9v4zcurPYHGnJtOQG+KoaNXXzNgqiFn0ZWZz6YVXAOhsL78rnMeGkR
NnTlvDZ3vIh6TOOH2SJ338KMH4uVjOfLy9FSs0Z5ASJMoib9hahyDjNHR0Q3D2wz
U5lMr81wMLul5UhBsJHHH51CWju4qqXXkV+4LrMrB+2NIyegY9ubAdtQY2pEUjQm
fknB+3W7tPaMAYat/6HNk9zYjIcsA+DKresn5zwkYQfqh5FTlTLoNKSi0Ui+kCOx
lyehEp89EWqsrzCDk6UUB4j07UsOCjDwZmptwpQkHPw47byMSDbtXJrtP9Uy1eE9
KBsJ4d8zSO5p/trozGEr145z+k+wHzw9sCIGwaxC9/RcABQTxoZiGLfzx/xmSyAC
+ihejNUg+i06dDiWjobe82gOLMQ/IUf9gOeMd3BCOKtFpxqbrDj3d9DUEMrkjXCp
zEswd+soYNBOurtheuEUqFSaxgjEiXQOTb1jQJYnLSJVGHZrGlgkrWFry6Iu9ZMa
QxLJ9zOTPGLYmMooThpu41zvY3b9qU3Yr6EXUysHmgzWyP26an9vfE859l/UvKyv
93foHbTCxQ2oH7tCd+iOSX3XhbyHUsTWeo6LcDZxmt35NA8yWBQMn090YNuVigTg
ZO+K6DkiQiAfrZau+Je1UH4sWMyrxZGhQb3OIqikZkBYO5Gqzg7oxbP/bzW7yAfz
RC79ekf74HBKP62X+gN6wGV0mDmmC9JcBWyfGf9lZTUDBy9vkMET30/Gx0qUfIRf
F/Oz7O620cT3uVdP5H1tgZfl3NSSmHL6r3juQ3SWjraiDNSfO+67wg610Yv7s7g1
zbi2SOaJOIJ6iyTBLvbQisrJy5Ad7voq0YZ7R60c8YNxwsWP+v33L/VHKGVDwNMD
tcl9PvR9jA8L6O+TI8Kz2vhzN3SOYHV67XzGHURtnbC5tzZwYnU9esaQbBXCGzza
G1Y0yyREijU95wsg7XOrhfvXSPLwbJCspMwsMs5SMl1/RNacnSHJEnZAzmi/xXa9
4jwpENCgeAQDCFEreGdufQ5cDsLW38q6znKo8j+bj2VkME3PKXlNp9W0MniUt/Sc
zlE+v5ylQVGzMzrmKn13QahJCyaojmRepqq8csp7SeqZxiRBMz10rvEazBWDLxfH
xvRnlpDlHtrDeOk/9h2F/2hAnh7TvaW88iTgUTerXDbcC4H7Mc1wcbr32wAyYQxo
mrXdlOCtz8IJvR/3dRmrSOd3tmUYM9TixoiPy0MuYvW4hsHTFUS3EUX25hD1mS+v
NrE+1wtISbyAY2HeJk1sfTwRy8yvYHHGR4OSN2jRx/AncyTpeRA3JyeZ8SFfbFN9
CaGqGYxW6VWyatJM/co+HIKzC7eIWPvb5qxPRNCmj74VXZdOV5yAXHGutrfZE9jn
P51B1KKQPI85dPDbxuhPEsREFkTjXPeomGuzzSXf95FqM7H9HcL2+T4T+FR3EsXq
o2m43AH3jLCHLFQVcePowWo4sSJxOoYe+y3WnyHSS6WaFSILHAJUZ+0jlUhEHRfM
Enf9MGLwe/rIpzyVm4psFmEe8ED6qu/HKU3ePisqGgGpLs57paYu2ABUoX2/3pFA
2x5TTn3pooq+VLQHc5yU5F4R1mx+Da1Vtyy84UUZkMsoPbKPXAZ+lC40xZCt+ojU
XFjyJ1c8Ww6C79yUvhSBQRmUZ0Wp9NITs96aCLQVKnqzYTFisMku8qZ89xsmqdz5
EvJlDnnpTO70rC3aaOp9bqXhLJ4LQ3ixbhCO0nsgAkcEDOjadzANaXBXBxDvCOSI
`pragma protect end_protected
