`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Pn/IgWp+f2vPSwB0OxvlTTXXaMcI2OHKDqvs7POkq5Fqf+5LoUh5xiLIHhvUF+T7
lHrSxDSEM0XTmxMkTYsnAZQH8h0imXJmJtD8uO/NyAVfeIg5Gf3Co5yw2Xi4l+ZX
jOuSGXqz2Bl/HnsFxzEgJY/WBRjaFHlf3gj/F3SBxV4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27680)
hEfQC6eharNIydgoRFQ8Ep6pRpQi7DJ+TzbBRQGdS3Bnavn6cwRq371I36EtHJo7
8vfOzWlPUk2Xdpmw4ngRHosOfJYduod1YRbYiul3n3hDI3d2f0GihYgZ9QgF6F2X
1i0llYIcilu5vsigecwJLGGhA0D44RqBocQrrdfL2BffOMlPKWO+vheotubDYywD
H9NDNyXg9TYeuh7HSj7BlmeCWDd/Yupn8bk5VfC8ume9scWLepVjNI+hQIFz8c+E
iF+ytJAm4SjuYQ2eyN35iG5eCr2C63mrQZYwg4zo7XR+JBDu/+TWVhUMLbVeBQbb
mt46WGXHO63XMUreMXX9VDn4qQFY75ZxdGbqea4p3ReYI+ugjswdId+2lwXPZA/h
cfHwyyxTiB48Hof2fPJcveAVJ0hxHmPHrBBeSkEcZbZRNL4Yjyi5ohBU1f1g6jf0
4ZS2G0Vjug3u7OVbxNtMAO6vcXCiuVAFSN9ScG+G5rlmdRsjnyII//xftRmwyOAO
jHaLq50WLyTo9MDTuIWqs5xmPUIx3ve03ELrazeENRIWd5gTpgWB84j2waThyim0
LyM71MAWvwu9ehT5fC7xnSiWqHeXO9Op/9h3LRYMu+yhHq8LymOD3l7dOSDNODUx
RX9/pNzO+8GWDPT4hpzb/Ex9vuWttmlbau6mZtiHI5XUmfcTOywaBP6mO/RUMTEK
os9prCChyQ2z5R/eOXkXkR+C0xibB3Xcikn3JZyPJRe2BDMdeOsrwpGtLlWLBYL3
ki7vZPc9gbGkEd6geuDriApr5H3wQ1Gg3rOAAY2wERcsep0Y8TpNDR3SAxvAkS36
sDRjaeWauuwj9THI005cI/DeEFo6cIQUvS5RatksrfmFgpSClcVzY4cYpDgkFIO3
QikOgMs874xXuDDmcSVB0QiD+2280I0Ip4e5zMa4u7hz/H014X7cimf0a/82Tt5t
3v4WPpoQ9XJuQ7rprTcnstO/qxRlI5PEh0KtZVWzolUgtaJWeSk81OcnB87Gc/Hu
Hx3Sa69vHp3mgX35JErwM7YhB0d+9IXGcVPYAHZJhaEO30xcr2lvVax0iYEGo+DS
g2OPqDrMSpqjIbYGJ9/vVKq83rte9W5BNv46tPM2vEgRJOVLbx0SD7vN44CZH9Yz
3CI18MvhRRQfzVMKR0oE96asLlFzZEDS9TiRtwEkUJJ16iIk2CQsZUNTXNSGe9nI
eXLcGIxN793rsAliu6kjxcE7lt4/p+l/68rOYqHr678u/2R+vbj/HelygaDiZLdm
EMHIQ8NuAg1fXQb2w1ODvvEfss4pN2ayUUVkYKyX9Vgky5z3G0tgNDDBvVglTxm0
PPrixH+GdyCcHj1OfdPR6c2xh40LiMj3Hnj0QEa7E/9L0RWnL6d9MDdmGPseldwA
aTWDEhb9iN7eJIDAnR8vvt8JTlLZEDfFlBCtLt5NbPfg2p8EtAQsTkIejGWvxDx1
I7FCuEREAByM2SSGC8V1mDn6X+DZV78nYQ9dM3ELByY8X8ka+XNeXb4u6et0TNos
6dlpUGABOXae2/2JArwPpBSS9l/C8F8L5y+5EHw+UabGTQr4Iamk9gZTtiWuGJNZ
zMnRfAGq6jPmdfOEPSFdGlQNg0nPNk4iOxqq8YMQn+1ZmrwxKNXpnhD4Oa/IX0oK
ZnshXw9mIl9W7F17KimLwVO2/aQY/pjmWMWLyAMJM82cEjk2m+SyX9ZeBz2dkQqt
6fKJ1uV7teXsEnWKZk7tInCoTjt3TqrwE3GyAkGtv9fUhRzfVBqDd68zjGHR4r1W
fMUkHib8Mg7SfDjfrC/2KSmLcykVTYy1KNFUxIqBfe9/UQmzhQxCPWVJNmwR7Lar
/cBWf8SHhCmEfKKrLzi8r5/cX8E0RE7IrsZPwNO8Mn0R7ipBI4jqd5nX678i0gCH
b2C7OBsdUvTa0kkXdCQVVHVgTmwLeU8dbVWHa/17Msj4RXrpti/TYmCJNDXP1jHJ
ZbvaGPcKADB7we51xm1B1Gl0G7ao8OgTwhCyoIcZIoBaJHJVu9tRER1e7qatISW1
y3GELUOeyYnu4qbI51o4xrf2KfZHeYQExN5XTQsYAhtNVBy7lKok+Oml6NiS3s6y
NJbG9GAFrdBvYxw4jj09mxiZ4ugjDN1jD8H/OEusQV2DC+9DrLtrRyWu0Qwa/zKg
fUBz2jr6AzoZ6CD7rwEhJGfU2DOHieuDVm57JoLG+nmiqHirFllyDkDTXCUnbEyH
8bGPN1nLeilS08IIHMnOvPGavM3nzNCmLZEOuUCqQ5gb1hq5g6544h13CqZRfg2Y
wyi2bAZ/Rc6KzuUPQQg8KBMCFU8Sb4ZzFLEmyLLbrZBzo30IM864IjuxH//ghCsZ
crQNMo8KkwICBU158zMJS1NH1lh1oEETByq109T0Kqv9ZyTvhlReg7wmYC0hd5O8
tOrWhRTcpPUbgZsYpRW/tOgPsolgdQLby+eReOBm0NbXldtGXJhRI3bbI9I9kgth
q1Z3F9YDG3A8aEEh/1VTL65bbd011BHO7C9Z6zYchnSStGhUZeFQgfa2mRFtoBXD
zLisQ2kn3qpEozlwKkig7je6wuhXoSTenp6ITFa8hbNO1oOqQ78UiTPKfvMKKklG
ag9Z+kOU15MwYTlCG5zgJcGKWDXL+ZZ0G1tseA429TW0+t4PYLyI1bK9TWs69y/i
vYbxsO/1bHrCk38/J/uv7nUf/qFGTsopUytG7fwYXpzG+OrIsR0uUAtRe9Gm+AeA
+2sYsn2VZqE2DpgDtlazgWauUzPkjaK/1ijBEGGUJjhejziNEaza8m4GxkLQbqf0
PxklBemhEXdzPiMxfvpOOsaFPA32xLRIn7z8pAN9W2jUu5W6xV5ZxFDphHFc2K/D
Q3nykCM+JoNUfyC8g0KQgwr3ilIEnFoK+mWdsdBxd8PON806oJvg9cl1sRqNC/5S
6S+HFKZPKIEg/GPGwaBvwNSE9VE162J0diY2M4kueFrlWZfMbLC6q816NKRkvxKf
oRWkDYKGVAD9oRE0JvXg6uRHr4EjSKojKC8WQrXiS9EURxgAEk0gdLzKGhsxJqIL
UfPmSHBvnCPfvAnCVxRIbiNOUOo4RhjFYbH5Ckc5OVeMTiQzSPwv0jSoYUeg+Sp1
eRfIud0DdHDKXvUocXcSvCcaBIQ1IPh81lKSsbTnMauLBYkIOgsnC3tniGb2Wb+3
btuHxijfotqUb8jZbGg7RobPNjZhsvKIh0m8MXf6uB7Y4WQI1/HOUrJ9Xe3L6uAM
PX4AliMYXlWzKkPuDWF3Mzdd9rIwomWv+lPizJezUT8qHSYVozOeiL9Q4IpIaHh0
+v5uf8rlU9gJ5VsnJwnUwFEWfD0hyadOyVcidvDQB/Y5fKvs2oSmo29mKle5ddqX
jEAEIwokjs7PcBCOzSSbRVq8BUbW/970eWtKkEiFUZWFDCt4QCNi577Xj/Ra0YoZ
+S0PHtNBr6QXhRXXaayiaEIiTIOUQqTq2yTuG2bgDTE3Miq0PnQwuT0K5DfZMtzb
yB6nvhSvURerOES/5s+2Y30xLDZArAI/2Sz+Ku7QRyZuvhkj5EtFCLK/fBoXpw9O
TF/oyA8WdWbh7HZ2BHV5+iufPeIrE5wiRZwp/KAEiEVxr6FvW8ounTijJJke5lMw
yKbSOYJbK/++bEFYhXKMpjreR0Lmgy63JHLl6PINQUSpi0FIguQJ8OdVuqxCu9ks
XiHF2PQVrFlEM7Iv+lBlQGIgNzRXu4mBqjMxhs104SGbn6IU3C0y/W9kZlw1fT43
s6ijmNKqJlfR/T7grlJ/p6IjU+ykUVPBLkhODxIYLRb5Kj1EZTiB3toueGvy1MIu
dG3pbW6A8HgMq5UbsST6cH+P3UDZc9UgcO2rzan+jf0XxVpcAWSmKWhMXiEmxzVd
K3GbQxvX3SUMZohnmQ2ZIVh1eOTpeKEA6A41VP/1b1Cdv+NzPIWZkBX4+iy84NCO
LG8whjuU2FxNMPRlN4rSoT265GeB03six7+0m4TCxsRy1x5qBwdA9z8AcBuJM1B+
74V1Y0I/yZCT7X0In+RL2tQd+P7gc3h8BerKZxwKgST3N3PSJmJFPhq5O/M4Sdvz
6kssNDRruFEEznRqzjwQhU65KH9wB1S6YnuVTH9JNo7rPuejM/CG6mi8WXT3fCrE
n6LZXvzPTD8yPV8bmRwhuC0dBQeO0rpodEVPznFHKKcXq2kki38BMeYnmDeMxmH7
SFDJD5z00gFg4Xmfbpr9jfEYStr7TGKa9rj4Jz6UGtzXBLLe02j2/5LjaEWXBjSZ
rl9CY2L0ZfzwTk01EfyXrZduXwMQv1G3dYxBrXwqwhXN7Cj+IRYm06TzLS7dYWUA
slA8vPOzS3D6vN4mEuzVH+Dji1ZJEiADbdf4nmfJLLuBIwaQvXYlhZjA8breG9Pp
IeBRJKCxaIpVlRyvpq/Hkbi7Quf1+TkPv8t/w97K6awEbfwT9EH8UnXim49fWih4
rOdPVtnsi6PCvCAT0lRq7OfIw59z1lTXYHHMFi4sumwjiNwd4AwEmFUamXl2Irr5
Dj9I7VESduNJfzrdnNsBLa1cH6b5W2yJE139ZLefrCIghS2x8Tsa6AoGfsu+FwqZ
kg/eTIEJ2dHmQkocclYz6ghmcwuDzj2fea86JSkcfbqx4UvmNehs13jtvSspOPGr
sPYECnlIKDrqJeoIswPuOhVYebw+9WFGDf6nsehZfTiayLnDQMBYFswdgzyTTmYj
FdnlWir4hmlvqR5gC0/YpJCC35VP4GX8FK19CD6v2ZqS/EqbRnjKNmyo03XcAZ3a
RPwiJnCQTVTBKuD+nMebYiCDYBx7qCRbskkVXvQDl4fk62PNWPHS+Q8jV6GMqKPe
RQ7sNxCLswzIcgqXD7VXMhQe1ZVwmUU0+N4M3DcBRtuvFFbItMoQno7JuuLDMdW9
2wjbK6wH04tMwLjPZEKZ651BZMt+81Kp0LN168pq8W25cYZ8hYvKzTfsfijuKQ33
YARixjsqTPYh7CXLX5QvEDTLl8/ANhwuJa40Qd3zXBraN5NBNmh9S6s5qBZ7lmeF
K003lqLUkS2DzYNVtM+m6iSVg3r1+63anEWOl2e8U1qQIFCuxhWxKQlTwgi5o9KI
orayObLB134Puj46ZyBjhdKKCEykcSp0jAiwukvG6qxKKB28Ao6jTOgBc+xoR3Z5
7/xqQYYS6wHuCOjVE/sV93cTre69rY8cvVHoOUsDaNOoj0iau1p4P4G7xnqPEchO
ypGltmO200JwjPxgLdmybj14awEN0VD4JbtD1Lj1UyexKSOcQooGPTntnXfcwUHF
5ZcAwZjrW3vpWuvnRDjlpXtp1KUieqWod+6oXHZU6jAIGLR+0JZ2DGx8Rd1h/FK1
qMNEXql8gxkFpYJSVp8hyeXxD6DMkW6xvy37tKggVUJA+vZmck8xoMpJxRTYM2x/
RVUnu4qNL6FVtIM7+j+dTZu6sxxGBnZ4+Pnis4yx+4hX0uEysUSychr6smKTin44
jMVxJQ8oVX1oNw6oPejjswoAewyG9t9gtTlRQqPx6aTwGwJw+DLYUv3EeYz/06DP
3DqI0Sm342gtZItp4NS/qpPRh0aVFA0iAuruVR0YxpMdI1dV4Ios1ATBqHZ3KY0O
2f0nivmdqnr6YMdKZ5pULMyRx1Dyiw83Qi9fIz10U3UXzc6paIgkI3jlJG6OzbcZ
xBLkiPC6SDJ0t8ApnA0srIUBJV7O0U+yXk37HpMB3icIk5n8XyS1tcADulLUOXKy
kv6jtbxUq/w8OMNQjbDidZKxs+XDgGHz/Ms3rQqQop1N18/u5UbK1v1PWTMMutp0
FU+Mp8zPcy862jUyr31ohtPBaA+YHCM+cc4/EHsO1A4Slx83YRx5bfuESK3dbtMj
/3qhxysEXyegZ8fZ7O6fv0j+j/4WSr8guOjEtRHzpfs00r/H4wdPqk8O3vMvwDgm
eQRD4/LeMswHmU2U9orNrdls2FiP736GdH+hD+SeAA7gqqS9gZ0CkKLzDqz81bMz
D8chpDUUifIrSRZk//u8FVo5YzC/iPtI8Bzt6BoavpBswhQPxTqGMLJmh5kuASRU
Rd21bKKWHW6XbuDWXP8e0Zlpyrh3ajgCXz5s+J1LtclVCm+9mc0ErgzXzgfj4tCK
sIC/8ixm3CfHIzxoAWt4BthTrWDvLtF6k53pcvwcfIu133IXJsh7WXIQgzFeRzMe
7IYLVpMIHL46T5i1qKex0ZSUkKc8IhL0hZ8stvM9NqEuhXvF4qrKpEsUpM6uqpdU
wrDOxfSYglMjei7eVNVOKsxeQN9GV7Xcf3UI7VYo/156fkwaUcsYCrK9sccFAKd9
ZGizYgTEyELX85lb0noeAKIR3LW+OrBpEUe/oWkgzSsOu/oiQO98xI/ZS36ikGlQ
VCpyof6CC9zqSislB2zcfDjEFcQSznXjr2fCjGpVmUYmd65BnLUNOEMgp7tzKrid
2lmTE0TslD2jDqB8PVXN+Wdt8M2xZa7/o+/BoQ5YD/hZVsrx2bS8KylE+NOBd5sp
gzpqsMZ0oLbjr3AavGNnO94+CJAVMtluy3WucGcaxBdXfs1VgTvq3b0LxN+SyVlM
yOOkXqgmPj/SdBvbYZxeTmapxU6coWhr3C4He8Dm2cagc/M2bpvZWCXlch070mvb
K42p4g9fjy55x1rBbUYZSOYp3opjvjTLGD9MtEZbBX45UT4B4+HSbtj6lSKO5mXJ
1wqYlBPoOgiPyVgwBM5U14vFNuIiwZ/PDaha8choqb9S+AVJuWF8tWDALhLcvixc
eTbBz2LPaoKK3ghRMk+Dqn05SbxBOl1wgHFzUD7CtQBlikR+JxgXLM2P7CRGIY+c
kPxIlya4bytyNeisJMlTKx2v3t0Vy+ajL5skx2/OxCvgVKqo7a9aBYAY7gniv7W7
4rzLVghl6bgB/D1Novc5LwojTdL1jfDpj+2dFrKOiRGYuP5r+1id107TTVrVyhCJ
zRNkCHVJG5XlwdorpJZUwOCWHJHMAw1AJRR8nTWgRWdEmdgj0cl9Oc3HetR6cww+
Ru2Wwn6gntiQlorkmvaovVaZUNviUrx0K7G5Ka77a8uaokZXRqoPbhTpHT4IEF2N
lT4ixF67thezzfppOMXcwH/gJ8h/gieIfpbZrQ2NH32mU5fn5njNq0Y7Bkwu+dGE
vtdDlWq+cr9ozk/xSTJyRhCc7UzC5NmoMpyR4j1nc/pNC7thiHvRHT3pe6FNhK+0
WWSArQEk4Q9mgeiI8cPJXj80upKtFyJ9u1KTnrT25FKFUwU9wu/sXfB9qoyTCLU8
jEGsA4cm8nclbBk88n3bvYy1wrk/JFwO6vi+k/u1halhq5JfT8ECAIVZ/8+m7V6C
OLgjN/EZl993Nl+DcCYTA1XWTfLR0MvfXIWl0k9hUOm2ufjqfjYSSVVzlxVADkcV
sz53RQHmkQAy9oxNT4I3u3k+07mKK40ct1C8gcKe4gWxg3MtBeNKlcthh1Uel9Ze
A9CWPP2e0TsEE8FiFZavk74bsq5+w4vgwC6GP/QUsrv0zYImfYszBE64ha2wcB6c
hKPDmbLjPAcMccszPX7H3i2fWDHosAgSO1btjbsXKuC35o2cxsxtZZG8x9kC18hA
mIYVgN0CXHK7alHT4iUM51GRlj5MUBmGNXNpsTkxw+X1l1d6YVTxlJUlGJfqmNef
cIUXfrbGUt8ky324bmlZZDEZ/XIBMQR2lzuZr4jz0Or9JlJTQ8a/U36LI17a5QNN
Dj4WTYbpjFBGbXJEsC+m6e9edVc9Qpse2oo+tkwo9F6KoOWf9fuvd+VkvsuFalzW
ZYWXCWyikWOtM11WxiUeQ0AnHKtO3S6KyN1ZImfn+OD8CSBtH8XL7KdPCO/ZmcsI
ZGJkLmBeSqGIEe1pZ0gXgwFkQkOrqEJMGCPz+lUJ1WKWCbQfJN1lGkTJ/X4++U8x
zBBwZA69bPTOT2EF/zKAQV3TW7vNucXQj3WDChZFlZRpm6Ql4TaKnH6+2asSDkoJ
FELZHfcAFPzpMEGT0jdr7bh/jM7D8w9WpG0JUFvO1rtpqB+vF1CIBisaqIJ+jEcw
/B8Uy+iu4RQcgNN7K6K+R3bbxlOcZwQr7iaveB0Nve0198+AJLeC1LVyTPCOx+vT
wx2EYXHIJzGutIvZ38YPoVQfVRISjfdWZi4zYuFug0pwIY7ivPJNAWHMiwEUMk38
rXDT/XSyAf5Q+mbZ+UEio9l1OTwHKQlO/BUx7eu76/srVAjC1mEyuWLmIJdzYn+P
+enrs5Kql6BXOznKp6pAC5SlxVcWkQlMR0XGyh6t8d8nKf6sgHvQsyaGycroY1aD
sg2u2EHI7UOc1HtYhNEJZUXSKfvXKp15Y4uLV4FOQnLakgMM2uKzXQ82eZz8BeAJ
exXDaAQQMptyEQJ1xbB7qyLoMwqekCk/bTXTpjskb4bQOtxzQSlG2LRXT+M1ehKZ
UE2PSbEYOSAYxZcV1PKlqeJqcmqMVFaQwGhm3BtFnDEQ23kQQKOzv7JYdJgBgWSH
6r0blRTQw5bmJcGLtJ5ks/ggX1FInDgkgzmPgdME8kQCApMl8aos4ki6wADZD4HN
08fK9WwG3Ywn9/ZQF9bakEqDoK3cvMJiuARsnfi46LRGwnG2vUnlzZ1F6bKDAVMa
QQByqckspGn1D/7OQNndRlOh79M+i1+iYKzeQuqUXS09wnaQXUo0Hdu03grn9sZy
aj10FlEcGUK0Cxd9mjgivON1H9iY1E9LTOwTQ8DFtuEQxbNfxKI2LCMWlMuG7/Be
ZbzSt90aTu9Jjq+X+GqwtEtjCwJ5ppsJgLNkdsm3EgMnR0b/XnV+YCOnZa48TmZg
V9x/3BHuYXBHEugL7CH+/Kc9yiVhzC1zB9OxPCkdgPYp5YKCmRY4qZRwInbeBgn4
AUm7lkK3wI8ZP3yyqRPxO5YTbrIXt/bkdMwbkb8+Wk0Q3eo2xkqSclnwevNfDDF7
cxMdjIXU79g+rCGF3fmd92lSZ4TqxLVHOsM5/rutj3qPb3oWplbcbB+yebOPLpIK
4HVGAC1suQ53SOBI7/kdPH3xjtpE7xVi6D4CqUGIqEDdVodSPgUGiJCVNJYnzFnu
yf5co5j+L7pId2DYIm6E0BEQJD7zrZ94aeyo8GkAMGEpJgoIlMDEa2sYUVG/m2Wv
5+IkMFLXQNfy19/piVeDh42cG1dQeLMOTi13ljF8euS8aVSAl9jQsG6aRpGyqVsm
FATnh7kG4eX/9xqjC6cQwa58l+hUL/FR7mquJ2IEOsGt6HDf9mx9fdgjdca9Cbps
GzgEKDgWJlPdzAr3YGoVID6KWli8YtTLllWi9sow7mxiC4S268BjrS2nZYk3QpJK
K04qrFWMqBOlhdJpy7/IX0FSx7LpWetT0qiw+cp522aqrCuNvGgx2LyRhOBMxhXZ
GYaCCyf0XDX33Y5+d4FgkzyzNXiNg7uA96qeiZ+LKlogbB9vHWpcjCe/vojghwJR
AHgeyFLWr/i1W9jgDnSOk3nPbVCpypV391icMxiFU4Jq49AlxASAXInX7ux8tRGv
pYHLtm/6MXFMbQ6s0wwq8K1hpN7UwKqPKeDikYytTY2aHEjUYZVVHelftMhhH6b7
DDe6G8ayl9YRDrtUQFecnttP9xIRSYtrKS/atVcDTK8Hxz/mbQ7eKHadXNSo85Ot
9vKv/w1O1yGt8MEP8k1sDuGiFKYdXZRxXnsDPJ+DMCWeKXkFlzKXb6NUrsGm0JVe
HQXwcpMc5Rm7zqiF2W9lZomhJqHNi4r1IHmiF3Lb45j45leR3+Cn6Jz920k4aFPR
5b69wixv3KZTuRmLtZxtG3Kfd/P3kYoqNmaRww4nhxVEK7OdXQAY5OePfpGRXRoC
BIWR25lv/bPivxVFhLSKj1J/wqjPqLn7PjiMIJomrHTLkRYi5JRr163hwbTWjPPy
9RE8cHXtW0s+UmuILvaLoJ8mdNYsr6Cyu2dZHkppujAcantOek6EfG0kR52QiWiN
CPZj8LVvPsUN7Q2qtjdpQZy0tPlIFsvqGph6I8B/53I6hDrGc+jzJ2abgva+fqrk
fpQgh5EgnRWNNgff7OrKLOOLNWN2Y78FNLUe6tUr1qisJAs/ruHbZ7sRxwavoxj6
aZ5eMTkRP87THNnvQMwk0XpGE/v2g2E3Kj+Fm8h5DIlmMm7eQ3V2ydpiWOUmjJQl
GaUPwkyuMKCil0Kdhiwd87M/U0xJv3JB+E4GhdcsjtRVWCFg/C5TJvf3rLpyh/L0
+eDZxivWYe1i8qL6lJAjUgkOr0EL+YlG85/ILTyw+V4VAdV9w9+cvUq3kDCC+dME
aFbum2qsiz78wb7MvOAa3GL6Kuy4aTyvWeIWwrsyllqbt3L26kxh4jSgkqV39QwG
fOfOaTuwcnnPkYus7JN5+UxIwZ8zuLX6rXNxG1DeZ9Q9Hqs+OdKeFUtMRFjiDO7l
Wxk4c2+ToSaL+4V9MWQ6nuyo2SeFNj6cBIfpUNpZ+KOS2xypJ5p4XGy+qQBlpmGA
pZia8y6ts/obBZC1Rit8ecUVjM7lWLYfPTTx7Dw7H0PcpYXyck8pCMR+rA2BPwuK
UlF0nGQ8xf4xwJRD513IkoQopOCdkjAAJcaGv7fZPhjYs3r1yUsRa5nSQFSbyHYg
IYSuyRF3XM3HtaUwlrgIRr7ODQDdcXKPMW1a0/D2TmYd+3dVOtK+8hgDXHzDmu0W
tJZAY4+9R/ER7ZMvp+sNm7IllG0xbZmEpBN+CTzoWoVOIyo/tdcf5PFTcL/4DW24
34qVPUNjta2qDG4+u9wcYRAYSV85PUbJhZXcVWfN9fbtvFtA06zVumzwRoje+ify
HCV4XVn8/PI/Ze4hCVGppiYBP3mDQ/87SxMk02QSZV/uaAD1jBC+1OeW/Qk3PFpG
ScEX4WN4Kd2uo4TDcxjhEcksFuIBmLOdoQ58IfAyieLhE994phggy1xptXQxaLlj
MW9Zw6P/x9L1VQeEwByy971yNvmpldBAaUnqiUiWu2uSgmJX0mkWVmAr3swpNnk4
eJRjLOvjmNkuigyCAQ/DCh6NI4o7ATSmKf3SrloX/nweJj0hQ5EgRJGuDux1FI/T
OXfgZ7EQ24tEjlMVIXm9vWy2j2N6/93EFBe82EH6R+0oR+/K/A6bBoTMjIApGe0k
MRO387wrcaHbJ+yde+10xTYLY4CWCOHNPBouB3vLzZUoBIKN/8CCPDl0v4+R9Twj
S0BaniRtdDPFaZdnNp4c8tyiyT5pNiOfNBYWe2Ao2xI2PjFCrtpgeqe46G9rG3CG
IKYiKTwIxQVjeoeJ907n/sD8GRYffikmOspT5yor9zi0FiUCBbjMmnKm3XYvVNlO
+++GX7dc221Y6lJUzgbj13dlunYCwNSz2mF1z0qBhSZ1O8lG2LFwhtb1LWrsuynT
nfAz1085eVPz36s7g24xHC+F0+eDBLn+ZgLXpYbsqtd2e37e/HIYDFa/q9AHuF3t
+UzpiO4AFWltCZBlP/F5DOrHh8AyKTRAvz73MuB9aWGXwYXXsX8tpNY83w5uNzgW
a5uxKuv+Semma/haZShLc38hVZhox53KZC5fgwBtKjsPuA9yjYOFDnLx1+oZG7a5
oWfD/HoX7taZyqH5uB3y8x/ML7fECqjo7yWofjakmpmofvZRyZpj7McrhHAZRAKI
kZhkrzCIBQFPsTp/H3AVUEpNjgIS40Ww6CWmYhcF6qlBVI47wtI5IreosI67z8S1
GunnIDuZ02OLfbITE3LFJj6GQ7zaMuaNSoTwPgm1w0MXsGBEuoWF/Ed+FPGLG2qy
m7FL+C1fNpxaQpyGsbHnecv/5wYDv8zgd2nfYdnpXzsAobctAtjGurj2AjM/V06N
96EWGBR7MaAbSJtpmvKq0H1v9pnyqXuwfzer2gF5RAzODJGapv7t+b7OfwkDvfy0
OfbbMfC93EBSbhXEFUw+wzQLgUAWzK5TVLM3NMqSa/TEHFWHWFr01OtTy85KdlXm
qcTGbKvutQXOl755vZJcdxYmO//qm+to7Xbyt9BX+MCiJxgoSXEnenb0rshRj/tN
bx5T9GKZI1Jorj4oK+FbLrwkSB4o+f5a4ks918U0LTnJtZNCE/GRzfzv+8WJ4Ouj
1aKrZ1Avu+xUKgGc4/VYs7UcTfg7qQYLXfEmtpMe9V/uLAF2NS7Wgx2Q5lYE19jR
ydUt4XYhnoFkPAXQnM2VSQ0p+Dv7PsPCQn5v8Infx6BnJuOzFPDnZumQgXTER8MN
+dCyOSfCX69u8eO43OAx9xW07G5A04ajvHhvcZpXzk6CSsILn0JAk9xImnoGzgM5
8hauitkx/sQ8nF1NW0zYcGOhtH/Av81Gb+JyMk9M8M+8zOG9/jdxWxnqDrwCSUqB
nukdEBhDfZB9IancClniUuXAj/G5en45WjlwfBg59yCq7GBWRUWVJahwN7Yni3DU
7gVYQOz4+dPsXVg7S4gajYMIIn8HUu+/14M3oivxmGkru1L0MNd/PSDXUer/rvLU
lVzYTV7VBurmG3+Cex+hD4LILwNN2YgXgRRb2RAfWBJ3jk61CtgZV6PeTFBYv730
z8HRJEacUx6MCDd7whe493Hws4T9ZGJZ2rQCEZxyFT0awzVW2h3nxczhNraeA0oj
U3QyOBApXa12hhj6INtFC8YanwJkFEt/7KsfP+LP+OturLDefxdC8DcN1yPFE5JW
DbtQzszlJ+Y0dliYxAWlMw3U5x5YdT1R6jNIIEe8PZtysvEdAXWSXohyOBo3flKH
TdlIODn4Ox9+LUiRtkaSeLC4iXM4eIvZui9PPS8n0TWWxo/xdO839Wry8MjmBVp2
3vLOjdM4TuCnQkS+iFs3a6pA6b8uAfluW5VwFY1NlPA7U9UXLbd5swgoXsUCTabX
vY/R51MNNV+XLw6UAr4H8yRRhD74Aou6dyj0CK+eAFk2h7CXRGGvoW9wCyRT1+tj
+mcPsG3jOgBGelTdOx1FD3ayoU6anCHbby7R+G8zdJoyLtz+uHDoE5wF3i+hwIue
qe3wQKULgb0dCP7cOTPouSqFISYWDCxCrq0HVeMMlfAH83hsczpYMhiMiWG3bHdh
xJFz5qRWe8l/Dg5QBdzfgXbEcShdVXkOIWI0HIO+7nLHnI+wzAWc2x1OCgLwwZGr
MrxzVbW8DTzmbS1HlNkSBhtUVamj2zoCKsJEmJNr0OhgLI523lHPpmoobFXhywe8
hqlHwzQLk1XaFuF4wTzSIYssBnpy7orWqE+tbIYy1m3rc6/FJWy+IBoqi8xSPe+8
XnAgJQRE+yfsho+JiG6ecTjXoV0aienTKqLHq1+vkSBRvAYyZZCumqoOoPxO3Vvz
nmoNzf4FETvKqBio0VjMfixLfmF0HZzE7+eaqmbuMYt4sBWTbLaNrggMBgqRBDKs
BW84PH3Ta0pJc6HeypCnmNATX+aptv8P7CA3/uNPsxsP0SgZzSttPjrEqUSGKvVO
T/hKIggCemdyueRy8XrKcIlc0bPQ0AcZePmvrVmz7uam2cvLVayWcegL4EEHzys8
/ewrwn8v2Ab2PSzWdItxUWqeU7797z9kjNjl3tER7lqKSzgNupfN4BnZGZ2VMXOT
A0VpgUCGS31xnpZG9foNf8P6/F1r7oCxNtZrFCNHAan7EaZZWfbhbjo47+UNrxcJ
dXCpdf7sz7K237CAWuC+CwVIe0qTUIDPkDnIHx7PObKPP0OI6dVjinMNHRrVbR45
1DLmOUmsr4RuUKhrgOpTI0ff2RxAF/TAwk+pripGDOPSHoVIkb3Ke8HRwwhfFoB9
NgFQre6mCB+NJ3ue0DpVIcdkb8DiK9b92qsc+htrntK86E1JZSU6JzLjByWT5wfg
59ni3SOnN4AJl/1wvwGJYACC8kGArD+hXq4mI5PE3PA8KmOlteeit5nSPkvu/UHj
hkSOFMc98BI9UC6DuTzXTk+ksslvZ3Va9/QtaJWMSQoYGJRHKFKW3Y8rvfFFzJ5D
bU8RYrHkfzeGkE6lbqgsESbxb2KUGgWK98gy+q8WLI1PjaNFhQmzHBujOn54QbQb
ALQVoHbn/4/3nJs/8t6SqyIfXMHTEb38Wsy29YFJGDl1uvE0OtFtCDspR1mfe2OI
JBNk7Ir96ztZzRcuJuLHE3Nf9BuKDJ340MrsBRjbjBxZ1asQYa+oAUOcjYpE6Ovf
e7/Hgj12SZs5wId6jBZB89EmHPmX/KiLqP/EbyoM2G3E61jVhfgX1XCrqvImUwlO
2PFjktWmawYa25O6XTpybcuhRgT1YMV7LVFGMu4PLCELj34UAGKCRMGM73PHJ3XF
qIWjWfzaOx95aNLeu9TYNMY9J/oroOuwQBcBRd7NyT7VXzqRL47VZAt16xTsZYZy
F88+6OeDjt7DJ/kJl0rqdT5Efyqujg2l8kL/bjBdneieGOekHLU99sY2/P4+GnRS
nij+P6za0qrls1LCrd8k8sS6Q8Xvms/itribgsLAZNimLOpuRiZSQYbj0RTd47Nv
aeO+hu9x15iP9Hi5tSOXxdTw5Sf/oot+geMqbfPQKqEWhym/OKEdoTax5elLueu2
Xs45Y/xWoeaElvht42FOfudjM1jgVIhuc7lQUkU6y7h1qVBjqC6bSci7Bt+5kYmr
ANP72ebAEP1PguGxjFY0wIPWMjmmTCWMwwq3Z2ErzDcuqeYiMhFUbyT+zbEyb9rm
L66iuzO9+ajfYwLECZ1hIiVVek78RO1dlrRycXw3a2BEDfqC5tZQIfw/VYvZaJDY
6+K9d7s7YQsFKnLzAmH7ia6DDRjWvti6Pz4AP0I39Rrx5jF4TaECeaXMZjjOKN8c
PZJAm6eqnLz4XQhpNXiO5TwujezPIFQzZ58/q/IGTJNlw5Z4jGun/q2W4gQCs3Iv
YTQ/ErcfqdmQm3oaMBWgYqYGGphWxWz16EG3hCaAMmWvPnr6ONCx48iOPsEgmKYi
oF1vlIR82mOgfWFG2Gn712tkqe1pKFPLeGhZmB8eNxEfa1oHkL949ETj4pTPuNSI
fl5JKiLMUqvVd6qFXXF+jwuUbC36xfBd4bENFciuBgTsNUmD29FM0NK1YEG/KA1h
a6slXpUT2c7/Wy3j/DhCGmq7zPFjflAfqltdJIVIFcDLHMwWaIF8uOTAo2v3zQnM
5yNZrnH9DUSK+raA5qgxZbdcEXsFH+TOD4Efsa7eqvZt4yG9Li2wyyK+sxczQ2Ls
YV6eAS91+DChOW0CbRLhj49aj6zsJBcc0xbyMWdf48UjkfCaxsryf5IbVCnhF7PU
qJZ5Uxj/Vi67vey9JshuaR46aYIkhJrPkC3OV2mJ8/yPaUahwSugjHOZtAbJMu4Y
h1u8p6KhVGVklICEJEjKRDVLjtHuDE/XK/UN3WzsKyXt0GZGZkIBwPCjs1ZTdKLD
H1rUvvQaFJ5G9v0ykbtfMfZQQTkOZP8DGywxkqOYxzYR46hXnnkO5nPhaNQq+oiD
/xdfpl/dlm0qgcuu8iguxybv5xNG0iZDzT2fhLo0K38QozsjiLr3ejKkysGM95ol
+Yj2osHnk37g3WRuglBq+czVlV0ieMNIhmPP0XMxyDCRpLgFuY/BH/L36edwDf1C
opkW0MiRojim8PfGryCfW4XQ61W6n18OTiFfCxdhr04U0In91FnDP7S9A2qS8Udu
UAuLZwrtHx1xYp50N2HwOazT5US4sCnq5Gr3fgU5z3jJ6VxTKsz1BOI6/PnNreSb
IxbHFeNJNQTpl9gZQu09Zp12NFL06u0br+9olfSMB/VWk+FiGrULtY2Z0HXNz8MP
SE22UdlnODTfeB27GKVfkUEW8dxIF7I4Iuc4l5XrYo67Fe7SeHkCgdzxTYi+Rq3x
cORnY9DKfSn4ktHGeNWjzvsbaFhee9xr1hp2Rk4AQ9S1tKMqCkcbj0s7ao4jp6Ct
F/QLsjU1Qpg44YgF7qnVZq+yEQhNtpk3zXeeOgoonWFZp/IoFX9k7kXjmjwzIRqH
o7hIEvdq9savo/kFXHoJ7JzjOs64FKOMOw+/M8XRy+U4B+QS7RG2UnV+trhzt16c
oqObEcpbdhaqOS/gEU8RJ2ve5TnoahcmUc9c4Di5H6rtpHHHK73aAfXoupjZl10P
9HM8gQ58GiHmsFtnVwihAkjeZZjfWPXSM7j2hyFrc2tF8l3YBEQKqQVUkC5+RVpc
p8syx/RY+P+ag9Yn852pH4MNwspH2wnV49ql1y0hSHQKGg8Qu1+3aj1zdRm5/QCG
sm1Xgzixm64zNC1u9LcKJin7uFZY2iXiXCKhjhAvcWGr3txc8B4Cm6bgRS3YEDBR
qyJE1k7kjf1+2JE5lhEBC8bmDa/gHadBK3OBooK4mAQUSxiv8ExwQoquVt/ZXdcr
z/XLNsY+2Sel6rNDAyDVhhQjXewjlKM89gJ9Deyl+sYF6Bnwkc7iZNn44YicFupU
4ptTCF1m4qbx89YKIz8mhdsXmN5kr7Ej+akDHEKbXA0WZJUEcmfLjo5epl5Z8zn6
mEhbnWniYABFRjHiQ512obpPiqWW+NbR/RGL0MacutAFZJsWYJk+pUtRrlNNJauH
wHxYSGpS//Huj4doRiq1WNTI8yLpKYiEp98K17ea3eUJwC+gpK65WOoJkYqFXGXl
0WLLsHBcjamY1rFADRDwqIlOEaV7Wq2lTOjXjMidKYexgvGaThJx/Fdu+gsEwKjQ
5KzOrrH3o3hZ366q9CgrvJfULUq48D6WQ8ELFZF8WAGABNWzNOlp+PIYfHCY3O1J
29sooQxcC4GvVCyIWvsomh757CwDi9xgam8jOiSj7N+ChTVDT0ZuvxZ21FSPKzW3
kx2OBFn8bjFyEhjiNlyohsdgdjAMsjoZfB0kf8plzERzc9l0yfUr8O9Os+l/xbEH
bWDaRl0NVxBhfrqBysFZrb+MI08Oo3KUh3I5GGi0dN1tPE/Bcgu4JVV843e7PHk6
U+ee6CLoRt48qt/BQNAGkgQ5yoEK/ZOM9QDmvlmzREA9Tb9g8mopt5iCpYaxj86E
Ma+k/zOgdE1M3cE2pcM507ue15yOkUCJKTtjF3oYbbcdGICC5susRZlJN9XZSywZ
1bhbE7o8dBgbVcjMWDa6IbDso8v3KpVvfY+X3bVNqwW7MLZWqXZWUEEVWSiEhePn
e/4u0jq8gBJuYcQrX14nmbMAP45v1RE1SBNEn28pvkH9iLWK0C9CX5ZLN5hRWAHP
ZXPJnBQiziwElodxGneAFW05qK2eJkZNYT4/Qispp8sLEGgr1u7L9bW2n6wc0Pd0
x1RZEKXxlKUvrb2snBNn+qXVIrgMdYlMRHFg3AuNDlnp171k9W0CDkL7oZFaSc4r
g2EBvdhWoa0LbKK+zKZQvblfq3uJxEsinXwzoBD2pLBbCp5OPt3wgC7tHOADvrj1
XfzFmG4FKh32XSK7h1NtbFGv2GTdOjHi1LP4XRHygbiLlo+lj0I6PXmY3ckEo3YY
H49d4mmXKRDpAYfyxRdPdT2Sew23xD/nHAdgnkFjNUxKbzpkpJPRRBha/8Pa24sR
io8MiVz/W9EN8X5lwU8tE4euks2tCw33vdC5sLDXfopF0W+k4OkvIjAbTm4emxzw
MJUEVphCPv+Xmwr6etKICu74o7t+b9g7bW9qom2ZXi6boHsSA53Op908MEen5DsS
W+/2quxePK85LXIrtuXLwZ9wTiQE787CVGBx9rIW1sJ4/n1gRLiH1MlrFJfhFUmZ
r3EzzGBfoiuqIVOsG/NaJlhWPr1SAQdf/WD3S8kqngIE40FVTa8bSXmdm8U80W2J
yy4BQ7bm/1BNXbcQnKi+e9VXnm32woofOGhnSkDlrRgdBR3Upu+2ae+s0tFxG0E3
x6xy7AyX07bJknvAydQ4F592pJZl6H9vsKbYjn3uqK0K8MOiJ3R1bhB0pjWX+W4R
qAuM4+iKAA1asxiHfaNu9IOwzoKWQ7xeB6bW+QZ79BLIfg5AD3/2MWVQHunSmj5r
nLa5l4yam+mSuGdPJUf+twCop0nVvecBCFNw3mo/QlH/BK+OFThCVg8Npy5/E0a+
5hEjRolXRkC0JKSM+2T8MpRqTj13ElUJxsWtW9EhSM5LSkT0xTYrqGgUM9+9QtW+
PqrXuNv3ViKrbYpHIgH2haV+HRa484fH3tKwDEvuStIMNX5IMfm4zL0I+be970yG
eU3Sk6yvxSSsqEE5Q++dPE/dB1doaQKPq/+u6cSY/0K8k1MtFiJxJ02nwEonePac
urwRF7i7U4y0M/IzXFGjPT3AUYXlY9Ic2M3tNVEvmpKAw2VYm9WCXvAuazTMsoT8
AHyeCjXyX+Bs3c0eV2BpGgk6yk5eySSp2e17NiiLcQ5IvJ1EmE1s8cKeaq+1vdeJ
9VbA/pH3nTp/rybGkRIZYgZGZ78LRYjA+Lwu3QcVoWGtoOXI4jVErAClaEAGip1E
n+fKl3C2x60tPMz+CSjCR0FuRnkpG55F/WrVi/WLtd8TuWw/y/Po12kaoCsvc9Gf
EByGYfzUZ3nHES6VNZhvZTDi8K9wbTVIgarySf3JS+Vs1345IYEcVDSsrFn24EkS
2cGkSBSjgP3OGsOJNe69KuQFTPzFGbZ/snUIinpK2IXXnevqEo+wJXPTXnGp0u21
dWIcLI3UoxohTesgxowYCp/+11bvcRXIL30NBBCuhJ26cDrWCqPZWLor0gM25HKh
jB8S5kUaS/Fzap32v0Hrd6qNRfNFgKI9GKFtAlPUwVaDByeSfHc4yG6TOZHZX6SY
0fq74PfBWKkL5NrBSGTpOJK4PVnZdDuF4pUUzVnO3sjKQ1FZgV7+wlmIRaIV/b01
3zp80bicBJMS69Z5JjLnCPqsthRz0jcdSV5LBM1GvupzUW90cCBnYbu5/cLriO6M
9cqWsZ+VfS8kesDgzfanQwQveEV6ro8zGNAIKlyo5rq6bvBLRpPtALy5fX4v5ocX
AN0gxMJfeZKPk8QqfMPc7k7h+bQG1dH49xst9fQ0tnSWlFXzQNater6OTZluMxLy
qxsvj63UnpcOZ4BDcN9FA/8Fq5s/9gjZA8e/tcWamaTQkF6/c7dKBHNjeNwFp/iT
1lZViRewRSOyY/T1pkjmw5oP7WSz8Xr1s7beYbZx2phIaImx3puvtEEH7/tYloMR
J4kc+O2AvyytCXt2xcAbcbMOFNpRQNr04zZoelJhojVgHA1NiAnhbXbIUg+7m0ap
bqiWQ7vsU4RTIhC48+WzLvpMjuLAgxE8jXtvx6wF/dxqNkUqKF9/MOS/Tjnson1s
6d7ve8++dUTNsfC5jj4fFqEWyoiWvzWoFy9uDGIB8B/8IcIswy/LEKZ6EptP9hbe
z58Ux1CHvQ9Zl+w2sM/hJ7BQ2Nk4irCWq3ZwCrwUteFUyQHHm749grLoHfbiSXqF
dCTUj5EQn5FKPZ01pkREuvOjw2igp2wA40joazWZENRj63xFvx45xKWhG0BTuyvq
ZFp/NDxCIxsOiMo1k1/t9mdUayOeByOePDiyzVse/Ao4SKfg123PYtgOKZFFliGr
vZBL6NVDpzkVC7g0M3/9Pw1mQ2LXpihZBfDHU7SxCiEYOov7RXDaN3JkWAOW8rlE
bGj3rr7mnljo8D2AySRQ2+n6mY2iif8UPmotd5B3fcCC4tpRtyaFcgzVIfLGyrPf
Incmaa8Lany9nDIDD174HTtqXbyE0Hh0FUzsut7hA6dWnqDY7pUY7b1ZMG+9otL/
Ri4EZtTrlr5kbOZX04Qn7LCCmfVMB4QyAZtZaCh2KJbjYLGjq1sUL2Pi7LohoLmg
dRzf2n6oBOzdEM9c+5R+4NB0TmTOy1hiRYg6qQHz/RzVHitmmRUB3821AwVE8Ydj
iGFeya056b0Ai6Afb4uiCz/RpfL80U2xrL2/iNRpQgDj8n6B3ARBO/HhEQzGOGL3
S+MR9o/2eF9OtTjbGyOQGtEyP99rsMrQKsMNdwtQ6md1TUHdNLVH+hrFlkUOHCPe
S1FofUzTWIJs5r4WxoMDG9Rpg7o95tOOEJyIY82OnUHiR/Bohh1G82I6mDKPJGZN
pLibBmWGDpgjezyFB6Fx/c1UtDMSCoUc8LjK8HM+ufufgBMXyfqHfm5cvfw+onNc
uH/fKWyWg88mALSwyEHMhu26VhEz9rMFqaXVp8FlJZIRM8Qs4d22f02DYEJ/t9vf
z8iJtHkA/8R36ydgqiT3508r7/3v9I8slsaC6FnpUvBf6cWwWhMtqzhxeylf/v7T
wkpdscLcSuDP/xUbdWyoJ2xSd4Wfjks/vU8/Jbwgy6l9u2dmZCneLYlMsD2b9JeY
pglunN4AR4tHi+2IUs+YTW6YZdNCUV26JkFeUFcgYPVjRLeRO/SpXgk1RiZi+L30
ls1OM3v2DgNglkPUDNEjd8p4YcHqj8gjblt/umZLO42Zv9eMtYdQTr3WDSDxjtKx
9+8Fs1KOm3o7uefSfIF0I9inPwH76kiDRj1Pk1H0Ae7HpJuPZceLLb4lTVxvGBMp
mS81wWlcPJ9MR4kYoCXn1ja1I/869jvEVegsv7t9dySOwxMdaAkp1NjnLd5RPDSY
C0hC+mZYflUgmh4tOAI+QIAMQGIs8Z06aWc9Y7KUQ4e9ZgmWchvCtR5SK+C6BIaD
PJMB2GLQsX6Ih7x2yhPh55xqzW1U+Q4tu2X9J5m1U/kpp0vZtC7DGqrCZxGaYaK8
c+p59dhGbA4/NZt3wjXJqmUb8bIimACjCfHnTeLDO4P6GOHcmcJOnRQzToh5L1Zh
m5wI2J93/Dqb0V1CrKgmvaAg6N2CvR6APYQzpcqr1PZ1BJ/siimd24jPMXLVvYRL
yaw4Z2Nyjrl3SeuPNaK2bf4sm+IEGDy+T9yBk/u5dTj3QifD707OXwKAFTXLeJ4W
FhBxPGNWRW8RZNY4sy9fIEkUNTtN2td0jgFQA/T1yJ9HDh2tHiiY4l+37a0yALhQ
3ubO4nMEJnyPVtheizlFySFoYe2qobbDDZI3zMLtnGmau/ZCcJ3I6+am9A6LoFkn
2Bi3Bvtx52d+ASm+ZmKSNHLUD8Ps5OVauh1bkoQ/fLZ1gIoP1sB2fDrzeqW976Ux
UA1tEm+O6SGWFciw+PtH8KMNVpHfvHSnoywKO9dSvXiuws4Tby/rqHBTjh5Glx08
5DTLivWkcc5WJRObh+U6m8/uE5rHZ8cKow7OSE+yQdZbTVUEsm2b3a55AZ1YULce
sBBW/mwDpjaA3EMKqn8xP/7sRnqDnZ3lhJOgwjOMzBgN/cDDcw1GDC4AfnBMy4Wi
Uw+HfykyVEBUDJO72bO/288w4Ty1Su/XbIy+fb8rl7u2+YbPIi1kBpn80PoSHpD1
bS6XAc+/hFITpocXz3X14MRQY7J2rk6i/sDub+qhOBUYLooncAPOMDFyJ+QKPVxr
pUY8haLV7UdAmZoZfAqeHB+CfJUozSHwK7V41VzR3eXhs/lARuoQFuK1g4ec8cTj
Ju90MjAwxugdDSsFeI9kDw9o8EpdzKMUafLKi4a9iTVXSkhkJLpP6p4sg63vA2n6
j+eQcHiAnBfG5KqjF2chB21Cam6ltc8t5HfZeQCgdhz8/NV2GwCx5JE+W396P7nB
YUBgp+IS19nlE43AXf/6LkQbGiIphO81HC4Jm3tVNifVoC6WDZlZ0hYUWJJATNTP
8IJEu0/XVA4vSzw/YBzq7wCymeBWqTbvq/6YJseRV8YAt2ycHgbIPuiUIj5kfS6+
E7LksiznOpVSYP3y0L2IeqsoMKcjuwA29LH3vs7bu9KZmCBrLsTobkS5yU9/ANxe
vcqIs32xNLikGe9/33cNwtdMoQTcicq+I5rrRwpbzMYZ3x/pnQfxu1ZeAuDQjI7C
V2YEI49Gv/aKMcY4rr5WpvKnRhPtTarOUYGkPqNbjBDZmUcSh8N6pcqsH0ZMA79T
zvERHl9pUgWwJkPCo89vSMGmgre8SuH3njl0uVclD2US8YG/pymQWWR/455/85lR
1p8ZBec9R+3HirqT9Zc2XasebFNEsZ1/6y3VqT4ZpVW9SgnIZLj9o9vJ+7oelpon
hZrasWmpw47XYPRT2LlYOZTrOt5Z2AlD6/IxIre+Hg8Zs0DA4PUIU7HO2qwBE8d2
BQI/Lh5jpfeTXnKqpodXOa3F/jO5RU31tq4I4De5hL7mJSOqmlMuZMyQs5g57xXb
lNMvKtf9rGvHmqvlrJweP8UX51Mcuz5p4F3644Pm+YfLGv6zVdm26H3y3w7PiDcF
bWvROqaWcVAfQDxPSoflkiBwI4ia/eSSvO7U2ibr/854NXICY3WGBnmVyVKjICx1
a2qz6E5mj+Dtu7huwERWkGWxf4RPFflPie1ue8bprDYgzwWdRnW78XbzXcr5i/Nk
6u02XzHQ92jrtFuXfuzT1tmaXVbz3iBPr1ineKf9qGj1gmnaTKQ03+62EWdiZ4jf
nAd2e5sBnRnfywYnrNPXPcgbxHe4NeFDPTmOhXDp+hS2yypOHEabXXzstLdksVI5
aMl0nVszjtSCjHuoEh8oM/gatG/pHnjB9PQO9CLL151HuaIThiukJ1lgphNwnNFq
6XvEO6xoxGxuhnoiTdc7ed+KMtnl5qS4UInSjcSW9LXnGcCz903ckwNoJPSjgh5u
RNKm/k3E/wmAWYQD0d4gAffjcWgXpFQD93bV1n+eaMKOeZChV7xVv2gKNXW4Tbex
Q7osY6DUCA6kPcO5JxuNmsb9asDCIAtjQbFHScbu+Tsn2QzRkko0ZKZGHBZXgZFp
3bJdkQuIS661JFUigGsfYcqJQCEXmFA+EYzZy8PrAJ55UDkhyuf5FUV+hOvn4V9G
HGD0buF4SCncXzJmpwM8MAJ2wKNJCKzT9mbsCiOIL8z6F3XH17IeN9F4NqW/zj6P
HgQcfvetpRA/E70KpVeWvCiPdY1IctgdjV2fjwroMFKAUWfStvBlmm2lIPm5mWYg
zrcJSW+wRDMrOVsWMQk7yTb5tugNJHT9SDvHrEs1w4ymzBWbNpTzJ9DNjeWJ3+48
CnY0gZchb8/3RN2mM3v8jcACIhcU34Db/CUfKQiNblJ0tIvu1OTxNfxEDJ4ta2aq
3rLo6VFieOPLYwIdvAaYGIPuCN+dipN2rrE1v1FLYjbe982FyR9A3Hvn89sNIZgM
50fzQfJUZxfpZpzexs8uqR08NcSmoH2HsAPJ5Y7xW/nZzKEizWWWJk5sGfwo0N50
IksoziK5IHT7gbQO4fTCxwxw580BX2ksv4XYd+dKQ8AFeN+fJNSJKSwPQu9sFPw0
akfUMribk7miXyq397tJhYR2g51OFnQ9ahckvl7QxgmoB7oUWLVoDvixyLP7sqck
VCU/Ez1WCems+odqU+4qa7i/gVx18NyIFlvNxGGcTvGkcAVTtEBdkETuq2Chwkpc
7WZtySFGBNyY5jayg9/w4HhyDoCUyinsbdqe4NO7d9qIS5wMoG/SBCWiUU0kC8Nn
/x6NlqFWkvrC6sxI79YRqRTM5UB6HSuShqCs8yiVQ9fFWSdh8roqYdwh6wY61I0X
Z/dk1XNayZkDyspBg2S6qs+Jp/OrzQqmDvRl9D+5VrtsL6kfx1qzc6nO6x2jsjFX
y/lr451GpNN3kbArOGzcEMoXJEAB9wZVhTxQBpacB1zMczRu0JrpSBLsEdBbeXhb
GwQ75TdsKaOJKIeowDr2idz2XLZ/ideBlxP72Bjv0cWNdD2Ix5fuB+IVVl5aD28x
zhJJKc8ni9+CeDIQmbaci/SCwhnNqDfBDVVdf12VD9h8jbvLp0QTGV2fWtaOJGMx
U3uCC7W0L21OxOqZa8jy+bY19z03Vkf46wXPsb1pz34d7u5gzz7N3HB6NeGb/+BO
2TrlCP/9gpXa1xUHdm4QWyAQHDFHrLrGncs5BJeJ5awqXvkqvwNLUxykt/pHYGwC
BhrfJwNbTdWyptifg/pibKLIuTOY6s+ibWV+++ZsY8ecL+MOkdu3juc/7Y/IrR8c
cYvxrlxtFAXrXXkc7aJGGvnV2d6uIFy71czO4lk3zxeU7ZXqonUhhSCxH6zxwpro
CdyzLgt0IPEjSafXZgQubU/kbRjXEMUM7wE+QzSZB9sHP8XwcWWhw36y1dWTm2M8
Or9RoHPgitP7RMuU4GPLl/3zp0Uz03iugsYLehWApt8fNzWmdNK0vJ/fEYpmfli8
yyosNUQKgKK58VTPJ6xYSV0VncXZDcsxiRYBmzDleKw2rqXWEexJ7bf5580X2ccp
abVLT2d0BgqpE9UJbA2BUrlqebaZkavzwV8oUCSZ8OW1GU5Up5Ke+ip0cyGJ7unV
EVPFYnkBi39aYyk6n2shAsrCmERiiBGAjvxu0WjDtucoL2NzD7g+tSVvTldlyWir
28+ulLeh7QmSBiRR0IXkswywXsgIggPLXymq9EfKg3jdqw4Qx5cHVYTKIqRFCA8h
W9LlzbHqwxEBVR3JLyIPZWT+kDPaKcezcXxAWt8AHd5iqklpk8z+hW4+/O2iuLlm
FuNvezb5hLdYqoPBO7RzG8roI8pwxD7KfJMkKG0p0/+1tpS/wauDVkAGj7QkU0nm
hQD2YSFLbhwj3HmrJywEFEX7yhVpCRvSBWvbPe6pPaRMNLFhc9HOZdeflEa09rpQ
DR5tW25POEeAcXvPfZqQapm3Nno5uqq+s+H7BfaPhlHwRA7Ey+ytBywdukKpKnq+
dhgBKlTlqSj0bg/gBc6FE1hGlV+VVUVCrxLeJ3ZubL6IAe90iAIsecXHtZJBYai+
pu1BZGCOgSBM+vU6aE0goD1Ji08WwVxLJFJVavv1gcDtnavEIXqPpRbgce3ngTsn
bMCPOR22723FEc+D+NJ/HVsXRnn7XLY54kuNITM6ssGpHTzX6YBiSWg/A3yz/5du
ey1mwdcUxIavXSfSqEi8K53sFCN9l3LAAjchN5ABbdLQ1izRB+dZNfB0glENDETf
CEG9D4R7tbxDTviSlskfiGbSdpNIM4Q8E1BOaKzxWVlj5xhuMyHc3BGmiD5AZ6cC
QQM7uwRIt4eBtmuEFmsqhV8Oj2asfknOJeWSjHIXRXBoWypKkxtgO/GATekoWinZ
FK218AXFUrohs5bmSeizdee9myqKgJkjmIXFbaWBcpoStE37mEXNzb37iyelQwBx
nHKUMOGMlTXAnWdvKnQS5/OqfOGVzHMz7zzbDGgdI0rIVlvyj/CzLVWvKkK8v9xe
t0uyO/jMXfV8AOibyE5fnV2uvhbvNyVgwDqUKScoLqSosY3JwuMpHH5Cna27V7ix
yg2QvVUJyoWJHiMuc8CeyiztMEfD3ML1iIpldAZkXYPpeeEZklxa1yKPgpPr6NMG
Yn1MSSPW8sF+G5DF9UuFYCtMyKBFbg87TCbcr+tjjhWzhQH3pH+SlZf/0HJXWNZO
eRdBetOc1pvsqA2qtjHuG/ZaIqXDtAw2nAl/wmHkcb8kGHU2T7rU/YMU0nk3iXBZ
QiFl1K0vnw8wNRVnwIVjLek8nKsHXJRTfGD7y3UWI7ThK6Q4xHiOPvqcSSE3ImlJ
PJi8Iay4eA6kTQcAoetv04LzH6TYhu4+CgeBe3BUimoJfyKYyRiLPxgCChzjbkbz
udoE+WTXEE+e2+ER0FQ/Cf2q5u9+WEjqsHJ1LqcZwMiJ33rYyLQOeksfLXTQyhx6
r+xoDSCfKCX5ZY7re7Wy1uRy/IL8BrqiVWOQPnt2jvkIHDWp9pHXYzwP+e2C5Vn0
/4PudKB1aPYIGyK9QpkzoKgW45v7RSDM7T5EiUbUdyyYmXgHtXedtAFj3Qt/fVN2
mQiI39pq+dnhZqERLhZE29DtZqBepQ7AjsqwWRdbrefpwYkQCS8mMvRyg4Gv7y5f
6fCCZCCZibx8yR50d8kTTHhdumOk+oUY4rxb2uYqtRYY1twR/T/7pS04WSWWGUtH
apLW16SxG7ZmoIWlQnlMETylVZBBX/mobhSwve1JpP+LQTTK1dIIGzY03b2KMpOc
0N7ZTJ8So/sO3EOW2cPwSz2zeSBv+wvDd4UvzMwp0rMO6Ue46o20eJhoSfTRBiXh
ytZhiDq3lcpdT2Tz7a6pFlK/1iY4bAYaCpaZlKd/GxyT3Zy9XYmYl98FTdBheUet
a7X/nMk5XYK2rBw5/22q3PXlVZuZAwKWX5LNZYI8mj5bvE/o2aWPwt/CzsEUvwbb
ISnlAOWPAUQ7tb/1J67QXpVUV+lHsWN4DDNb9unYxmbEQ1Xk8AXOQUX6oy/Y3TNq
TRG/VnOABegD3w+Fr7OOsPMOo56vq/HT+ELu2fcQg5HJ1fV938TPGWY1VWbU8Lvj
ci3HPjBDFABxRrJ9yuTKfMr/n6YhgF7M4tLoSW+iiz4TFmfcbQzEE3DTgEnlMbuW
rnekETxZDLKV3L3Y6fjVTBMXGb2wrOODAoNQhypD4Jn0X6rmSexSXTeS1ZXdRVLn
x5AuAc+9Wqw6y/aYiiuudl+jqQ/fF63HRP05P3cENohxP1sbRXxh0qso3NyBUIP7
mBq1u42wxiUcFskrhGg235MXxtFAuXpBEfN6WfjJhyMoimHdrnoS+Ha1jTo0lZqs
0CaYrwORQBc2Onxo+KIbmVgnsLi+TgABv6ahgOXXxfNpDt6cBueRB5gM78ZBoWLu
2+me7wQe4X3GdoCBPazFxRudT9Uk9MrAgmwpPkiX607SpKllQMbIchqAK9XRoMXg
09AAPz0pT0WbRjln6MBCCcPlXMAO5EuZzE9s+n4HYsZVq7dUz9l1DzadmKXW+Rax
LTv4goYMAWiQFd+pj1ZHUFq3eP2lUJnr6SHhxIH4rGo+wkJwJMyQ87rsXZcnyMCX
EASO5A5IZArL1qctsuH/xTzBSCi3y3QsSWGRJISOO771yUx+JeQ5Y3CV05DFT19p
ac3S30IM1Lef3jgyVPzmad2kyqde71rnitpX+hywGJTRywViTWtG/CnU3eltN1nM
Us1NOubFgKto6gNp7WFpACH3/z33hQK6hI6osqfz81NQVI9Dtu8D98e+QiJ52t6b
F9dgwJAe/rK6vU3ov/vzvqaDWD0GzsxsBFuVu6hIlFqSHnthCeasSmZjpyexptv2
b3n4PBv4BR1HjViw0/eWWB1DxOzXqF6Mf1XLQc9PPIha4osyraxBRWLddFWltAwK
34MFmPkzxH0sMNq1jYET1x2Xa3ejnndh4lYVlyPHINj72fGj8FobHy5JhJOuBvL7
LqlPuhbYpliPEVKw2irgINrireoFdt2MWG4Dxp6Jw6taYv83N4ae9uIwXoqzcgbI
wXyRPMLFb0tgoAtEwfM5xfCaCpEdwzatw6jYLOLTy02WgqzcCm4ryAJYarro+ld8
eoUOBZmbTqRrMr00diV/AhUyUqXgimfwRU8drwPOhbF5HdZ5PLSfdtVA9n/Ycmkq
Q2ZmPDs9AaVySuvLbK8yVzRLEO5AcNvlmFgAz5sfH9Fn1N8JHiMENnF82FLVHypA
G9BJUGjP14CnXwMr5QFUWS+6pclUE6x3yOcopXCMnY9yZm5qgNG2x0A+WqXxh6YM
P28f6h2BMiR1pF7Y964Pu58Eu5HM7jZcg9tV19mZWzUGsEkYXNpdRVEEV/NFR0Sa
FMrw6HOr64PaovYMhdHGqidtywK5p8FUtXbEnxun+/YsuJBWD7QpYCwZujzBCVP5
vbfjPkBOsCmJXvTTireTmHjHykllSJpJQNjEJaUTuVuJ0jcm0VEFG3uOqTzLuiL0
490FoWaMYpwDciqaosAj55T+YJu5eZ6ac29iIdsNWvx0KcWZN0HLJLCw4JUemqQA
7SB/q34XojUKHuNiSm+ND0FLfdVTKZZFxkQyZjtXzEdDSM0YRrBFRzTJ4Dmp89Iw
vowDZztxJ76DvqxqG9WlpEQEIbveVT9NvXMIliPJoATf0lFqPT5Z299ZuWbk5aNL
Kk5CIRrAn+/yoDfPWFq90P1WhhwukzaB0R/XGVHmFeGdne0LX/c7eYIN0xNXIbpQ
TS55kRmAb/BXZP2tmmGie5nnAp4vmvkgVByinApn4Fk7ltu501e2JSvL5rzNc71B
jzgzVDjgWJfu0ojTYG7/bdUig46AXSIVYopt011SNwsQHy3I1HieqiFP3MbzXMvW
A45N2cj7PZir6EaC2WzNzU4J5TWv5ax7sRc6lbHL16zKnwWkZXTzhy1nlKJuukZT
zjN7BUOLd29ixCzLGX7ZF9xYy8QMcGRObqE4Q3VvLjaKM/Un45Yyyw4nI34g/hOx
JH0atutBX89pVBlG1wz17j4d9+HfKhKMaT2lyQI44Sv/hP6r++xprzxVfdAY3sQx
Td+GGHBJqu+SlkOCoSgaEj3eMKBhZJaVYYJE0YpBEq3ZrrTj0lPoa9++JdD5YL6f
K61I+aPdeMtoic/lT8evGsHnMVQOII2y2P0qdtf94bpTxt8vLOph2p8BCNC3bljP
p1bfkbOxF6oOlGjORION8z69+DFbx31oV6Po/kFPDn4RqRbU1H1k6Z9yWAxsfpto
wzjbNel8oxJdkbuAn2/1cxkV8m9fqSXsVI+hwYtZpQz1Qgnbp84k+cHfrPh7QYx/
M68QGHz82mYeoLjkBSn2uPd7iBgTcyc3OHQWIU1gY4dISfWRMvPW9jHwAAwCj6Ew
1fqYVkdwS76b+UfbPKQ05BtKJa9nITrfaC1fQTK47NG2t4PRgdgf0isEWEQ1zqLX
vCOPcmztsCGpHRtrf3PAt+0V0STPVDhx3wzVMQmUkqMnh/NpvjsuQ/aqOgpX0iIk
z1J1kJVvXb+So0SoZGZpajVRId7H6INSPjItqtmvL+SP2WKxVXFe1z1MEE/PslMn
JQi0kDpb+5S3JK/H7bc1/7Mxoj0nzJW10nQxBtO9X7fwl6uoLKgXJAClR2SifiI7
y5sCP9DlyDP9y+GyEYMm+8qDQ+bDJjkgcV7Ig4fhVmPshq2GbzR2JYPFCzJqMKqr
veXFe9dmbbo30GvmXKFgddicBfeHPZ3YfyvFX9QOnI3lrqKb6D/dBzGvpLA5DAyi
iOD5waBbi1Bb8XSHBE93E1nvvKNsojaqKlLvhveRARWRfg/OSDNal5QQeVOjsro7
NKHk58AfEkA4xhRIMPAzNZTNoUxwEew+KX5w8JXEctvXiiwRwnFgArep0JQ6K2Cy
ioNYStoAnzxb9zUuMJVuWJ89K1kbSDs2IGeIXUOXe0Di20APAgixZ2YGDKaqBU5a
waDU8RkKZS5qM4GFUn5AO3hr/E4HInY29giYVi2bhLIjBnLKc5Q1+aGww/64YIoD
H6VHrJv/d2O4avC3aEJo/988OtakvJD4Gvrq4BgIbmqUWwaWcylSjm8vk/K5fj3d
vX1kwuaIepITrV0uqAqg070eiQTcmOTbEEj7dVt4Tzel6S5sk2aZznP6V0GRPb45
UBdGR5g/CSLJq4yn0xuPHwZJ4ViMD0qDqCNhvvv1xH5+CKtbXTdhZu3DB+wSkTbg
1aq/TTYBLSndd/WtRY6hj4zrojaBoXUq4Kp1elszbZ0whM5S/O78piHT4DdWwe30
q8SWZTY3qD1sAq3mFv1S+tfTz5kEKf31Z/TIfFrS5nnASbdeeiGAdsBivNDCYnGZ
WKTUeDM3qFDvW9aDEILtpDwiIXq8BMHi6lm1cNhi83Z8rFJrPY3zPl79CT6oVhzQ
2VOe8iXzUyeR3NQlPQq7Qvoyjp17E+EOJ34Dwi75iH3nnY5BrVpFJ3cVO5wivdzE
BroT3Nmb3C6j5BYVqILsl0a3WO3VRGunUutu8S2yTY3Iu9TY47v6KNmZqjyhByt8
vNk4REuQsPlvpA6iB5N2vuTTiCCpsGEA9rCCftTY7tpiR976mXH03WOvwnRX4YjT
27qWN7xi/hT4MdtfCkUDlnjkz8SztsLsnj7pcg8l8XTnOHHY6cBzzgfyly1o/yDg
BO41Sy8zRkCGhJ69knkcl7zQuYzUp/Kia8WziyNUeSFmLV6kjLPS9SUUOQQ0JnEH
jKimsqkRCajn0uAu5U0X4+o/P1Eb3dYHftihuHQmzhTZvJqAAdqoAcpMSKzMUy1x
9Gjodh5gPh9321BAHfpwW/1fVUUinWMEZ4mbQRxAE4VtqIQsXv7ybrqsL6h8dlTS
oABgjEkG1gsf0XNe8yoPx5R4rz+9g+8yHSAoCkvrNxoIrHI3D/cQegi85T+JL1jB
eoLqm9wX8gvZjlLwVSORWPCy26TR6N1VUWotq7EEMzRj0lCtngtevp19xyCh4aSi
d6c5u45MGXnzDaBMoQijRtFgd0mLNN2UKK99mOu5IbIczeA+0gFTBsS+TOtGmQjD
6OhLl+Ph9YWEuXROKL6TS5IuJl2zosmjbdYaTuHx7qDTODrA6KBcIn8vGaSNUL14
NtMb5vQUuHV3JMt77XKsN7Xao5kiDgz+/O9MGV70C2m+woiZ3aWlJA7OPyD8VQUb
S4evcFPn8EIom22NmlNFLgFc9mz8eYxUJpTmWMeDzBQZnTwZYhxNqT2Ti7H4+IMz
snwe/k61Plgap4bJ7EejkI8S7xpOSOPbJvGURxFRPVLrsVHlEvK7ZqZqzmg3NDEz
wpbtwYnhd4WpHQjE3CiIly/fT2wwu9nfcRpekKrKBK0Y6Rswf329gB/N3UyyOiD6
UJhJa6KozCKfGRJqnAIQNLrOmN5HX/zK9WX4tB8KSZv9FOv8L+Y/l57MSCJIwPBw
xzLPAHiKVwUfm93eEA45Ahd2lF5gasqsSixNnDkN5YUVpSawrtayBE6sfqyqUCxF
eTGJB3F3EKt50hp/tXecawI0cZDViOs5FI+XRuSd74pwqRgiXQBy4N5xuEGPxW8W
EiciW+qSJezp2yJX4C+xYHDk34kfBWe55Jf4kp8BOCCl3sUJnE0xoL/6m+r7HCLU
+Y9gLoy0ZYNb10eGKiUwFfj9ksf4G8FMu6JOd3ASPRvQ49zOcoq1IASbBK7GC7MQ
Z1y8OoSLmjWvID6VRPMLR0aPcypEpSLaE54hLByCOuAtZF6mGxPjBvwFQ4BQaGXB
UVL63jlkjew61lA7Bz1AcLsJ+nWhcekgFJcu+x4CQMYngGNz3QSxMBMl+ee90ox8
vGdbpMGgdIIkppryCLyXI2OAmCuoNV4MHM0dCt34JiR0tQ3dra8VDhpwzcZv0Pra
BYScwVKm2HnLlawXj/jYzi8cxH3X4Gq2V6dH2kuJL85BS6lAB2j4lgj84Zzytu+k
Lc1oUYFOBDwYARweaPlk35hiTzX0FyY2tkj69+PynfNNNNzKlEf+tZJS/Vkew+PT
3gnUyTX4cF6m0ECS1xX2Oa4rXPY6TRJ5G/Zb1gzmIUBr8t0RxdjQMUpimUXt6s8h
wav+pEWvAVI9U4zTdBJRWwEpYLMyvKpOVOmXmOiHoYQO5iOjNC5zjjt3XEF8FLzp
v/cH42hjxJRPl5pqCASM6GEIaEBzGhEeUZ6kaLRVd2s5sE1ulz2/JbDvoXWjB13e
kXpr997Jhu3iBgIaXopSnUtg6bryu1qatsQhQIfTKiWzby5nBhPlS6fViVTgUzDS
NR4cl/3ygiqVtAi3gSoPLdjxvnloA8MMtG9oq7ztpEOztjviuiuRtfWZ/xCFMHo7
ULTgmRXoVhmq7Ui8rlWx4Wc72xQZtFzoBHsyQbXtOIGzCcHJS5Ouu3ucd3SB2ydX
L30WBVNLeo7eIYHaeVJZUnac9GPL4wzvhWUWLD6/C/5CT/hO0V16ioWSMmgV4FOj
8dheO8aRh1okZxa4mAiv5s3/9ogIz9oaoJxLiPkjm/AQ5OWujOCfxhGMEfk3YPot
w4uem2IMqAV/5X0SIXjcRGo6afY2J7JHtTMZh3qo2vtorzRRgKJNhvpzVkO3fnGk
NFWmxxaXfmGj4gO3D3c9QhrYwdwMfhv7xGJpnnxmeo22+HvB/G8OHJ4AR3WvGPnB
sx+ZSNHt2ZlyDD14QS0HQ44FL+p6MWgjS5FUXcuifyP69DEKiJwdzn5BKC8HF7t/
0fKpdqoL4PUGWhXkrijRLj0rYBe8C/08WyqCG63Wo0Aorli4lKGVOemsmyvv6X5y
RgBVE8zjdNuAa5JH5hSyK0X4pTujG6w3T4ThqXh5SEdpaIueaqPzo2cfcw42Js6k
Zf7VtpFG2aY9pxam3q3Z3/SSp8d1AXX/hIhjQc78QSLJp482dbmjYABKIaauMBRh
LH2B1jpOC6JiovQB+3QA46ouoYVHVPtLk/IEbaeNBiVjUIN8KuE6v8HQsFK862f7
hEGOQ2c5ywV57yx3G+oEGQhNJlLhqvgZNk0Ffieoi5ilZBDKEKUmp0khQcL3OSfe
wwEbttM+UJj+s8aFhYzrind6iXVbcjUWgn+ZiYKDxTfWApodq3DnABjFHEzwqpFK
e9TqfWOFWkZgd9qt0Blbq0xUpkKGQtX6mZSqhiyejHJwj7JjJDchpousXFBZTY8R
LrQyE79fZfq50Gqtvzkds4UEFrgOzCaTMjXHIIceyI/E6YLwt7cvLTO+G9LcLwCw
wiXBqnL1HL1oz3/DeUUg/LzCOchUlp3C8d7agbiZcCdVAFXeV5FDOjalfWjBIhW2
Hl9u3RGw8izx33P7hoxw3FgRIHkyRpQgwULx43LoeLCXgOmhd2isZNTmvSL8ffuT
3frBdOLqCvjoiX5Zpd/0AjbOEbBYfJODl1NYzwNjjyuXTqnRYlv/EdWVxvXcNuPZ
J+8eCqbyI6+NwbUdIDmGIUwtasdTn7EiYLJCpMCue9zNy9HVXeOCnEapA1cf8Ckj
jrJsvju1hUbg1Nm2phuISH2C3sPUrRnuSXY8sUVvrB9Irvk4JrqUBV317euF/oX8
c8+64PtopoCYVjgUF+T7F7ZBBKxjSDkbjPtUAqaKByM5jPOTS1drRYyRyeJR95fn
HrXpv8u0xL2HSWCa/yCJiSPJon5+mSjheFqfm51iu2rCRhh+BFqRgEigdLjdmz7g
arf/os4gS7CmNDbxu6SPpuux4Wx5c0qT20K7+uRvLisblCb1amvUdUquFJeHoF6d
2WyUeIlkseqX+/57tieBu4wzvd4cuKlICMzbwMNwPclPQLalJo6KBpg3y6YN1mXF
Xh2GVmqk+4NOXCloyoQmYFzW9GX46rYnu8/QIBkzXh+SR54q+goLO0/h3c4qPoI4
osJiPJudRQUi+FYYL3pU3YUk1kM1W5PKntkhSwexoZTOAUcLO8jF/3Bx/K3HTwV1
kiZk9imCqew4bydfXyg9Ft2+vKPORZMCB/mnUdESigNA1c6ggxyebgLBc4JJuayv
8osBNU2QBuHUbrCynCx8D1MAs2JXVmTzdw9ZupqX7RoK1cvJHxbDO5D/baxlznJU
vcVEbTlXW869c/8Mr3scL29fzJ2eeEKAiaaS/0X4md/46CxfdenbUQ0VLA/tHuza
L0GcTw4NfCcku1S8MmnWZasZ3+h98YWFMO1RkZn98TPrjgNdkRAcRtgvqHdjK+K+
rg7oI8dhg7ADT5n/k3SXILX0MQE6orLkEvLxN5KKT6I5CDhrKyrsSnIQUfuFuiiQ
ivqUUZDIXl0+Vug0xU83sZHzFZXVc1YVd1LHegcKTXSOS2e6A/BY/vWDXXaCgonU
h9m3CmcBWxoYUSlRF0N5cfI1H9Dmh/ijMctG68h4eku/Bzqc4pVBLu5dBt8pTe+C
lQTn4uJ8iskGEqwoSWAHGBjcu87KLMAGCPusQhwN1uHsPrBiJ+1UcMtGvbzXvOXW
3IOgN9Jcu0GIOh5pYWATetbzRNKcjg5sO8qu0ez6oajHdO647U8cU0FCHLuO+aa/
djnjkkSaI+Bhi/1HmkD/S6mTWlsmovrfmBqodjYXpisOIdxF0AAWuZYkPUkb5DjF
08tO4CY+0qZHAqCmtC0zTZuBI0BmgJX1WRHPpe0+IFHyQ0yTtH3Ct5yNKcDM3ydE
h9AND76FORi/MeAxag4PwEMIBcu6C3kvTnAyleLvf+qQ/Qr5lnOZRYd7aQ1NQ4d3
bDf2stQ8NBjk2CHras6K/QG6xOk6Zsag8vriyeXuTZnonWT4eLLesse1LwhZnNHi
rFi3NzQUiCFZeuejpnoHq6vDiZsoVap20ntHKQFPkf+T93JrtrJySMWHpXTSKxdV
ZFITLxxGyarxuIedkIQ+Kunbc2ZvzNhmAxD/PQh6pmedwhLb6qApD86RW9bXh2s2
0fWtSp/OMfbbKCwj595oJHEzczvAvlI7LJA8eGyJqUjBcbNbAh2BLOzsZt17BC4r
a2+1wCZhIc2Q9O7l00X7niVbs5y6BGsLAboZTVkjlK343E3zBx647/Tf2KAvADDg
jng+SUB8w1QL1mptU4nFwa6Y63ymvhQIhurA3CILr29NXN+TGem56PwzUMNqXs4C
25pPwqzi8hmn6zML+sztCoRFqNrDLZWLoIGsbwMDpmkrEIZcr7gQ9qpVMa0kOG4W
GRjmdFCw3/FdVaVBQF4miU5hyFZHEjCsRer4OEDl0WJtDaDm5WtgFVG0JjZOBJcL
A5PFO3rS/0roOYVTfREFeP4zggkqacuKeGyGDdE+Q+NsIYQLdCmHzqBw3T0QpmxQ
2+fcxgRm8xNT39Mv1MfdXCqCL+DtOercArNNlyzzPmdZ2uSEpU7JmQzdAaA5fACX
P/0qjCLzlNXPVvcDO4pKRhsCaecyiQIaHRX2sUYJztQPoqgO/DTjmaAp0J/6jnbA
Z+B4wOzkmtuAGGzIHSBPp5FebzsE26+Wl/xVshVV1F0qDaQIISSiepP2kEdBV46Q
+hSew+tPQOIhkY/o3sAhDxwvW5dkcLTP8fnR08lvN4DXmYblnxlGYhtJpW+i3SJG
VVqS/kIiyMUeq7FOd4sVIYT32TrQvXd72wR6NGhsVACpA1k4XvSEvXYXHyQ4m+ph
wlgakMjp6HcMpBAeGxBrtlNqpSPuOsrqDekOWRWispnS73NLsER1C5/HxMy9S5MZ
p23d7ZDf7jnDdHzWYNju3UeFMrH4JlUQGzDYJf+UNccwhHsYcLbaXKStYT9/3w+t
URGif6HY+dy/R/+JRuhsoFPWimgpSr1XIhS8XI3db3IMdURoEekxechD6M/2eLfb
Nqp1AHfzv5bvMhFC+/f+uLDOCBN1tGVdptVjDGPhfUn6XDrkevakaHs0ovFQpn9N
b14QLO4aaemClzLyFmII7yy2Y375kAU0rrXKGf3y8u8ymeN6a2aaI2dgzTQgPz37
xFB1mB8D2HBn238JFdA5uSBdkm7Ng1q8NSUq+UQJfJpZWvBv/5NBcDHxy4v1U0gj
gdhGY+tcMoLm+oZzmawJB8sp272pP3pjpeYDff10fMwW6hARekaudcYWshqkVrQi
gnUH2eIpcNRzlRutNIBIfjUOSVDTEGuQQrGS2OENbmyJzQBlPOZD7UKdFL/j3J7+
WRnlrs5Vznecs1hUiIkSdlIdCxLt/by2ZkAEf5plU0rumz0kc0aA+Ghnb6yI0HAw
XrsPfL5BVbnjP5EgVXM1eAGx8W0vH2jFqnXg0GGEN86ciP4t5dmObQjGERQdcd1s
/o+M/NoBSocssrSgWDjFcyMbayDr5Hnya+G5Tb5FhaDU/4NPY+S6F7/+2UL3e0fQ
EoNs+Fhz8ulRtp374p+QoDd89K+oxKS1j0DOTzuIVkn9JbNxSIVpUz0yQ2kos90y
fyldlPxMpO81qGTvCuVIbbkGmYUDf12i4EIsactBetD7jSxYN0uMxBAJh19zKXJ8
lT1+PkWn7U23M8O0A5A2yKiz6G7aLcn0/l13d+N/vqHyVb2hC8ESfapDgOxaCrhg
5GcXqpdOR95SNvGB6N5sj5TrAsIyRgJxtS+/mGDUuwJ85WkBQuPF5IkR+LRzNlkq
V2+EPk6ix+ebU2zzR0wY4MRqm61Vrv63QU4Alx7EiMjzWjC2goXM/wC5SaaQE0Xs
LeHgtEFZBfOH6rC3N5ULzYR6KE+KdYwFgfczDYV2ec1pYjfgUdwJ4dVGwXPCEO9k
9gKJWEu7FmTPzZJfqhxj9mcsPc0biqOSC7EJ8aM/D4Mom1ZHVYLkucM3FxaL9oFT
UJiqbmnwV4XbAJjNhCbsNerpir4nyXifO4QrR/5ragNLXXTbHvujoRdZjn11F4dW
z3pvIWwuttop1WUp7/sWDC+uoZDbnFGarWgeRMMsmGKJIKdGkeOHXCOcDZFEUF3q
f74fqBzrhgDp2N390Ocsb2Lv3gpsVKnvjYs/b8yRNRsRvsLJ1HW1IJnB+HuRnR1j
1tnl2Y9I/68czQyZ/oau9XWqlgol599LU5050SYVnMiTHJnAQ6+5eD0JzZ2MT4u0
4nbB1h5HBDGMDS2DJ10MIYOa8n8vg+0fFBmIstbtNGd5tqOZDanj0pzfNTKStzph
IKVeXQZWEN9QIUz30k+cIU3ejYMRceJdCBZRJ5C3KfNgtIDrdc3mZnX2G1/F59wS
gvQa24Ij5GImoJ3vsoGSSWJ1oF2a6tv+Sx1NIO+W8XVI8LEusWwjt3DHphxSY56e
FM7XUbXHkdjHmULjUzjr3qO3ospSXrG1s2kjuJXxEN6lB7gk3r4mABauHcyrSqQJ
DiGG6Sbga5+6EwDcus7GvkQXx4ZpFYcUhtjgwKgnfeyhHdG3r0cPzXYa1t0vuFFZ
47NkrYUtVXVkAqMrpllxZR62Dn07D8FX1jTnpf6UktlkisyksLsEmCPZXVfMaU5e
BQbrX5+/KENHG62LmGCPUuIKTtb8KrIXefc+ekUJcni6MgvmXme378XTSy6FxBZw
d2diS7/qeBNSkT7CAu0gT1ekLwcFmIGmXXOvMddeYQlTZ2UITSbudGBvA0UGxP2T
ce+BiD+5ResnM4p7znU5azRCKdfFFQBQXaxwiyGBEfaC4JM3+ibAwGHzvxfj19nC
LHxU1bPCLT1nJNeWFNXoCP9IXZWDE7mtcKupXL+FIDJAYuP99OpyG/GNki1c9zN4
S+JGcFfzb0QjddyWkHncaq7g57DiVilDZUlr+6WvyrevAj0al8HjZKSpBBObIRwS
+Eqg6KdHwl3+OKzGdlNuS64TZ4naWLr5pOdhkCe7Jk0AQZR4zgATG2BOiyUoQtKD
b50p+xJqEiPjTu0oS9Z4jmZNrgdPSEO4PBDaGCqHKSQ=
`pragma protect end_protected
