`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YSXbbhtRWWdTJPSsWBxNNBMrcnXucXuCsuUnYya2rgla7Uf3p+pboAnYTrH9Ve9Y
TnX6GMgSSn9OEhzh4cPPLBNgNKqYMjsfh6wFEd9CeBbgyCIwHfD3TUYVyYeAF/Ln
gKmvfAah4qr2MiS3DY+3OzobHXHq80YWHWQgIUHPH3U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21680)
uHnw92qhzzc3hDt/3M4UL9r2qgaeOyyRPgJ4JCu0KITuE1evfKHETTDezYKodx36
mc5Rzj3ksNZxqcEckwInOM27K8BjigGTbKvh6m8LoOVRjhEkPlwwar6E82kGN4hJ
Td+ZWkUWSUxlle+nU1wDVdsFd9grlIXoA46x6u5Q+GeQYhDHLKbYqZyj/TMT5TCt
xVH4Gr5FXbJ6fEVIJEeWMgbWu5ZtAyx6YKI1iTeeJA1BTAhEslJ++kp4Ohagy5uS
Y3dgexXrx/q+vgwKR1QiNIT2hh7SYRdt6OkJkiE8esdFG5i3iRC2Xh16oDolu0/1
/2cc95R58ooubr/3de7G3nvoGVH7fc/36ZpEVeZv2xBXL9rTEbFWNoBUuqPNvGTm
2AAOL6RI8Lq/BEW2ryQX0PSO5QAQNJSlySyAALpEXLi8IYkJMpYOiFbzNCR5bdqM
DKEszMEmM29EQfXLxr9nhKZ/OKSlNlx6Igm+86Oq6bDxDhof1KU7iohXdafKuaGE
tfy28rCzN/qnQT2K5oF+3R+2YFIjnvM/nNS08bbt5udmWqwFT9odk46n+ZdgBBY5
qX+Cfoi4TKuwMp8JH6E1a1NYKSXj6rlsXWV0tf56fXU2eJGVLJnHydXIq8lwxkoB
Ebxtga1eCm2qJYgPxOnRaGgWxZW8KRcTejyjefQtkD0N1TH826aHeMeMyRIYTXxt
vz1tAOzKOdLO3UgKV/2qI7dnHD7Gf13vYa6hxnJy2odG1Chlcyz4YUDGBqalkvr9
zsc5EsmQp9cOWkpqlxSmXY5tn427J0H7ClzQBOezw2OkY28A7+yzyvZ67nCCWLwT
T2berK/VN/WzqNtKkutKuSDd0crtp+Bn3sJscvvDxhmV/sFpYzV98ElL4InnmSdX
TymeaDYYUJ/jH0f8s1mPHpBXYWYmJUhfpeT17zZiWlvZiCE4ni/nd2zo+1u0dVkG
UGdQ2APTqXm02VwAyasxes4qGTP8uj4QSz1W/+wRc9ztuetN/uvkjIPssigF05Sp
h3kkvicRehLaHFLdhrkPsAofAchnxSH/W08vLxMPQrcikviLK0UVJDxDvUAUfcAa
LBiAorIypxOhGq/GW4MuK2Iagq6l5EjcZmOzym8fsFwWkSkqX6/mxKX4gwn7x4UA
ihbvDJmFo/cubE9mBrsGCFzQZmxYu+O4Mxcp0ZQ78XtnMQu/383FVzvrct4wnjPs
suPZtAo8eMBrJAk56oj8oSvo3JWh0KV+ngdInZAfP1sCd6sovkaFtorP1vcUdWeG
XBrP3zOC842khtKp9pGNqs6Et0JNyGODlUkrl9Wftad+TwZ7N6FiymXVVIx0usgD
6Au/EQ0Pf3263rnZRJbdbuk0gPQDm0vL/3c3NAzUoACFbhmLS0IolG9msdwW+ZNY
RsvkiCCL7JsBcDVQikziw7sw5UstCcH/V1DTulqMfhQ7r4F9WE9tJfvLwQPPjCLb
ZF6RrhvKMKW6ZiUkmTOXR4GKr/xEHAk0+gDAe6FlsNt0+zDU4329ipFwO8l9HOLy
vvFwnFBU3i333zYEoMj5zy6OAZOqcqmsVvqCiFyH6wS2lP4T1akyzeHFIg79GjBf
E2x4MPenDoAqqko4gBFv17kDzmGe5FCIqmhQ/wl4DdbWtPSmawXPbVdFeTG3se4J
wtBIHrM7NNtU63CklNbFBTB1iZEoSQymVcYau6Mz26UXzImj9F53CWN45MIDacix
7KS5H+bpBMFGCjys1ARfR10UsJJkyYAu2+6gOEqJeL3NxkXdKPE8b8r1SOzhW4eb
gtEwd4nQqV/meXYxrtnCos8nBqxVAJvndQkZXfyRXEmn61k3C4qtoupj8Mu8YTd7
uBy+qL4DINArGsgP3UDk7FFhrTkqgfVkf20toYw6EDvkaxXlCiDVhdkXilJi6GW6
ANFfDqV5mfV2U2QFqcmKMBfFMUwhcpf3D9cH9FOUO2i3qho68/RwVKPMn6ShSXtb
SeyIm3gYMHSFwRFFtdpTFjKoz/ERngYMYqsUjtHx7fwon4niZXMF0rPWpDjzkItp
WhGlv+nZjW85HLPI9So8HDJgUy3E+lCB84O0Q3NNRxl/ImliVfOGdf3xq3c7+WNA
Z/FwHwvzxFhTx+tb++wxbuQyn+m6y16QnGzKzJaGUsTGw0NliYg8WauOFgOndNNQ
QBnv2gWg2ZHkMr9Xcc/FuNgmZFPBeZm2jx7boB6RKbLzMjQF4hY9BWAR28Q/XlEo
RbXPhmBcmJp+vak7nQnH52JPlGQZbcRD11ooYNffUzPYcc4HMTYs/wqOk9hJ9WBu
evvKJwIMbIBu5x3N/qVJRQZ7gz0RIyN0/XnOBqcqqgcAmJynHafxtqPp5Wu1hhHG
NHIOii/wcdobf/YUIfSS2K2lzlXxJ5dU1AtCEWpF0rQCdvR53NKm1ltZTZQ4WD5T
mG+Lt2Vw0F29iDrpXD/r/BR41VqQhrnl9jx8NwepNe5UXsCPs80LMQg6is40MAcJ
9WXBMXrvfYmUBwZnmt2vM/v70suTX7Z6hjg1DPvGt9EzLELPWZTpA4Yz5UaT0qRC
qCCpJtdCUJFatM2pDbVHVv3Z7snvamtPB4+IUOvQXqfoGkJxRMaJi/BNueGt36+b
VlDyjlvfjKlXO/6+QjZrxnVD/VglnSTbn69r5bdyKcHrVv7nxJ9tSOot7fQDKFEG
Sp8zFrinfJVpEJ17XDGCVPTsUPkVwSvq2rBy/eN9zcuYoPqTWtLsFrKJ9lWetp1w
zZ505C3vIA3CM4isoqpNE1Tttp+MeH4+ytexdIbV59uDEVapg2wPL/d2mGd9ns8N
ZHauNeTueWJxM0Q82Ym/GXSCq1fGz8W/3tPHPZfvjEfG9QaBpvtJI7M9TTweu45a
D53brvLk08xr5niFFd7u7f3P5+pNFnFK8JTa/sAuPTfPMtOWsK20ZDqbdZhIaSKj
KqtxEY8TwHwLi0CZ+ijmUptOD4+i6GHTDqPiK731zPp1pGnOjCXZR3HQbKHzQKvo
x287FIiVShkI7WEl9Qv6HPSHlSROzPfoF8vKDhALS4EcHyw2l669qLDfo9wlmYDr
R/J0B1+vp4eyEqpLqa7IDS3RYWpD9VHfylcfQCg2/cH+UM1mu3zY5mbHW14AkcsT
MVMU49v27g0uOZ0r8hWSjBK87e65QfTwQ9YuYjycE6c0qg2RmxPc362Zf0Q3hE0H
iufJ5aWfxxal0zfW5apVdFaDurCR3DUzpKvR15XZL5BqBfcRUk+p1WGaYLb2EqDJ
HwUMxt3JpFWoRVQZ3sYUIskyBi5cBWgAtiBAzsNdgpx6CVyE48l9YxwvHrNELnqa
/pSBZdXY9FBLg3/mJtZHZPfwh/pZATH43KuNykEYAFiShTzYH9VfGJyDZgeuk1rP
IzoAtx1mYZ8bEDpEutYO3k2BUJ6OBCOzeuLEhVFkCgFo3gR1KaZrlE5dIO1BEZeY
idlR9UVaYNo7Q6XeBQrGRu955KYWwrviocylEwlLd7GvG9g+xmv1ktf8P1ZXCO+8
4opPdiNkX2TwX1gg1a52rS1f1aBCZWj9s28wa4YZ4ftC3Am2k2fIzKvfvxJ+4VwJ
degOkW+cfMyUhJHoPfA5Qw0ygien2G3b+xfx8f5uKNc0Y9KgoXFG3OsyajigmwNs
Kux4qduCJQGH68AuXPFIv3aPYnG3lRJQZpNCDTGXUCqHSk8rHI0+ChILsP6oUP7i
WZ9skiHzBac8hCzWkuz6YS9CVpm7czmv5ogEhlHiFcli9IVlH1wd9XgrHOBUxOKW
6Uiy9DOnmx27i4k75Ii1T8LZJXi+9lgwYKnb1VI/SLd4Rq0s27TxsR2vdWOAe7kk
ZjdrvyY23d0lOd1TUunQZcgRh5ibTnPwqML2puyAqjE4TxNaIcYO6IsKEFrgm29J
dA8YfStUZn1AMdmb2/NNObN/L+PAo6Y29uRVEpzIYcV8JAOkNEK5/+pesS1qi1Br
DzFsfRzgDkKuC8vfPhY7Buyz1fzD4MJuOyWdpSDkxmfzwTwOJR6B8/oNq6IPpTdU
1qREfvRYkoK+xfxqfKySWnFe71fwI7BWO8cDQLSBRoQZHDqzRuMRyHxaCT+ltrBa
WiIpJhC0IKYREf9Pe6UYjhGxPmPd8mmqoMDnYs5vsEpP+xtMfBs07ZBYaC5vDvdy
0R5+6+/wzOCzKd1UqG/dCkZZijeShYyZhF+MyC6SHhisCdJXAnyeHDdWxhdi32ne
Jpu0VUHIYSi4yVmTgSpzorCm/5ncQ4LhXYRZa/v4LHkf1Neqt1DzbjpmSOQdJHN0
wLlk4dZr3aFCOMqE91BvJdTiiMkMiX422XdFcmeE9vnd0rEgIBdfgTWx6aSE14oj
p07vJFLm/702qHD4U+9o30GXpHY+1UuK2UxSoVZJ065/BZpjoWup7EXsbaq4yf3l
VtP7g6DgJ6ooVo99ttI/7Aa6vu0Gbi+uQBy/hYLcdzWaMtkZMDdwrXI21L5tyFFa
0c8vcjZAU1/j1RLZ5R8tV5izK2P6F5GQ0+ISB2dLhG7sqpk2IqeFBYwkzGsoA0pJ
AIAiPh9MQ4mEAgnfBOZ0/kXw5/UlzGrZcmNfzk0qgGRxXAClyYXqf/esO/iFycts
YXZ/7fw+sKCGzi/PqHrrkBT2Uj4NAaOpX/Q3NuaYu9QpzrBJRb6xveye8HxQnYBH
0PZbgtW/zEASnJqMllZzTQnd9k7ELtvGZc37QpFeugZ6fmquDDI/XD4ckObbR86L
fGx5y5yLOkDoAAAk2zMMzdmrab90LaqQlOeR0x0YgUUH1HT25JNkNtEYmd1DUg4o
qPx+Tozm3+pxUxDh33Y2UOnHNkftHlwt5tnEyPCYqahAchii21DV+RnhWWn0JC77
woIH1a+CfXLXwxMt8yngbr1chV2CcsLNAFkNOpyy+sq1FPuC7LZmCg6fE4t7pK4H
uEiSR11grI+RENLy9k7Jr/lV0d4rewbtuTDsKeRZvdu1k1frdFSHZeWlxdsbNecd
e/cnlNNONiLjnk6QO0LGvLZ0XheCJ+JGdf7vInqhKkedpVusHK+e2MDpFWgrQ4Jq
XPAeRo0i7xU8dwJU/8RJ6u2HYDxF0AiI7aKBr8KcWzt5ynY7G+TSUzL6maVtluEc
HNHzmpT5wB6Rih/S30Z+815h35pYWfP7XxYMh7RNyjeESiHyYNSkZ1ZHlIYWdUEZ
m/8++VFJnd7C0ZGa0MGyOvD/z8U1rZE3aAc+M6kjyh0ncvFmziZVqynrAv/EGi+D
LoRsPA6aVT0+hGvRpCUKlqRejHWDub9nATZYS6+b2D9p6wxOxB8OlSFW1DCKhFzh
iGWmzLfcMYe8Cn9Py5/halHqguR7sU4Y090MinmQcLOCW2htnBEw0NyM6WsE4mcB
q4mfrvuyx0VJ/9xsa4rsdDntKz8xhPDDcVkAifSkTy0tHjfJHc/0X2zmow44iBWk
agmrI9981wE+4yGem3IwCbGlv31QWCTYemSvjOPHtKXNX8sQstPHgbjtxhf9XvAl
DTVjpGzdc0X/HIhuLbizSWmrLwKJcqJfL+S9KF9uI8A/Yee8wtoHlLSHzWAzrD2R
R6HT53f48r5qbOkCRDqVcYtP6FfcfNlVttX/E2/dM6sbjYWfLTL/d4/7sO9Ar2RK
W+RbwRzaBIetaZwxyT+0rjNqE93F6HyHOAqjtS2hOLvPB1nzlhYQL9+10E4Uc3yR
Ot3yQgQPM+PVM6q1Aed9h041QhMfxZTwdj/stdGI/nXQ/fUjTI8BRTxP9aUZI7zF
x9B4LglySuNWj+DWxnIEFCOq3lX29QUIZmV6cS5GnykBFl3Fqp4kXA8z2rvkH3Qb
HFOX+eDNHrMA8rziu8R+RGP5jOkUH/QgjpjJwSFutxWxGnbhkJ1p8y/bo5qf1J0k
yP4bwa+1EIhV2LIcGPwTy1tzRnilyOHwfd3eOuoMhT1lHC5ZcwGz27uJYwM3JNqT
PzpdDi2cxypnvimrCemfFhaMZPFmzNESgNHUCd9bXuOaDwzKdfPMViDuW1TOKg5l
E/TA2QCGMmvReGeY6gWITgTz4BjJfWTtkiF6ddZSz+ynxy7dSQQGyHNSyCJLN6U1
cFeJgthRp53XVvRg1KDRvOtckbhaXCmXpCmCzXBYUV7OVe1AtMfhBLLLk5RHPuXL
AwRkaqMzOQ0OidA0ElTlQdF1d8m8avaOKATJq0sNMprGN0TcbCFVfxUKveuvCnTt
vxt+Gqd7IYMfWTlxFyodktd9/hImbJKOlkiAIVX0CTNBrG7uW2MRCG2HqpO1EVZl
9+hk+WFYG479UVB8dMsh3x5aW3Ec7lgHoPDXZEhg1EYfkTKtFICRd+vNo7g1UVXW
IlBcwSoBihhFbPuoXtIJ/xRdUCKKc20qKbhoML4rtOxMJSZg/0YJ/luJGOYH/3R3
x8jJ0dBrfxo0qAnV4QYnW/LXDvzFpxrM0b95pkBXp4hz/9KVqVw0xPdOI6/PizIL
BYdrpIy1agwClwc5USArmSJG0R1/KRSid13WCuvSfNqcPUSxuDClibD2hsVDrn3q
ZLVyaw1LT/M7bYbEo3F/p1ZLR6QmHgqb9WxuQYG6ccV25H7NCJj3BgGRzKG3v8rv
NYQuYZskS3Dq58dwwpOu+qzaYeDtWCXkqjrlZRZECuUl1BfgPFoBmJjgdZDS90Ch
TiNpoJL8gPnJJMb9SpeCKaDqNJHlitu3tKBopS2Au5xW15wFpLXaaSrn1ZZXy6fd
drZGXPRnsbXwlN/Z+fGQYcOu1qCF+LI3Krx723hn2wp+I5iV3GzRSNK9ttqBxaGz
xOcarXKCueTO0cwLh7HeCr4kMQd37FMihfQBR7Q9dT+lDL7DQOG2syT/S6wN3Z7s
EV9Lp2eGGnnZ9cTrOXkssPsGrY6ak9ym04OMijjoBs5+cGCLM9QkA+N2vZHoWkY6
3r74iGojlJbvoIaBhhqoVrdCdRgr3UbMt/rzm5ybU8LLj7zx/PvqHZ7lEH07SaNB
eXhzSw5l8nH6Pdc0PsSJ7tTCdENMb4FON3h/qdKwdas06EOV3Ww1YFgcZCkNRknK
vvsSMg1+doydMPNbtjfbZBxK/X2PxCMSLJR0VSECbX914kxxnQ4LdjHavScA+QBl
fCgtQIh/ng5r4oEHx9GgGO76Bzwa+JD0lrBIM/46bwzkINzuuX1MJOJrh/MSSUnW
DbtuB7qs2NVZmKMSdRKRGXzGE6/5m/kBlCVCJoDmLvxOQa3H+yj30Oo6aUqN/7fW
VdroO60xxyTTd0JaUu7kzeUGWDVgQaT12DE7wAO++McFjy5fkKPXaLW2TilY7M38
MAXuUGYcXgie5keHQrJj5N7RLbEs99ucMNQVtw9aJp06vyNhcmTfjMtYoLCu8DSh
4ZQZtWqTJMZGwTvS/ksyO9JXPjEdKK/r+FKPsUWIEdov5/uR4ZoRAYmXKDksm8M2
esY/IPD/aiVQtZwyMQnq/cQ90tGxUdue6XYgQte7qHPXIfL2H95GdHCQpObRn0eS
zf7TV6tNaoSZEpwCzuD778AKXKMG0LQucrjiAPLbR/r5Wl0p8NEo8tNQeSaIemF3
0bj6c9wa79OMXJp1qUhQOcKVzcA+T4LLkPOqAMhzm7XoxzfpuZ7dE++rTokRcfx6
bfl1k9gKdM9da/+cnmWKtPXROOw+KKI85t/KroC+SdWa7aZS5K6o4W42hF+Y4DjZ
bmHdiH+biooSJDCNWoUqF5dlz9zskIPIDvkzOnqLeVnYbtHOdQ83vXbZleeSHuFD
GH5wGe0U4jRHIFUBAph0FGv/YYMOsL2xTGZPrs+8Yab5/A0I2Mbn0Mwc6+UXWUND
3upBt6orn2jo8XOzNbJZU6tYSXOpTTaw09ZFs8ddjND4wQmnSdj895b/yq+RA4aZ
S6gn4DMze7jBSMhdYvmfWXmdDbhB0aZBTH2X3z9BnyOyGvhqcaeJ6ZkknvWOz9md
usa0wQlSylmEOCmAD1r66hFMBYKIwulJXGSUD37dXN/8ZAAMExavWagqPO4M8Phw
bjf1M1kt59OlOD0ExRmnEN2AJGdy+CrUSkfyMpNVaZSVO6mz14XniW4vhPaCGB8q
7A9sU/xIwfeMguNm2vdHnkfTU5HHbXjBdbhxYPuRnG5ehnbZH29dxHAb1qNtZzcK
+kf2ttHuTVB+9aEp5Y2Iex0DUEVyuKnTFx7wdZmfrNHm34QOb7fDoqAxka8QKRlT
f/Wgasi7McKGJUTcSMBaZkRNL5ece4QpOiYoVRvWlzhg7jaQG4myE5m+NrF7lGn8
YacpOOD61WMyHmbSrqOqq3WCV3ut33wSkSrpbjO6XX13sToxJkiI1XTMs+02SF4a
f46cWS1ISAts1hPaThmH+5Y53BZiurg5NGKNP38WBp4NtYyMtCz6bZFzssRvyOMp
0DL1AaaEbjQYB95FAIpxHJ3p2FyR0d3zP2t7mgSaeVnXSjIxurbbX4XjqXPF31lx
rKhxfwg2GrlohN/9Y/DIIYpSJF652kHoPSqGdaXoifaHeptURfuNPY2r1d2/KJfC
Blg1X2VHGWhfjJOadt0ThyiaKZoQa2gRcYjMTBDNQDwoWJV5ZmeTjOMNCevxYsaG
ShAJ9SlEsciz6Is5z/o3Z41NzLaUxRzJ4aYG5R7wBYvFOb2k2FLGN5RKBe7c5A/M
fYL3WagoobECh17DJ+xbfkVixCp2eaYNXuUetIe/2u+mWuXN0iRI5Uc8fJJIKGe9
xe0m0k4W8qTl08EoXUNMzpfqjIFdwHUmcRhVHptvErbST8vvzglz1J1rb5HJB8ia
cz76V+OWqpZJd43QcU4IxNyP7A64AORnpNVz+dLvlOArHC/y+sAGeolAr2pUX6rV
MOuamzQ0FAsiU+MEkFU76blveftJJBwfJOQx1l4WZ19zDzO2RiSGEkAVasaCj3NV
YIN04RA9ZftDtplSViqKCVB+WmRUChpdFeYW2T71Ft/uB6z39v5AT8shWDdVXKV7
hzfxgG0I0oswSJsYNUA/swKv7puL++Maubsb58/SfkenKBsEbllz4cFHGXUNweBc
iskrnJ1Y/PzQuibyM5nXx7k83hcz9VNNwpVCoqI5xbe0Lm8NHC+jRlmplY427U9d
KRP5sgvmcszBeBND+f8LOpEoHyzk6JoxAEF6+Rp+OZ/bIZLXohFMekho2Btl9vM6
cdSNjpxguW8lJGNujZ7TGMkysYNLpC6MvkIVNuN/ffgw94CrdKM0zGCOfavNm3/W
NUsPboEMy/MSLnAT6fcTK4s4VT6JSOImHfgn1tsvwXykuk/iL2mdR42SmP9l2mdT
wVWQ10VCDAhfYs7v+ZX3/z+lx7+OFGGxnnQOxYMHfelPEUEEq8+fqqF7B4r6z2zQ
TnOI8+8ZAIphumtYp9mF1q9ylDM92PE5qhz6jQ1Txdb8zK5ewczbw4BzaY443Ouj
Tr+ZrEAC4m9WmrWzoWmk/aFta1C6nprWgK8vVernWKW7Gm8wP7gkbniRNr4d4cIl
bjVqDizd5SvouFfdXgrQujw4cnf5BFxQM65dCxYpkhNlhRtcyBUvjLHQjuahHbr/
89vj0HW899K2VwkZLkMFEPEw6ILsi+TXE9XRZtL3Z0jP0lvKlTc3ioRNGanLDHM6
ezL+Mmeod9Bs3sQERI3C5vX2qo1h+5xxYnJAQt8QqCvr2bkjzVh7kLejXD8GQwM4
y9zMgjU9+BtRib33Qn2/kRIX/0rrHxsLeSfYowNeXDHcWyeYF0vvRbedtS/PHtqI
XDG4dCXA8dklBGGttf8OMopDL2erVk811gKV976B7l9oGx7FyecKSdP1cHZy6C+e
sKvaeKi3OQPKYpd8YJd4L3kdyDPXH59+9wv6dLKDA+CMA3msCGULVgTAHWaps408
EDvTbWErBK2jqvQN275vdTpe3Ce9RbyS89qs54oLln55O0UwVg9xLAkeUUoeG5/s
q43hL56d3Pt3ZbbT3hvvVmUie8igbLrr7DbBs41Gs0cHG3NIvV4IbNv0eoPlz06M
7H59k4exUdnwswH7Qv1fTBLvCEb+JuaIDLwb1ZeV6/bv8nM7qPP+aSOzV9F/lGMs
LmSosoSRaIxZ4nZcpW5pHzJFe/O/l0836orQ3JgQKKacRB3elgQcw+3VQ92E8LkE
PRKBoi7bKXQYV0dwxTa4aYwHLj7LfrAr7MAFZGMxKlNpa5JLtEnWOscyqNON+AH5
kTS2N3fzkRBnGNlwBqYBxdHH7ilnWyXshT2gtIE41IR1XNNwH06dZK/KRudxVAV0
CSQTc+XEGWUIEdONqnONi//A+MkUPVuaqmqBWNUhqqh4tqjRH7rM/bd7ssLIZ2Um
+ihHzrGILPG91Nubc5fxYGxf+xEgFduxQa6TQHoImG4qKa4yDXRsQB4Y2Dttia4M
b8y18xPsdIk8KHxYAy8K35VQUWhnYYctEnO+wQGxdkWxXFP5reUEgDB3hc7VcgUE
y1EjN7a0WgF58byaAqy4xmLSD2GSV5Mc413KzGD1AEJUeSrBXMlJusXiYDyQJMxl
cadSCV/oVKjLJMRR++UG9+JRj+H26N3zfLk9ba9ZcmtIgV0CPO+oFUmT2pCOJMwZ
SaF8K2/5bU8ko1uvdNHMpNwBxGEfNBHw9ySVhFg+iirxSs3NVmJWbyiWo+xYRzA2
gqPCyJQz/oG0Ns5AjwVJoZn+WfR6eu3o/bQua4NIIup1Zzrhx8Luhz11IE+S+yrE
embhgyXBdNOn1BWpxpB576vJmTprxQLyG3ye4QAxaXq79xWjztuGj/5YJuwof1Vn
ZAhMIBDUaAyNZ3Bu0ffpitDWzinFiZ3oji9kTdHqYXHUr2hrpjS76WfJ2U6dTGS1
Gdiy+haIfm6CmmT/xnpuWMReioSHzrUuW2QXSow8OIve90R+U+H0914sPG6mtrHW
AFVnZVRUbWg/HiNTesbe33vJ/KJFQxLy6Ob9KsFJQJ1RjI89ohMD7lNnHLUJgAbg
ZCZOKIlOVhlzIn8fltUUxt/09/vjVmWlUf/sQ9GDOCSINxQ/sbQ/F2534/DPLC/5
JKf1y5M6kbndD3SPbT3cwHUuwoZRx4kHxhNMALviWUhnJimnSD9pyDRd07c4hoB6
cvrPuKkg6Pk4xJGsdtZaWf9WNsiNTueGtkTgskNOPd10eFmQboiaT1cemo7RgrRc
go95sWYN1jIZrYU1vpLTWAOU6lwjpduCdaktqQh6eeSwYGsk0arYEO/Na+EhuPew
QYIDo7170EhciywEw1nJWOBLKlT+3TrgZrNMIU4Xx+bzoCs/DjkU4jRsdA4t7GFd
i4fdHT6ZUfi1XFg3tN1E/q4Y4LEDOJ0pRB/b1oMKHVarZcegA4EB4Dq1vg6DXZM0
MeCuUjEaiwHRQ1L150uWSaiQS+frIsMbS3yLQochVdxecvIuc1tY+rE1ihuEXGXa
+Kc3D+ySZeBW3nGGFMn2qtF/mxc9o9WR09EdR39F2nXhjbrSIJWu633PTxBZ6iFA
0d/+1bsSLHz947Biczv88Y3qoB4D5CEBtfnfbOdBxtvosg8XhhwpVHnOvWkL40ld
FbvaMLHY9uI6aq2372HuIRujAqO5ohj/UAn9bmUz2xJu6IPzNz6/zGeHCFoBkPBF
8FN9XvGumand5FYNLXlJSGSaOv6K4ah1SX0zmEIrCfZYjPr+YvJSitcaQlJf+SqM
vwAIKFF60vAko6MgF2X/3Fwrj0nLdy0mr+GngWol0yCs3chsTEXtjqaPy9OGF202
Ws+I/VQwzyuHhRMszU13EO9aR27QYOcxPPrrvcYsBfWT1zPR81Ut3DWWr/jPOFEd
VIlWjsfE14W3RscdcxLpm4NGXUAvxJWBgOQNBY3HNSxwOiUT1TttVAJVVEWhCA2M
F6laUt4T5aBr4hCzLQcEml7Rno5tRI5FceIbHp6qpPpPyOMm2ZYMw77DEhg6h7GN
5Wfm6/JAJlkiRuwX98e6koN6CwVZSDc91On+cAnrXJK5GFGRVfjgbLL/b/F+7w64
cFsG7sD6aXFQHYA82KjN576HbB5rB5dEalOlgG9bNIGhHvEjeZ5qJV7Wp2f2hDNx
VrF7iuNlHXKcanaJ2NIuAfpKL1eaj9YQGVXFjcuiNatvGc7GRhxtS6cm8fFC6ipl
Aa8x6TZ8AzTYYzhQjhu/G0LoZ1eDkVnQFz0i0XENyxYEMYyIb3+8jASIuqjrP3d5
BhE8Y8CXoAXul6+7cogqCMN0AeEq9FaHj94QRerv9tU6FifDe6nMwexyP+343wN1
Q4RdKj3wAK9z8FBcowmVjFn4ONF29lE+rsxiijLYRrY2a9T9PO2v0GSXjPgUkzOn
iexz8ei9sPMuorpQDtCQ0SihMBdh6xMVlM5nQ9CYflOElkUvSxjcLCIdSfgCKJuw
khoE0WUKHiw9g5a8105W7aXiXUcQUOJnG+JvJCN9Hy9hE0BYaBcqf3Jk/MEKK6xA
ufwZlnui87h++wWpWY8kf4gIELZ36dPUAoDi7GX5znsWFP9HzDervyP7qx4YXUvu
X1xLFhIY7TfGmoA5zE6Y2+YM4XcwQ9kLNB7/LAj/0vnlxGjBtX7yvKHnXEoQatQe
XZgBI857MFhJ4yOevW4c+Xb3jwGk+91lmi7GE7TustYLmsApz18ttf1Fz7y+4dLM
X02I78ONLeThIhH5/aXFhApBK9d1bv5gjk1692rIfpRyIDixaM2XjKJjqzodkhzZ
kywn/qU+FJxcjsWd9sZNvgQi/SywUM/nkklEKozvJ8p3sKN1EV3MlloElQUvH2kM
c32y/UXU/2xBv4PMCULIfP94//HRugH95VbfREbsABuku9ZlGkeMXMgJdxnYywF/
UIpevxivLXJvIDprpBxDwQTbNs+1Ig6GCxohXzWlMC5aArRCXDpyZZ4oT+Rtpod6
I66Y+ExbwhJpA9ettRv/et2OjM5F3Zs3Z23JYXSGzVqQww81R2leBcM451ifFUaU
DC4myd/C8BttFv5xfqEqHdA84GejOExxgPLecHgXHW1u5RWfKmtrtmy31BfdOQ5a
jTj26eF3JXYgOUmhDTUdc+CfrYe8DNaq6CAK9Wlqca8O2Eple3B51HWah/Gng1bF
8pdv55QMBr34gEp5VhTcgDbpRSc/TsbBn9vXzwPucoYavknEFj39pc5+rTHqsu6i
KDAZyEQacCWDE4ifpOWao7MoLJ4LRQxT5f2jzzR+oMg7RpYBJH3s2tQQ/QyIWE6J
qD3BaN7wPMnQ4ptxFSoNih2xkbZnsIhavdtaZUI45iqV4uOTvqnQ1u+j0SDzRD6a
oc0vPnVzjTzxuigXySgcZoSBvlM7QOxmUSAQ0fdMvOVQ3XShHvJwYNhL3AUdbE6/
WYqoG3G6hVgPR74W05FTTZ2lDLWlwbxHFUT8LcKlljwW8vEmlnc0Q0mrnelh8bzt
l/l9Ls3N8ZHN4+jHPuBcu/D6NCrt2qn3PM5Esl0OEw6NPthlki7jsmO4zsmlMx6s
Sm0c4crxQphspJVCF7n3CtBdM/OvgNmrQV0mlKJfR6nX/E2lyVZaBJoko+hyYIch
ngRyY++lVuZ0AtWDSg7xzHpfLe5S+yH11y2Tqu36D3cQdVmUN4Ixd1mDfLq75W7T
hGG187LuPqQYBEEj2qUgad6VziMWaCeEiHxtu6vdy0N2G0L35N7mAJjjvgl2LnJ+
G2aps2+bsEPnML/VZlY/e3OI4+Yj6UT+SSBy4ko6MeN0LL6Bem02ncnxALGCgXEO
8HMgoScS4OzOyZwgfDq9JPDnSae9k45MrOJJq3PQBHOamDAX7D7WVV8xL8AHz8FP
5E9cRv+dU8gX9w2kvYg4zXWtnjSeSm+eKqe4NMBZv99DgiE1Lo5JMvUgFOdVJlUE
VNNQkTdcKWxEkJPM9ZE83Vur6ubc5Y73CfVKUvZvVuGvGBPx3t/6ah7+KTwIl0HJ
DQ4dCHmua+KqInieBXhaVl9IMxLLiJW8rf4Pc5k60hzTE4+oOUB/cOw5V45zVBET
7Y3Ko5rX8mrYkttjxRJ4VDx0PSYFOacjiS+SI+tLJjblf/04BVINb2w6rB8nudTP
7Wm077whExYBSGIiV/2wyOCSWfx6uWHM5T/L5ErtUoe/2apNciVc/OjrtW2CIDsz
uM4LVifq/B/DNFarXaajsf5ASCdB0dCrs85gAzkVg6kqIVZWwm1XXxl+CJ3D9yWa
s1gQhQpkg2Gw5TOFDzY9/UFgv4JCVCbG0TA2ywyntONqHBFWyEfDZXr5EsR/h7ic
+E3BAPNxJDZLI2wvgyEvxrb0C44q6wz9u6EgmBVsk6qfQpm7wHvVYxI/c/jCz+Zf
pal05qU9gkv2lJ+Pt7w47Y4OjOlEGboHiOvHv+UVj8dbeeaT0Y0Jd8fFGhcGI7TR
gQo7XsoRFDXQr0srsYG8cEV2/Jmbs9xDtwJ4yMNqii+ARa5ajugQ4rswOHCDzkDD
Rijna8mtvIwJDD06RlF8WV2sEUFC8v+N+nPnjonqMQEmcAj4uHMKT9JkPmaVbmsg
LOdRJf1koM7MqKUJv2PIjU8jB7vqxGuKlY7NbM7gn4KwSt+WjYIEMDWA478WUTeK
EAnKsDKerYS9oWy9VfutZv6igh9IkS03trt8T5UzQubbfWP1EeYXk5GBw/bRGzJl
0Li6a1gd5aEWQz0CZp5IA8voJM0Xu5Z0EcFFABFu1u3i212dD/kl5fuGvnP6T+vy
o8GrG4xIWigjk8YGYXmPmKHZn6DMA7Tq8A52oDK2yQxh0k6yNZcSWdfwdxPfsv+s
ZONXrvoMlIhgxBcJw9tG2fYMePrdlwdAChOujTyw5qzhYBVZ9i0XlCV7epFuP868
AYZHBgyalh4IwSpwZF2QSwtcq1XlQ6UrBHF72klncYZ+Leci8Otpw0Y6i+HaDWSz
1hM+PgEKN7D6VehhK9VfJBdchJQKyyoSYnWLcpQhDKtB3JVnJYLVPPqkjdHKOGX8
NGNI4vlmiazw6LNVPARyoIeg/pc8Jz4qLQ5PGObMiTHxTjArEgaGMLFgWXCkN6dR
tcJpXwYEmB/DMu+2zhXONGIp/YEyxKHGmIlc8Th2UY1kBz6FhP3W0u+7ugM60/Kr
etOffY+BUT386MRyvPgy4QrTDb57Im9YebmhOs6eT5QvqRlCEHApL5vkI/1GfTxh
9kheHVkiJSv6BRdiRI0mwFpURdkc8a2CWwW1Nd4zwhkHVqZXYNZVF8MNmA702oA9
3Rw+myGD4mzy9hSry9khTbdb2a3IB68+3VtQtbY7AbiV7/WWYLIGtH4hfEYDMN+r
YI4wN44XZPFCxCjkkz9SGjuPGo/iD4HBQ2+dZfTmq7SGNxbArxvWbi//iNbqm93v
WhIjXtjOeIDrm8Dduc95zWNuZOA9RaJhv/SJev/47+Bd2hhyQoAa0tSbemKZ3VOc
zZVRccIo8JLMwnEUoZ7HsSe4eHbmAOXMW5oic2V44DO2ZzISZA/psYVvDpt8Yhmy
K59aHoq/mZgi+KjQ1OXIgTR9ARrPBb6DxWzcjm/Zs8J+LX4cEGOowI9bWk6lEbFn
y/czn08DJpEEmCa0SPon5sVJdmksXSSTP5JzRLueNr2FIcScZm7ymMt9ktANH96u
JfV6Btdbc8uve+S7Ez1mNQWyYjURGPa1yk+Zi+TtV9f3sl0E+pdBj2+mTwda/Yjo
PwbsxTTM1nI8OS5cudbl3Jtq1r8SI7gYFmWR6F9ub996pnUAb0x/ldqThNuxfuhs
erw49d9S+YyBHCcvQnyLBoGte/VvqkaapxQN2VtAyo1pWpW9+SeI1MGqJgiHf5vw
JoGeLxnhKnq8jahtj6cUd06h0AUMMWaZAvsUCdq5QiXzoPk6hmFJ/MerFztm4lGv
GZIDz4xgONZ+9nyge4ZLEGBj8KmACT4jK2ToDmtEkgeBS0wRxuGJ6weuMj2dNnkJ
YtZHg90wCZxwKUbG42CrRR22aJm3RsT3MpEz9KHkUT1BsuIeiWLyagIQGTZBLKHE
TQI3Y3fk7BVduTYFW+3HGUDgdwOGlzqoznfka5824qDDA/e8LrmNiVVEP5K2t0AH
b7CLWy6zhj4L90pBi8MhgBLUJd/m+6EP5FQAvLUHfmXd5CRLUIZCiwu4NZiVrpPI
/MGakdpIseQZWA+c+zlnFbbTRkfMkm2xlQbaVv+64PQuv5/aIv+iMUvbbLQSebOS
3B7Dd4pmqujyP1PfPBONdvtr65VCa9bVQVstr70Lwfs7QhxYOzJjiyvjBw0UAFay
m0xxXUA368/x0FAIG0OXl+/2NJwdYTfhRzqNfQr0LhGpwqaL1af1YP3r0lr1LF6F
8YvNoPsKOwHgICClrNyEDkgZCIClAcxZ3v+ViDa9uVUxNu20FuZZFroy90sxOg6S
AK3lmcQxqt6EpwxLwanNKE1S8F06hcR3ZErXsiD8j4Jsqymb+cqz0+hKlRXmnVF0
gMoqMCK26EJ1ADB+s3gaPxmTTN5BJrc9N4v3qpL8wgydaITpkXrWqqb/fu+mcKD3
9BOgIG7VUsGGsGs1X4KfyTvTanNRcSj1l+ZuMSFXAh/J0D8ZzCFHNsQY1opZ50f/
THGKukDEW4f4CCOnvRwsUpLLAIh0DjWvO4I5r22LmHPLlHau0IqccOGGe8TYtG6S
nG7HfJlf8R2qHt8LkThfw8uVkM3rogqiUkwN01G/gyOcMwW5DB6gZpRhDPZkvkYL
oL7p+W9GxiMmLhI/gAf1bvBJXnftiysqhMGgpGHozhR/7dyRP3RzM0cCsLojdbnw
U/m4+/8jUO6y1AkaV1flf50we7KQxr8yo+YTCwJroE50jOgyDKukSL5d6p9iSFt3
dLl51g+o/EEKdjsIY+Sf9nlK1wzhgARhcEmn1ET3MmiUWQZVYFkT9Ks91JZ63Btm
oz19/vE4dKyWJo4l9zXMMv4dzOFNZt1mX9lwfUcjqiONes4/otczMAVkEN4kz5nQ
ZJBbhkYajBkw1nz0q/hf1j7qJFqECfZSpbLaq8CYk7XHcHe/S6EMPtd/HMN2hsdu
lHSjVwotWTy4jp9u4IA4BEvvd8BEimP+e3FOvvwiVx5Ip75J23IH0I+A0cxesvnW
3DH/VXzvqDY0Yxf690xMDkamo+8APKmkuQ0L9Wae2zm+K2bcvQFjnSFaqTERsWax
aSAr9tA1bWJdr+BKfbb6Ri20Wm+Xfz6lQRFMSYEhQOAI8l7llsMZdUJe/DPc6it1
WRN++6KegK2EpHSppvTCLsCE4ozWZrK6ETrFfm8FJ7y+u0cNkjcEqyK35Hsuv/QK
vtMGEQHKUD8AjkeTIIbbQCitqkJ/yNTzpsPPxS34ldCXxMM5+k8utjVWPg0OW+pG
etGx39Ni8mCwfuyLBjDBUCcfERj2R/8ldl57wxEqosc5IJYmBEgrsgnTyF6UdlXZ
gTr2bARbOqY1UaLsdzF+CCIotrNzNjoACnQLjkWLf1ou9rYH1mgXkd25Mwc+MiJv
B600ZmnSKWzsAPkAYf3iMpFL5VkttzbiXbKuhNCyzSuMi6YW9huK0MwEUFf7JKRa
iBWqQSfvJmM37CypfECugImDFcmxLXk0NS/U4NBhw5sK9HWjdIeB9khnxU8bpmWU
PuFghLVe+R3VemOmeqEJ+4OO98XDA2aOq93FdLpmx8aWt/3cVPQEeA7ulEHjPM2W
QYm8ekrfC78fCVw8wdzKNjftJHplCz1S3TIgGp3/z1LN98Ai09kNMEsUXG6NvgJk
a6AC4JfUBuWW7b9NS7klXTUIEOnVkj5ZcTesB512GpUIBjM+7sT7G9/wbBO0AVq0
sTQThKX2bNhCj+YhmBVQJGyijiF3VSn5JBtj8y6E9zMCI5sWkmdbcvYYuUhPWr3o
Z3vu99j78Q8xJTDEk2qBSFOkQg2FD683YanST+Qdr/yhAfikEg+XFZNjRtG/Nh1B
tQApNURfNPmAKrmvzK6YKIiOpA0Qc7QG4/mtQzIG6+vg8hwKThHPtgV0lgsbOpj9
NvBhpeAoOOuVhbLqqkfl8u1cXuy3L/XvMYpNcRR75BTJSA58nCpz6+4vrhRXnSwy
AHi9/ZEt6tzPD58t4v85pg09hnGs3iZJfhmTVb6LytNYRMQEYgpYeLi5F9Hdms2a
IkoCFP2K6irJEE+AOlgEs1dYOx8hNN1pcwe06+xWGdVycrYxKwNgJMHYghKlkxdM
d/WZt1nMiLV03JzzqlENiSHF3C9tmmq1KlVS5pBr+9i4vtQFrv/pYZ+iv1eDwP0E
u23MnsLzvFF4hpndpB3WOh7bzL9uiKQdB2AXYEu1/vcji8YCNuGblTT2J1SLtM/U
dngsw9V2jx5wy/YWrazWE4EJTMnX6ZJ0xPnJhSasgtR3sz1BDRsSam6FRwN9o8o/
Mgk0ThJKTlSeassqE4DuxxOVKgsWMbZEi8+3lm8CFZE0cRw3FYHr8lE4yNHBLMoS
jdSfPCE71E03iTBrBf0u1jVNGWi1Ejf/4drW8tHnzd62+X9BA+KMN+zGe7eQ5baP
LkOa0VbahvcqQdX1iwnISYrIP9FhOboc/m/6pPTiN+gwAx4bAjr4V20VTU672urQ
Pm1EZhAvgdps0DdsPkNndDEM8IraG4wIhiMNKB1sVRvN49tNsgVVpxFM7sT3zIeA
tQTe+NwiaKNlNmWnXvh3IdSeXsTohJ7DN8gW/YdQyN0ApeGSxUsq0KDWEYQhP4pQ
ZdiKnVv5GrvWEa0gYpfytGPrd3JNSSaBOlnamMF2naatyFtdkZS3pVvhJrd0sLWD
+HGiN7zZcyo2YhMJKwuV1bBo9vy+ut7X2tl65CQphSWq869zlrxom3hzUnMO4afl
qU0Ezt1WnbBx80qeEV01Hof8vGTiJFIrP2FNgQ2Nia31SlSwsDkLduqoDv9x+ysI
vnGmE3gltbEuIS+3COl9ZNGLB1eCzM6W7nMvAnOZW/3O7LYCAQin82TuYiJb1gw2
0it1HQmPSrUlj5U/jNgbM7Uj1sOUo0sUnWLD3yGrdmDDl7EgJ1IAKVKzZJfavqwl
1f8Ms8G44bBVZsdn54CL4VTR3d/O6gmXG5m63qzJjvTi28XDmvbfMLLbHYXU5oUc
dJgFJePBzdNexlgNOMd0vqExvtfkSegFlJhvr9GeOZA4PgWK+AhyFyy/TXZd8Kn3
h8xKflMaPJg3Y0T9ZOAmH9qDe7ELfeVu2zT2JDqmD9v0WBwtGXRlaSOgDS4AomD7
cCKn09GOwD8mTG4tk0xixP2xeaOqRbvL66QaA7iN38LXB7+vkoDl88jDGkg9sgRp
TrdRUQVyrCDi7UWc6PNUBnrY5aI+SGek7wTh/ClMSt+Ln5PUQB5q5xIzDgx3nVd3
xtEYZYndV9w8aDgzua9VcjRz+gSOxFUzCwTaAFIfBXFs4kF0F51Wwd1cws/IBDuo
7W+uPEKKVteISYOUZ28gLZ0qCfInVPAFJBw0zf/nXMDy7DGmGXkQHf+s+Df0BgvA
mXySSLOTqbinSng6s4lzbedA+AH3d+MbcTtFISidKFy0uN+c7YCT8EyZuYJh5qha
JrJhkoyTvnPAIbSv0+v1tNKiEs5U7TQDK7hu0l0fRr6WFVT4ZQlHYa2FrALHzbWw
E3U+kWjPYRkm3usm+vK2AqdC6dGEk51XX9rLii+NeSo/u27glr7OwSsQjt0dnOgG
eCFdaaEUsAI6fYHrBeQM3+ooOY1Nuj+YIvrmww7443FLiZOsUWlGXaMgQrzPsOzB
pBgd+jJrrVdn0pgGN6P94eodIOhlxFZ37wFoabHiMrHafwD+OBeDseroD410wApL
PHSDbGetTY3BRDoY/UPCBb/S/Zpdkl/VwXpWhPpgTVi31Wu+Ky3khZsWc6QT24vK
470wKV1/Q9oigpQp8Qm1GFYIDoBDC15OjYQXWPBiIhulOXpkbzFkqYHQvHqvoLOu
E2Vl+fSZhwSsXcKeZnTiB8bzgGAE+6eyQMsAU4iPdSei4U82DqBL3exohbjmnnAQ
qsTqNi4izBBphnb2Wr19e5H7f1bndMeIrB6+0Y6/IiBVNsMXOKJQUBN1AL5BfOcW
ajIGT5t5hxLWlzOpFbFdrZIV5rkOXThCQ2E0HeR+D82jR8M0OvRT03R40kGWLKsX
t2MUKIeLvtHrc534gVAZ8ki44PDXtehU8BinyRq2p1e2/JUNIZdIdot4j6za6Ndf
VrslW8alzk3WJjA3FdZi454kOcod/yMj8iu5t6t29syGAjbGzLoWcRGoM1blQFIA
xsB2d9WeXZXLNNrUBEU5iZVjsgMHRnSt+MCJYRcan3daIqydHna49B1eMN4ZWlMY
eBEwb6yUpQ/0tpGGkp+QHro57o3PQB7RPxX8f8lcxvDsDEx9vcYXOrW4iNy8Arlo
lOyMq2uCNuNT5ylocs407qzEBlKbQ+Pdxe3zF52c49brVZlwyTktUnYwJQ3zNXQs
pau9GQ+HNH5c4QIAHs5ddJLuRbKVammjB37uF8PiQ3Xa+suetumrBbeD03HKQFpH
5Y4mYv4jU7UWhDkQSjvWrQwC0fPgGXBodvTxKPVOLt4TDea0+qDH/QtHss0N7NsH
ygvI6tt8q/9vcG3BhPadhqOb5ExxLIJU2tZECmj2Ygs+fgIslQoIKkOFmd6yVbAe
XpSpGUaTH/zcYHGdlVQNxZXsXms4wwcW97o6T5lx/Xqj8t0gYEnE+vq6jC51LObH
iHbEHqQ8mdOAhzgbyNix1CvEkxyeIJ9ESW65SE2T2ntZXM/Ch92Whp9i7M61CSOh
peAZiRib8mpllr01ZkNb64kpuveijcrFtpkCaeAKInQVdx7WH/SzAZ/29EZpihdv
/QrH+NnVg2G3epY6LsYk6a5YIbYnJ3nIK3dwp33MZl4en5YhFzcRwhaM6qpK385w
5hzVFLHWK33Bx0IVDCaqOOHIXB0ilZNa0ljJVCHn8Q2rejL/BeBeIWwep/XlTlcM
sz8PNZ9tEj5OxWpL+II1Ns/huOimy/Q54r2nDM2cB8WCiDCXztl1aXrXHzEESFOw
F7y+UB5zH0EUqzH824d+fTQ2WXebXzWINFOlw5tFBsQW5Ma4JBhafkrFFgrOWI4w
AAJ0yzZqx6yrb1v62KNWLw5aFWLnRV5ZqaA+HtGjw3guUQqV/ngQLzCdevn4/evG
p1k8gmta0vgvu0n43ZFJax16MeHKI3+rVf1z1RmBspZoG3VtiXkphT0RqpC1evL/
xNAtySPeuYMFjEPNy4WSuDA7SMBfT+TZLn3QvNBUxbL9gAFsnLDIpd6AfBBfMKM8
riZ+IxAYj3nR2XxDjcw84ZnEwUOxfN9J1hmnC6xh9cds1gG5PMGipGM4Wr2zb4tf
6QVIdOWt1iSlRq+t5bqU/lxw12A8v0KrCy4Zc6Hl88j4rPsOBZAifGWhBegHIZL0
D+gLRwW7O8XhjuKQibw3IvHeeJtz7ZIizURl2npoUm7aZC9RSOXz2zrpnDCd2a77
x5xXzRBZLX5gbyniPYinq2mnrF9QTbdg/dhNtMwzXSFsdoimt8IHnsYVm5UkCIGM
KRTq4UQql3Z8ZGLexw8Wegk5TZEGMZxSe9f6c2Ah0KcAApbxfRbDU+9C8mxHHiQ9
uoCV1ux0YEwvs9Bo03oFgOPbSJy6OXujluIHnbv1XpcoaYqt4OsRbscpqqtuRL/C
Oi1D3LeRCWbLg1Rurx3QCVrzbb9rQe8bjy7N9YXuygr5euB/A/aLm24FhlOrKq3C
pE5KEfjpPpA6YSbl7EQgRfXc3DZMSkEBxCZWc13qWYJXBnvsQ20EewlXNq3bbgSN
yn4oxvH/Cs9XV9r9IoI8A9RZDmT+e61u99eQCe0cSteFeH0xv7MDWoQKqMzwoXAm
nCMjs4aABYH15qotlANy1tqcNGunz+0pYtW5Cua2ZPJ2C5UOcB6QGeVAcNwAojnW
ozeErHjsIsW3d9RtbBmXtrQtogOnxRTFmEUUgzDt8IW1HX56qfcZ3UkWMMyHFb2L
dB6VPAAOXE5qExZnoLKohqwSC2ZYzlhaDzx0mBnprl/gktlXGRIUl4ei4c4opXFy
WdjJs3dp2pTpEkxRkQXy2NFJDQkmabqL1PUfepdbIefc1qdmoX5L8xhy7s8eGiEg
xUVc9TiliUTLCXXUS0dTYvXEjp9S4Ycb4O1vUbizZQKBX6uLAdXjvgrk/+vFOM8j
lBtmfhLiJAmfkNcbWZU0b3arGR44u8Uf05yp9kkDRf6wUeI9Unf4++IrMbqUFb/6
qUn1e8wYk84nArJH8KjrAQM3dQ3o61y/tQBebQs1NyD22cwEOBZZI14W6U5vwiTI
Sv8rhJ+cgb3SGFOl5OJ99PAyLoCUk4hi0WcGeaSh6zFLTQHo3C7sHGsEaqUWpBVa
K265npsn5CAKUlX/kxNRZxzrpQkHsZDOlxAgBxat/Ka/B0HeNekBJpcOzFIkUQ1N
MmibGchOy7Ija4o4jTOA0X24sk79pzxteQK74urJfw9zi4+uBmWvHG7YRRGIdG56
0NCATHgwClCAxIndiwagXKdjG5Npb1r5fYt6b7Vkoer4wdv/hVpYfPrirQABu+UM
aFqGob34Lg4Vf3PiRJc+wdMoQtMBf/yZWqz+kzYwextpPkq/jhMUTmi/MSC8TroJ
+2rXXhLwEy5ybiPNxemfGRCOcWUefvkQPKxhp91C9kx00iaTocrZ8LGpfcHBo830
+3QBE+d5MuPAc4yK74roeg5HBTNnS1QZ2/g29NzUpSTPN0O9nxac7pVanabTcloS
Rtu8LjEFETvu9wlY4QKRnPPZ+4rlg7T8UfAfUGgKZGVjww0ux5mOpUgt2RzvphFw
CRVKzufN+XmFWbNzqmvPhAEn3G+QfdWGX1inKf8cHwkKqUbU2GFcs9hrcy2XRprn
Qp24o5hYqUqqXh0TQAW7Pqjw6BoDoBRcCExrAYJ78jRrxTVkIygRbZeu7rosPiDy
MNDPaPy3GrqtFW0i0jUut7oqZ5FdL6//s/to9SBZeq8wW7Sxlu3RQ4LWBC4fSnUB
qoTKYHOJp5dIenipOh8MydEYn/y/cT28IEeu62KSTJ/dlnd7eACmjwyPm+x4O+6W
CsdR9v71hlHCdEVqykSeMIG256P4dyGLCfkv5acYN2LtMU1EN44Klm7J0bV+ipe+
VvTuW+fWhV+mbnpFn2701t5HMFgdXe9AS68ESYRqr5NlPXauUAj9iRqJBmMJsZnx
v4cGnUzIClqU1+cGEydi5rIKOCCip5npRg62cAK2udpF/WzJFZ5roGs3Ny/itT10
ZXe9qrnGq4yYk1AbWarjKUeuGt2MMVDwszrSqutXLXqpKc7kgi7FzJo9+2q0Gikf
lsmXxmLgOF5Wg8LZe8+oWANP75z1+HkrFyI+tNyltnDOuc9QOE69Qmy09re3YD09
KBtISIUG/IHykbbCSHJa8izWN8XB7MiGbNt8dTvr7KBClM2GeXy8xgDV/4dxTfCD
uLKEhI91z0u5okBtUuNjQwQbm6QONSs9Q0PpWUvBo14pm4NDL2TQ61vJC2kY4NmL
N2kYlIJdzu/jf+5MjIzHIwnVVctxySyAUgMGiBeTaFfHAKfvgywRYWHZ4apuwH2D
mmqT/ihM+XrCEIVnVVJSvpmWWnb8EJkcPhhVX/MD5tqAadnkldupTypzE3sSeArd
oRHEOfPW98oHci/C32CydZ/Ie5+L1jLDPro1uVOR13CZFPiUe0cBHVk6x6c5YNow
1ggfH58HbW1JU4R754sU5xw2IwIJTUen9SoeA2vIjEkGOrYCYJwEZqvQjKVEwQjt
t5edDZJ5FLdr/AY378syD67q5xZzt3kVTDb+xSanYCliIvU7ftVZvvQI2jPXoZ27
Qc30tlRKdyVkgJzHAAO4I8zbH8xp5FIZc88RCMzQvYJNjB18qMpK4YWRL/Otjt1d
Eed9kiY4nxSO+e7y3FLjmDiro4MWxFmqBJExKFiN0GBvvLH0DkOwTWE6l2Jijb2D
LhhyZusGIV5X8iYVjV9krTYDCgT9zForSAJcs16Bz+uXH+tTFx6ttUXlgEUp0DHd
3K/2QSKFAKzwcSk5aKf0Yv3a3H8a/ewEnVziXBd9Y80v1X6ioij9NlXvF49atRdD
lLnNizvOWmzUEGF08NZKt3C/b+5O4a6cpPKXNHQrRN2gmhbnglsEKMKmAZRj8gpH
g7agdiV36n2B/nc9EcDx53A+ZcpdJ0PR+0tztXsV9QRAp7IO3Abotp25BfndETSx
kUEZNpxaOpzzlud6C4Qk8zsghp/GBjnxcJvE/JMsYH963+rVKoBkpXZEa6cDBUGz
NcGltvWzTNXbzeWXGlY57BgAkY5O6NNFzKYP3+n7s4BXXsDo+IUBzSXKjm4THhwr
I9s1h3rIyz3xWcDjITU86TkYRPL/zJQ87+5Ott7ca1l1pSbtDYoaOUAqZs1PFKtd
tScuZDBeX+IFa19yAVFJqOylmWvJLJrTg4VHnZ8uk56WYLnzHtXAaau+2FFd1X6s
Jb24hQ+RAmCCZGhVuQE1+Dy3pPJPGBUDtuCTvdMOrUR3twKhSbhMd3sT4bXBU8OJ
XvrnIThUYXaeSBH7mOphsLcAQGSNNGBEetrnC7LkJ7c23glbHdG6HzwWFQblEyra
7m5NrOe1TX5SpU7P6QG0zWiK0MAat2u846jkcs2AeEGfKiV2nQyfHMunyIgZqMsy
biizVMYNWtMX2F14lcmsHVYpGR/7udPvmuoHVJroE0Girn46tbn9dhJ/jmWR098c
8/9PjJ4pXtsJdM6Doz/QxcUkJdjKyRzH5tOWfhp5tMW2WLtYdvbq48LXiABrHWHk
jHGZoEejVMc9E4F4X6U9sTIMXMCtzHYeTyIiKY3fqjhZfSMaQID+ZMAv798J61Z3
bllrgFpu6DgbIIJAeKdNHDn1KoUkBIWwgdlfkKXVAgMWb6G8pvy9hKB8lbvWGELe
oYIurpU4UlJ+ndPFBZTbXGs5mHTrvXVe9uYksUauxMGO1H7SAiqPNJ1/iOUHfiwF
J0KnqsdQog/2+urkdveIJBQDA7/N4Rrjq4V+IY553C9v+tHhThKviKhk+aHe8/zK
45rq862yy5YE3qfC1/AFB4vT2kit3HVeMfn9BNsR0/IeszpqzfggN6H3CKbld1aI
5PVmW0ftbH1gq+yofXgGjU84ctmsrXt42sGMtEzkU+3t3YIqQ4oGIsVvZ4zLxgEC
T539Z2JMNjSZpiTrbHctXQ1ImFVo/PjGL7JStYQYMQnMmH4WT1AF8EZvNgGcKBYl
J1kJ3XZ2RCnWMD0VYrAmsvGtAABYwTa8VoJbWZcM5iLAC0/ONVyF8ohkwI1Mtyld
GI2BvkrIYhdv74DkWqRrHuWcgcFoOV3/DC20kxUKvHOGnb3wvG07NZG3O7ZV0BLw
nDgNW7HEkzg2m85x5VPTvQs53daf8O9+G3VzbUXK8W/h6KLl4hIoD4PzGPqcgbf0
e37AixAMyT+CpGtO9tPfetEQ2+mbLGXrLbxIPwYyHvccX0TQbL2PSWDhVTDN+bXT
974z2KYpunr7pp6aGt2N3CpybXA89k/7at1Yxdm53wiNIWc86tmUe7hSIG6OezbK
FpOJpPLzKDgLYA1OndtxuQrBx6TyRTA0FUvjGcin39MK6VzA7AjRORQyDD4aaDhR
qT4M07WUZlUEzsLvZBf+/Lq/w9ORCAc76diQ6nQJuCAJ9BrkR2im8TqREbACTk/T
FVTP7zZFvVIePmggXEFRg1XMxeqZ6yYvWGep78lSvYSB3Vpy4OabOkjL+pPEP0OK
t4pLyG2SRj19MdK2rdoGs4rw7nbimGkrmQ9AgfVWkZfV2G1zRkqDIQ48W6kbBhiL
YK/2fzcd30MriU4acNqNlN5ZaCtunE2f2kDUJtD/mIV9HJ6MuJ/znJj1aw0tJzoy
xSEHGmbTY4z057qt1/04fFanWoXs5YXBQe/QRZoxDG/g/hpXLCk3qLyBx1aoesbC
8bdeJj6m1Ot0t6b6rVCKFo+W5e7t2uP+N7Hrbk5xwo8/oknU24OsHLaZDcmGkLt/
+FFXDQmJe5RGTV3bDvBd1tNJi/KLY/UA0X+sJxGIzAJURFH3FAYmt70fT531CxO2
7JngKSLibdD/+mDvxrZB2lKnW5AXL4E8B6y4X7q/K4aIOTXXGpBAfQkka2BDMLI4
c4iiNQeQhHSiCkAhRzXSBr9goq7KQMefAUdUPZQAa0b79MBzVu8KpgGNpRBQctB7
p4jrY8co/BpjgeDrdh5nyi4CX1UMUAHtMFIt93PfozOymvcpFX297NH+wJfcuvNP
H72HO+0M7LpHU7tnBw8uQmDDxROYyMHEiPp+2ljjES4tsHf26RSNy8lpTeImra/5
0AnZMb54jD+EWV5BPeoe8WCMZhha232YUhwQXV/9PkB+j6ZCh9joo68J/CP/h+n3
vs93nsgXGXo+cCGsg+IofT1yRF7PKfRk6/LJQXD2RxN54kuRIRxkxd266//mVVh9
xw4tEpkxS7FcfzeykrefWsHJkH7RcoagVg9R4qvhWvjuk/4td/9dh7G3kXJgapYZ
N0RmjjXmgEk5LXT0StnYN1+Ef5OY0EUFOV4s9iZ8V63nvBCCypN14z79x7hfdNr0
eaJrOVXRmPtVm3TQECHONcNhOZGYiEp9VWlxNx/441H4+U0yOXvDbIcFAkjtA/kq
paiPexqW+vNWDtNH0cINbyfBn9E1+TfRBRM906Fbo+IvRHXu+4ewMdOFoMeQz9JZ
GSuxgwZ+dKkNffSESgd9EN8I0lGYUXdqQsusuk7WHe/pDmrMseT5WKifIhBK5Xc1
lvZalgEJSCiHPN9Apc5QfXBFcERFOUBcrPRd4sAYjXzHmasn/acvfuZpshXdKZbq
iOHY/58cPsJPqkcl9yRHs6UsAO/V6hW30CgUaNa9UsDeezEW+gLPCuQK4IYjTaUP
QXo5sGCimmaJSVTXGo6vNGQQEgqg3P//BtjdmMVEcNSEGFXefr3gxfuvsZUCKO6V
g2VnDAu/imiXY2m1JdMqPP6CwX8YcK6XDf8QBzj6x9UptXm4zq3mu6EDjpjImql7
tvD3/2bz4KXiaffMkl8ysEKN+c+Ma65tOucgKBBC/IK4mpt4903bR1wJEJQRJCXi
gEoUns6Q4TE7uCQuCTCDvoLPyw8UFbIMbJoDbGoaBpsaaCeg/EA3Fgi7wDR7WjW3
B+QACkynwKoV3o05qrZzs0l1T6iUih7bPlXck9SPXRJbiW25bV/3w8LB+WSm9vUZ
PIIHtbVSMScZQFmnGrmHp5kZ++uqtjlhyjE3taJ/iuitLGoy5ZUl+qeOUn2zOMqE
qhUHDjVOSMxKYbb2wkvdA77J4XTNdMfJRnMfdDISRArWgPpwqHXfU6k5qstsiKtj
eHmPCOJQtd1RvN5gEZbydPDRAbFas/w7HlQY4wmk0WcD5NLP9mKILEN1Smiq+PZz
Gt+6PqX+sGqQJx8gnrlzEuiR0PjFeb7axlUjru2hUdaRaByo37mr7yfoMKOkVSLd
MK/b0BmQHyRca8SlPY66eDBfI7qYqcKGRefpKfaBVjVQuvGW6nu4FvLf7KrERbPN
+LehfdRWSyI69/vPeJsuzpVnurGLJ4bmssOHpbRtwCq5BjRtw51CDgsla3HDdZaA
QicHelCMrtXEwkIYUPVXIVf6i38LJ+5deDxMBsk6EcXfDEC2eKuGnbkfZnBmh0Bu
bvyZ9QnSIweBBwCD/KGM//cx5vQ0M4m/66quqg3yFmwOP6wVWXhcsWRb2Iqll0KS
w72VhX1fpYcwXuOwfZ3N+VSvC8qWcOOzFAizxYDoDo/VZaIQOd0mYoWLpwBjtSoq
ozqZhJTHEUPgnTnJINpzlzmg+dKvkcO2E5h9s6OKtbH1OLyak0fw/a9G2OtXeMGb
dykoNjd1riXZ3DQa1TJDzbWNzc+utYxdE3uMh64CXtK1cVr+QO0xWxy6nP8x4eu3
qYtdJIWhKInbk1dfbcarH4sqGvkavvJ1XF83roLMsMMN/hwxBhrjV+jjRxTrxu80
M0xHGEVawOaxfieqBJ/vpdPeRJDbV31ioDf/8Ts8PaGcQrmw2wGujBSAWW6CNhPt
eASQEFAltc6e395FvbtI27PIm5TGnBQRz8SqCCfBhGSqotLIIWEE6Za7LASgaW3x
QYcC50yxvFoiIRESsZLul8YSMtpv61+orA/uh6Q4+KdhV+R3guJbPOc9CkNZpoQL
xpYNWx+0iACwUJWjAv8z60ryKbCFrIAhQIIB3bCTgT9y0bmlyUoeRM9So21RTJlJ
0YM/bPkbEHQW48/n8OpylLj0i3hyAKNfAQrEA4hjiRrYceoTi1DrOduumKuENj8d
MODUrb2+e7UXkoQE8y6m3d4c0paICtWmXqeEiBE4oTHtBhC36HV4GY8pTGweR8B9
gRIGUR2EgA6HPvA9BPmybXtrfnAUlMi7/MAmLlK/bA97vH/osdEyAyv1DBbMi1B6
uBc5bXZWwSTr66wALYYII4MZQiidGTXa3iHsAX1unlvhqAgRI6HI73v0uMF8wOpR
UMEAcjRy9r5URJornM/ZTg6GxWKxXx3ihHJXlX5s+3USyT/YgtUdldezQ2T6w4yW
GU1zUFXTVrlEYev/e6LbvfXtkfSX2zeAihl9o2G5+OTuFJ5zErA+vOra8nyBNi81
RJIOfmTwqXVQq/vN16tkL5WyHMS7b4/GJwKqJryEX2NUB9Rc08W99nZ8uq9cvl2c
Md0/HzNp8qdMQqrrGmkR0goWyEMTmJ1rvdHzXZIVnu5c0puOVT5RCDhYHazVT3V3
9qlffNQVY4MvKsFN0Le4Mp/VtOYITxI76uoK+UV882Dqrl3C1HbWDGGg8E14xIt6
zVZBfOSr5OpklL+aTLWftX46Injl5MSAM+9vbLfkOjbP4sn9HWc1JZ4UMFaaG0ct
apf05xYWTv9aqfVy7fmt3jQFB/OP6JFFW2fLsapq4WQLU6uloWAsLt6kQu/40fW9
l2cKRrmLRk1CDtbpRQf3GUfE2sjcq1OkaR811llJfZA=
`pragma protect end_protected
