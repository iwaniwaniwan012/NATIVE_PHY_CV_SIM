`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JGOUyibRvA6hxOVYb0l8tp1biIFpv5nw6luR2yWBElU8JI3Jtjt3+15ZL5hPeBDU
8+tX79e6LrnhCCof7OtVV3AfqH7kh1IsgkTiISbMcV8SGxgXHkDvxADVEiGxY9aH
YqDxDLSShvmA+tGg5+g8hgw3wxNV0xPHh8jI3jz1mqk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9984)
nHaDLgVq96y26Mcc31l3futbkvs5MEedXKxv8rDC6C8GAMgPya+ZYete8MOCBmVN
gx89b/HRNYe/Ichuc9N3HVoXmY7RgynI5rz5aq0zuIwzI3BScM/mbfQfXRg+/6D4
8Zt63bp19otyLalGF/3rQ9vaeo3euiZcUv/tkgOTysG8pDkTKc2LYeJciGby7F1H
y09CTw3iLA0wPJxBTGiQa820ThIGMzz+sJH0Lcd7WiG/fIv5aUHUqRzaF35PMmMV
nftUo9CEfw/iH/1ZgEjxY+xkgwVaGyKeyrSwwQHHfpXaODDLw2gNFEd/Wv4mBmYv
N8hvmbvxZ9BN0r2RB2nN1/2L3XOVMdDXmrHaObzYaQBYKNOuVvJqbMNixUUYWOgt
nYfltcmjNBTHpRHd2j829MzCpwRTvkx+gzZQ5kDhAxv386Fi/8BHMJSjy+5YBG6L
gtCYxp9vg2Ea+kBpGJYiZD7pvW7EgSKGy4EYvKt/lGVkwo5jjbQMr4fgReHfsjWi
L/RwDqJUXlhN9JqtsRCeq7koseR6KN98gAW8UD2tW8tAG9V+6ZMuFxNOwHKh+E+i
LR7ppq2DTzWFPK80YqDIUk5dlNs4DPktq4Ug8oAt8HSUcBg/wnI7UXBTMIBdEx5j
dVxRLyIOqfq/TtkhttaxlXVcW03dI30cP2E7lg822hZgjUENr7ID3tMYEur5J3+W
Zxh4/VQWWzmrSCFaxMdvQ8A+rUtxySJs4tj09hHD4jR2/yrETmdxqaVJnr2XFEh7
/sdft0hjoJEcv8+ZoAsarpoMZ1X4yKMockIvd2xcT7bkfK8BqRbLhMKDYrNH55hr
0i9BfbRE6ulW6r2R2xyiUcyQohds3hAB3mr34/MjOdmBvZ2tvfEDIoyiQQ8KnqIN
VYg8B6cLngyC7e5n2xF4pGF4Zzov6PB/2c28d96LdsuxB6jx2OjwUSFLc3vJbCpg
+ENOnTy2GiSvKVXvKdg32+PJi1+Kt8EuZGyRI7pMMm4XBwc+nV7A+QpebS1uwexK
lmACLVkeNA/S4ClM8p3k/M77YO1/xsYDWYtLeg0QUvAnqqFLKPYmcbbNgavzPYxb
YjX8kJ1xotlbZXADgWMdoao2toS3s9dv7wPNJfb4z0M4R1n7DcL5SNfW6OpjqVZd
lNad+++AfUloHwJ7SoAZ7Od9ShT5f7J+VLtPA3r5/Vo99iPRAexx2v+LV7gDrgXY
0Iow/lgmKOoBAMtpAuLWDcuwoE/QF1F19kLC7KQ+IhtEnOUNrhN1F/V1YN/2+yaO
aKP2P4tHXMrNEdSkZEGnyaNQsKpZ84GD9xT+OhFXFuOEZI2AF0YoYiNQ98g7ZNhm
VRQyjGsXWdtIhUQbEKCZs3mhP/0sLtcWrPqX15Q/Pdwl8y9RvjleFT6h2Ogx98IL
xJ8DdUSssOtMRqksH5RO9XWajjw7z5c1hnXTncyVHEmOKuasFqYnmCGKM6Gzr1M+
NVCHwq1QrsbNHDWqJY295UMuGjxoMgwNY3VoT5zsNndb245oFEYugxA1aNtLZ+Vz
Bot6Vp9MYwL3eWB8nGIEtEzs0NzvDOWQNsj+78ZfNrcAbi0uA4ZAleqHS57srBwa
+nQhDv8zBiaxNcQNkZOmcRCZM2kPmMyiV6Of6wVOQ7y01xETxMvP4i9pL+0yKKaw
oCxZfRGvhywu9ryOfV4Rt2byDG+6lfGpD9Agne5BBjtZa7Dls6Lz5r6vUGNZvFKQ
f0GLk/nPPsfmRsaR8WevlLe35nyBP2+N+Lh1oDsSg0+XcYigxk2p3OU53EXmeGQm
OadQgoWSQYtqKw95w/J6BscpUjm0cERLRAATujw7LXSOyQ435O+PfLLfYo7s2Us5
bYLMyMexPHFZJNuvawC1hMP4l/FFzde4xQzVg7Oh5Rf4dZuI6HNiOBKxBXKkSc0K
31/z+vlRhTB9YWVsAtdcPWxHeZ6cUUDCco5T8glAA20OpCXj5MNr8bqvR01yQi2O
0mEUZiHVFGYN2cS3nKn+/Uxv0HJOxiwBsiGXsCsLMe9THmJ+RJ7hQfQ20SXBMbZe
bIRSczGNZmdWnxXUX45q7j3RH1g9ILYAuMUXmvA8Mf5aHMaqWXMwM3zALZZoydss
yaVgS7jTLAkSsN6DHTRCxQnFFgKWyz2fCm6uqq8CgWyyOC6yszBBTqNSOQFf/aG5
z589DHx8ZQS3T2VF0dnx0VP9MxFg8nkm49+WRuo/93QimJ7ECRKxk4od7pkQWfkH
1Q5LT9qc+fEvQWB+7XBCWlDcRaaoVEN9AoYH4o4qcvc+awVUHfb2RKiWzI+tvsEk
/OJaVev33tYvW7Svxx7/mBKCtS+xr4qCbsV51OdzapXdpuwEJAfRIt4AElgyqEln
5TgPmYay9k/MRsd7SSTHOt/EeSjDroJcna3atnDGYWDUvGlmhABcoO3ZJPn8MUYX
XOaQb5gDAg7E2rluG1LKv41F/4y+oxPyg8u/6smh261ypKl02fiRaLmkdcYHiN/j
1IV9vDfLkjxYhqeSaUdPBFr2QenxlvoEFsiG4/YrvGL2qOlTD27zTH19O9TWGG1/
miP6SBrbzHnJ2rt5ss+kKr0+D9APWpLRfhLLNzFLXo0TDKP8vDU/gSBxGgd57d95
9RA3WkFTa7kt/sfDAdYugrfg874P6rvspm40SFMY0dMSJzzgQIUke25oOcf9Mtn8
X9a9XLQpfxO2g1ghJpCanDTaFosTHIxrtUhAcLs+c318vZNCUkWnNSexIq/9vrF0
5RXhb0tShqYsFXhlfi8BAVO6WV+JSUHx5lIZD3NpcIrTUOyq6BbYzeJ1hRXrKYV5
uzK9cL7sJGo2AcCncPPJUfjhpvjQzRKAWg8EfRhwu50JM0t0WSB1wGQgFEQsS4RV
+7/A0yAD9SAAhoooQAfTnCD9LpLfYxIvJBUbq2i6pOiTvGSr5TN6sDduDryNanlZ
6N6Vezh9iK1wdhEXsVAHnd+BzEtvXG+BGr04U9bgh6ovoG0Hn/z9rTWq3ufPXOdn
l274nmUtoRoMmx8IAK6E+UzcNN33P98L89DX1Utep4Dc6Lny3DRfSHMel0bolYiY
WWoQCpjFy9Eo7AWK0aJtugJ3cpH8MsSAIS2oCRfxWTTu2n4fA3VVsRR9Ohmkf7l+
1s121+7yEAl4N5aeOyeAc6MUpCzDM3BBlvdOUJQl+HOqUa4xk8GSnC2S2AM3i/Ly
Fqdb5fE8pNr9aFWfrKBw/TfhdFMKbY7fswQyY6qHAjUIWUVBWbIBbQbHJNh3FZM8
7KqqLd3vhtu8iMhbwkBKmzQAMkVxAlDbcO3R8kxZa7KDYJnhAD89xEWdRVoTYuhr
my1E/DsEKFEhr1hAxJ3siZDuE4I48CdSyfqjKWcu1/+csPXrmL1d/40xn5cDTabQ
f7pEQfwZ6v5eBKLBb+tunb6WoOuZsmDt4IU2IbpPcrHx2ZMJUsWCteA9UDD6/PTe
AFcfZZhvWY+WsgH0iKS8D6DmYBe0htA9DE70BYvpl7znGmeHGHzR/FW4r1UT6/10
Av93Gr48chZqgFA0UzNsQkk6LeRPbIQGABvsDJkNLpVfC+gcNbQfL15lmRvcP5sF
8vvHqs7gkuCxDo/ikmSaymo4gUd9qdOJrqOBtXONrxKYOnqZ4uQbhmZdwbXdif+0
ygLot6UokcrpFAuMYNihHjzZxEkvJ6imVUueeCu0f+4S5x43uPCvoY8u4Chws3+4
WsPql/9HVGchz2+/kFzJy3YbkVdZNTjBjXboKdXAqdnozwpGTGbDl34SaavaszNN
+b7uEIqmKuJ4Rp7TBRau0pQj799Ckcst5/5LMhsNWlnYUVp2OUmzrq6D4hc/DY5/
1ftbZ6rWzKKcgl7Rcnc9NSsk47NC/+zj1Lg0Z1ui719OUBgJA77Dali0Wu/CtnVw
GMZaW3B9i5rxoAiSVgmOqJ9MnsbdtoCxjmCOgyMAIBAQWSc7lH5Dt6nKa7q+5n9P
KNpTk0I8KDXm71FlILUgJO7/cPMTbeVSt+VWika7O+4+8YqPMNaY8db/u9aw+zD0
4cYD6jvwceUSWgpv73jHF4HO3WzTVZJQgnxOVy9fwynv64Tgrw0y/qCNrIpZDuYe
uyoCMsMMiMSVSUQ5zw7kNVtGVCNN6NUhBXcrLpLXvlTuFt6CbTbdcH+/O+5njORW
lk0ecEgzud+nMZW2oalF3ga8hHispthkkfHHugjVfQC2VARjkB1wYtoJZ7sMs1gX
28Kxt0uWr0ZBrnovrdZrSPo753BQVZmQQ9j6PNI1s5lkWBbbM2Uk8s7FrmYFqZfV
cMkzW/3dnEoC8lVb/0Nueg7qcDpLlCc3uyNiHV045tF+tpreYTDoXZ7aBZ6D3sL8
iRxzkTiAr/ftxYJu4lxZ9hKsx6A4SEs8NGGufy2hB2BPuF655IMmlXpAYbtrS2AV
My8f9Aw63j1Agj7jGX3noJ5CslTB1rMi49Z6XMK5qwmVZesu9TxeFRBe1sdupwgf
qxeRKwaAXhU7m2g+Xgh+A3X1/jJNwjA1BCQTZ3T45lP3+PXiVJ+GcfRKgs6PF0up
PwNmrv2GM4GpLBjN4ywjH2mQXSgzFfXpNTx5FuooSbgxqb6xybGUdn+dYh0Oo2pq
K+sq241xpDev7ku/HKaewuyPfI4NShZZ3GZpCcUb9UE9kY75K1+m15+bC2slCjsz
eHcdhbnlHwJjIU1FOb1fHkSA42VNoEqzafje9pnyY9B54Hx61XJWWGV5bhTqajhz
BrotuTvyHjPKn67+50w5qn7uvncfTMs0EVxHb/N7+Pd3dW1UUGtshaSzFsy4n7nc
sguIe35koVIbQQX0jNCEykfKMRSC8/0RWwPThkbqMgqwweio3yirrzc6CborB3Hx
t/0TMN2lgi24e82nmdFcvw+Me8tAUS42D7jXo05NfcnoQhCzwAlKzr+wul8tjYVQ
FVGau6gFyWsNEocVUOu1MBdq6+DwytXj3R68xFsspgVaKHJeROlIj/39IwdA9TKl
jZJxRrj45gyCHFAtu/fWFZFcW31SE7Rzv/phzrsimuFKOvZlT6TGPYCmcHjuWjvG
jLSrovaDQdZfT7dstqL+S38EnZvu8oDbbq6+ujaeZ8d5UygjewJ+rpVRJ35v4sKT
jbgQ7xMt/l5R1CzsvcSZ5uiRhhg4iOtOGlobA7rSsW1Am2dJOA7GJzYF4rjHwhpT
omi88w/vIWJqH29jG8QHMDrhXm5ilaNbWPUqpu2DwQXXzPtkfXzBMZckv7sG34NI
eIg7a3gS2TsJKvkzQOcNqSO1XDS3LXuDYfQFEe8xBmoNBPFI/UNFta8emjh1ZoQO
bHintI6nxdbC2Y+Rya1X1s3n5/ygGSV3OdyPzgx3YAk0ne8IQ5TOWfTm2QW54oIx
s/BHuBfLJCkADNsCn+PeUsp67pjofztH+0Tx6TIouU9j1sI1IzDIv6vLO4I0u7HZ
evqyFG2RGbVQG08R7khwMfuT3BqcaI3rUwMryWCIBeffz0wYF2WRzVljwGn4fxvp
ehfTXx6wN+JwJY+MCYk7/GqmGlccu3NvqJsT4goSnhHciylvMLi8uNWwnL8jm5VR
HE4Qbe5ldomQijqBg5UFc8ikGMNWwHvK/HGiL85YYtkRTZyD3Ty3eVs30064fFMP
+wjL/WjPvk35qHGDjLPhxY+DTAj85/3vC9ZQ5pzF4uLfiBlPLGGTe8FxTlCpgrIU
jx+0HTyRscaflxu34TU6R07daDzJj1yE8q0FrXGDVNa3hy4V2tEHlpjzG8PDvI5Z
5w5qf/0u8SCsCM/NoUWxeczFQ2FPAeMO1oI1Mdpj7KFo6NXF5y7yG5tZfHhR0cCe
8vMtxeBvRyvobRlphd6Hg0CRDNGYd8zWEATlw/Lc+Rc12gusgDnLt0VkikGkS5gO
UlGSWsrSIdgytENYAbisFNk+85n1cGrWwcGJcJ43TQ5iPxndNUxYvj4mMLIT+Gw+
TA3e2K8KP9fE+7MkWjy8/hofv/uSYFcdLN7vdhuvcYuI2726ZwNu/VVGXIMQNqc/
BjfO0wHU8fYaoDgy8sdVLZrFrQux+v57O6iUnm/vyRR/L4Hk+BiycTYslyENFu9d
IJ0/LTRyIfJTr+atjN2PbElLaPkLksEU3Leetzs30sL6KVvA5PaQ61Grv+Ec9eYT
dLr25SHKhdXu6lgNo2dbNARWORk4+l9osT54fX957NOxH8zKzC2HQlwB7tk64E08
4yhewuYSxwn460RnnozauZV+0KhMZYowVZHNB1UncZKvGat3Ba1WS7C6fi7rep5A
f32Ysh8sBILwXOa1CWfze4UMyTQIDoQm6wyWEeKxrvyyPYuM1NGXnsEB7UUNn4te
DuyGLPxHqdscOiTOSQzFXI+IfoXYhx9bPNXAgf7hqc+4cluyGpUVT/f/7PpMEQFG
bB9E/ccgc2Jg755aTpcWXQ5Ys12onK92089iAK6WgEZ49sGd/FifV7Pb6OsK4C7e
A0rHP3FwbzKjuJkjSYO68UIc2UnKt4MEgHCgaQBXESgovdFjd3pya1QK0AR79Yod
+Xn0P03QD999sPva8f+G64Szq3e+j1Mmc5U0QVvy1W/8EbGjq44ZY0tg6w/V2dsW
ROONhrnPpHpu8jIb1Ya6C2WD3zoaqIeBoV+yukLiUoTzw9/wHuUd6LQfPuN6KbYU
IgdWD7M0VCgRGFNskoJIQoBv+6TmwWUmBbLgtar7OVdZLZPn9mMxrjiEU3aSi9ln
606HTVzrDdf1oq6SvjRbI4gjyzfJSdYzYg1Smb8v8MglxA3XwcsQWW3S5OzZSMvy
VR18UzPRp/H4u346G4ULWJXFfLXn7hBlC60Y+tiqnSyquJJHSw69/WjXnICXC8NF
KJn3GlXEYvQI4wfUnO32wTOFgxXDLB3gX1exULymVFlrRo4X2QhvVpEFJD9vnBfU
r0o+I1q2nuBD1Hln1GL/LHuUNs62k0oFSy9hXrnQ18a4ilI+BcXbFJuhde4mqnQe
Jf2Cc7ximl4M6wjhgm4xNY0GgQ2Xv/j/emvW5peUb+MU/VZ5BnTyOj96q8/vHigJ
F9YCHjulvCmB4sP43qlzE/pUNIkDBg/FXQ9MeQz9hg0n18RIv/ZLypj+c8eeRwcw
fm1VY8icTIZo2k0wBAPNIiVdPD1sJ+kXU6sXh0ZsTeTWho072rfkJCWalyxoVT/M
F8tcoOmiRQUp0p/tB0Zeq1dmd/GklxylhYxRsa8UHb/JQeM1xznNrGOO6YwJ2Txf
PFCo1gIIgAw5qs7/CYx3V3H8I50Aqs8mh9hJYLeTsotcDiXWYd7wYpzrRnsn0YnK
CxP/lOzexVDeTR04Fvr1d4fnmmz9k1ZOilafBoySYldWQbg2XrE6sdZNSmr8WMBO
tvT0MTnfJKr1R07A+DLxH+n87nUEfRCQKO+p1/uqEHyTSB0Ac67qkWPCkg4Ix+yK
AbmdVgNirvOqDK3R/Debj09f/uT5kZzQLr4mtEIxnaG3jxIzQzGZrUFah0KMDarz
kpmmnBqwDzc16M0ths44GYMQ6GehQgkINUXwB+6t8eVjZVTT9Qht0aWrk9xql7a3
qofSLLmIdHqkkywn38JrTnO3itH7uKKoUENAN5BcF3Um5H9q3mRdUAPLUIHLkFga
Xyd9T7hHhgULkeRhaD09RKkBZTBJt3Qsw87oSMZZ2TZ0q6UVjXZgjAXuw9MGZwhG
g3AU8T+KSoLFoVGsvTAfFbQycGQW00gmj2p6O10rlPzS0Mwy4qBDKAaOa4MGvotI
bPD21/h5wExQ3zhxWaAxEgCivVHerSW168TE7D0NLQ1xaTFksm1Ek/CyGTbh/vw2
wOQY4E5TXo5NaXA7Ep2hamY/yC3kpywpIvQ4jNwfG5xhwJh0gfzkxNRh8FHw6iHr
+Lya1Q2Xt6VmiJCL2Z54o5ha/rMQ3chVRX3eE8XISseUwoLyYQR7Ni2iWKRU5ZRe
+e6jDqL2LrV/DAfJyTX8fX9jWTx0yFz0hPAGQLwruwHT+8WzrOAsZXb2iSZmzm2m
Up9l2D/HgjfZF0GZq8gfLH9f6k339rDGqrvgl59ijr/AX3B+2+m5Ar++nfvN2Rvo
iSYBY8Sd5cFWKpB98MF4eyg+/GC2riNR8zECq2+ZRh+/xhnQbRmZRlyvLKKVWxmP
g5dCoxICVMR4nPhQmHLdbesIr/UyYqQjqYXBlE7sJa8z3AfiCf0JTTzuPpzSpqC3
2lH4aC2mrOjg15F1kUnVwUhQpf2FYH4xLw23Ey7uo4hWp2X3SgfuhOZLEYzJziG7
vxPzRU/l0s46MfrcrteVYveMwOXllQ8esw8uDicPBZ4dIMa8kv6Nf6PNVBuDd5fn
lQ8muhRu1TFy211oZ3/SJ84o/G3pq/+ZqurPLyXmwJCtMvfKYMwJBwND8kB9misB
UCG5uflL9c92rRDgQdhlzXgtkgQjiEkaq9DvchodkITbprE8no6WxPxh+A9Gkt9L
aQYW+haJ2J4ss8+brbxKFa0jfJWpKQpK2MdLuyIj1wpR/jFRHcdO98dizDFaBMuI
Gyi8ExuDAFGTwnR+ryG3NUkjiM1SbDEktfCpB2qbG0J4N8FVKANiIZCyYcDNqVqD
ISGhn4sTTofKrh5LZk+ciAIfi0ZX5a/va2MeasqtExDLXvGkzGP1uJIi9uSJji1k
vBhKeF6v9Rmzayrrg2ftq7rXNkVdal31oJlG9s+uUp40RVxxOrHYEb9iUkUZbHTk
qBELp7LTTqvH8lGCO/tnaFI3nHe2fxawCsX/wT9eYRlX983V5uyut24xPHk6Z5bD
Gt6f7fln3B5w4NQbQb+Qs2371Pdt4yfHSSkfdq9agYtopbvFBMi1/oYKIdk2D9Hp
azZWRzA3X6QTgSCmjuhISIyJt9eM3JaPIYOPerupNLcFK4hWVYBql/PBo2NfXwE0
rk9H2mJeF9I+vDizhP+OpcVnFvcBc872tHGP+bq+RKM98jvhhuM4RajDicZnb1zt
vUthXt5irEucyrXoFETnJZQXOwj+v8uh9rTNt8kLGXmCUAdUARaR7xELvsmAWUaY
Q/TsCOWF8ZA8eM/MDmMT8ZWB6H/TpNu/NHRm3vqo5xnD6o6Lk/UJmWQ4ovjjJjcL
hoVfSxykb+ZbvDmbLP8R3p3HTWxyXQDUIZvXKfcMwUzIDhvSR7XhbdsxogpuPtLf
wKDmXcuxvwRm8yJtN9heu2Fu9HOLAgmIHGloYVjVezZPYwWCKdejbu8/lRYfxR5J
ehdU3vJsfxnYYL8BmDSLgLjZlVxNiBFHjHmydr+H11wCdusG/yJQ3revaqTQ+ETZ
Y7Xai8kkCGMi8cj9UxnJcOsxhRRV/kahAOr6dDbSJDj7y69XT2w6YuyUHBIIQyeW
NLA10sjrbouTmzVfu7430SRQDdDhPWqxdtUrEa3hal/b9K1+lZY1CXt1ie3K1LgD
wTE8RI5YsFP5tH2BICbOo64qRkx2C1kBoU3ySx0rMhDNgq5tqLq40u5U7b5WQNgr
ArF48SUa2fbYXY4+N/YxiNKkzY7Ts3V3mwnH5ABBGAfPtovLJV3Ejzg0teNagp9o
xMqrbKuQqiq0ze3MbebBYpWaadmKbz/PDp8MXM/5bDP9cB9i0ro67JFmFJJDS8Gi
L/HSyo8xLzzWannW4P2qE6GqsJYIlt76meKG1LBaP/AcwyFjlye178fjiGEQLtPi
JeaULzqeq+oZtiHbqjo/oVqhfsEbpeOczly5cr0FX5wZHZlVDMTO55e8f9wB+B95
VVANg8S2PvF0Ob4RMYwP3G6ua2r4SJ5IDwENshotS6yUggtrywlyYeF3QxV8GWHj
tOjj/M/jx8CCGxy/1WFYaCb0qOHMLLKPryHMeaiQP/nW0Rga6k4GTdXNPw2evGgy
6aXQhXRku2Zu5aHJ7ImYifzLkPyv3i/SAXiZhvXhCGXrzAhWWaCLBCxqPpx9N0Qo
6r+tb8eBS5ERwoyZZGoQ+NoSbm5DebkRVfnWQLpFrMcIyzP6OHMF7/huoV2nSjTd
Du1hmszuYxuPzQliYsP1AbnSp9cs3RS7KqH3OdTz+RtdJvk4W1fHYmdw9mRHUozl
vnobW0kYLK37wcqS/cX17PVzNiP4JmwTFBexpexGtT1uZL3d5BycrD5CBLxvrcF5
iTHqzhlXOTtcyKSmP8c4GINW5SVtrYeZoSwE0umE32Kur2N0bWV+x3pArCLTvQDW
SC1jPtleiHdh8oTkGCyn9BbLJJcavTKSH1/jTYddaCce0hwZAt7aA26eN//WYyhi
ahE8trSTvMEpW16xsq1CyDtwaM7j+nm8krkUZkj6YpCzzonqF4/6U32TQhlEozRJ
09GHMcmrc86wiz4XAoHrX+TjVJ1obP5+nhvVOI9pqysBSf/ajC/zATzuI6J50zPJ
PP9yN2uWnHxlNcU9s/cv4ssjxhbT25wH3Ivdt2JfTrZNHX9pn3BSsSe4Mb4kGpIB
7CfEMvtvNr5rdw94Ktb8L91CdIoM4wzduy5GLAGNwjWhk/cT0Gwxso5uth5XE37t
CTSkAWwvyGTXUE4+wMKQBzj58w0p9DbohKPTNDXgJvUgpZrjTIhqMjMkSgeZ6dFB
yblYDM90Mti8K4vgnQoZFw5K0oHz7mrPPZMp4n6qN4Di17hwzMh5tnJ5zzVAu34j
ot6ysr4XbwGGR+YvVlH6lmxzEfuPOBAhuch1h7G6ysd8rvDQZIFAExofUI0eik9C
MHiyyAvMuTS3x8dn1XadBrG1fbuWWbTBMG3XCd4aZjxEXNssapbraqjzzq1PKwVg
KhVngtGGh6EcaXowVfxjDVsifdl4ykWyfoyJFYnJ1AD6WElI/6ng5GbM+SMQfPaH
4Hff7gn7FC4fOVIWLTxHu58qma7Hit0QEVISMe5h07y2xyUptJgMCNaf9HlE7F3j
FrQA6cdIdHci++nbk7hPuI1hEidkvXLoa7GtXxb6xwu/zFnTYiGuNjfhx+MXWxqZ
7jV34lck03o/I63a0q+feqBwxv7TKLq94BisOMqMNHGa6s/V1ma9rKf1W8w6BM+B
POiU3dL4ykPPyctibESfs1Ldh6gXElFMxL8p/w7fFs0c7BajqJS13QmdkrgFBECc
Psq7pWf/FTDOxludkkkn7AJVJ2FWhNBjCxQQvqSfEwm42vr6h9xcFKz6Qs3fNpny
lX+5CH6htH6ODk05SMstYcC/Zth2gqzT9TuryoCGozEQI5vsHLMuzitiLjzLKsZ8
tJMkoqJ15q64DFH77hr4oU6+2azshpIgr/rlhoxJSBZYnTu64mkXkDVUSU4Lzvv1
9ud/Bq3z9zg0xJ6dUJkAp4z5i9ka+H6iNCtUS/VpThv9y8dOK4z+Szon5KRR0tvy
blbdlMqxCieTUz0MBCJ5faOAqNI/My/vshIOkYytSXNsjs7eYwlzv7AJOTTNfJHV
BnxyKiNxyIjEDrD6fbsEDaRKS4PwcEij6nHK1BRBToXuOCB++TT1DZ6yG2+NAl/A
gp/gdbsNa7HwTxWcGGW67X8Kdbh38z1XDLHsSyG2Vs9KOshPlGsf78qs0y6tW2G+
6G/uJnC7uxZajjDeNcpyJoka9W+dUpT694uVIWNwax1MvzA3t7zoA8ADyQYKJd1O
1ZE6ERclm/5MUzQg9EeBB2/NKIH/W7hRBdJ4XNsNHVZ7wrn7qcaM7UBQnO4HS4gs
3HQEpo2ghxAJgzkCBNF8LoQydVLxPkXUBqLwC/3346jC+4TO4xIIDqtZkjriPK/1
guPVOJ+Kv283U+yMy/CEB5gUwS+qCKNg8joJXU0uk3XtqSYaGg+AM8uiD0n7Sthu
jsgkn8zmidgFFvn2+yJhzUYzIosNUBsUBseDCw8KmEVm25jOx6eRPIBdvDFbxqwF
+KRcQeS8e44AZydOoGKUzUqNbhWa0TTH0QzEWVjrV9k6Ma5g5SghLNlg3F0IjB0s
wCOYsO4MaaL10yakv5tF6Lpvsn4vlxsV1gQcF1qZ5uh6g+IuZQnXqOeOeaSA/H9r
EqVoiIl6nJ+XtT4gywsL7Sit1aUhXhekAzgSjyIKIZ5/NVnX6t2RFyNDye5OHTas
Pqj659HNWKfrh0Ct1/KXqup6656yDeNcZczRA4RGb1EMlWjxwM6hD0/zB5lYyHLn
GHopYtzcOlRjf7+bcrPQjn2AuvBtzGpUFmqpkovi5fbJOszI4x7Sk6ruptiajPkd
8CSpF7MLjuDdXbgKs/Loq9Y4ULBUdguHSBRmXwfBqrrxUm9N5d3lYhl5hTMtjYPs
b913zrnMRDQshRc31ROthUHMOvcWk63xalaJ5gLxr8WZ3qVxFAVu1S61qTsy72wn
NeRQ13q9Ajy1xWvb+CNT1NvPnwYabv7SWfcalkr2Akb0LiA31VsQSpKKwRvvonf+
MHgEN5Sk+TR9oWX+F7M2L2fX0fTN9SUIHbu541UkaO2rd95wsOrmaXTLBuoUfqMC
zAg8k/nbjlxBviofHnQkYribB3fpVoekpZEoJmbAf9AiUsh02ErPHmaZfLiDcHav
Ige02jGoQBH+piMGge+5nvqJeebu1/5l4Hc/cQK+q6n8XXQJjoPnIsqEmp17bGSL
ORexOryOpZCNcumqaRBmO42ob/x5djH+6tYEX4+KcwQlJjBu4LHUFqYfnM8+HS46
UzYajCf2Lut22HFVVoOCrpjenf4YWTotCYYmBUSZUke/ba6dTg/oxc62XIj/9zPi
fQ9ySgbIPZljvij7pQvixQkP6LQS2tHqvMic3YejCsZB58J2JVIqitljK3HcAWqt
Re51ge7ViqAN0AEcVh7xbQhMhS+PD84iD3iqWXS4ad7iVEI4dX2GlqFrg2PGaq0f
GddGn85+ELi33kiSl61TiWkzQaL0GmF5h7V1SeLUnZkiOVVJBshgqpznjeJm59bx
xBZ1g0UrxxlTLV62yXRxSZBN/2AGY4Hi786mXs9CQlMoLO5zf1BHahO6lNsSdtbb
HD+MN5/99qA/eIWGstUF58ypFHzS+XVIyMB5xA1GndjLpHAmKnsQGVsRELy6sRaB
jgt93NTBHi40cTJ+Q5zaTTrF76OVN0D+u/GRJ1RXxD/TTkS9ZN9Po6G0stoLheg0
2KlCkrOFhdOQL/R/gzN/CoaU3zqc+LCjUo++vq+ti7HTC/HeFK9woXUS9KoFKRQq
SNL5cHXpXubRrq9Q3pTPYW+kofEcXrAPF5i6QEVcv/gJZHhLQSR9myPrGc4YmTZf
e5PEurIrHlq9SHWfORkgAW5HJtlehzznPQ4TSxaIzaBniMf7A09EHsDOsIzZcv2f
6AdRAk0orMDwpQygEO4FUdQvc05x3krsln2JzClqj7pz0SQJhk4xPx02f9ft2qa3
`pragma protect end_protected
